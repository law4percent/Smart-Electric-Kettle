PK   �u�X��j�  �     cirkitFile.json�]Yo#9��+ͫR�}����>��l�@�C�`�٥����-��`��L*#��5=%�F2>�EF��l��^���������<-׫���/����������~���m�?~�}�>g�?�\}\����>��r��3�ʔ.s���.��+otq�f>}��x8���6\цk�pCna���R���,��uV0U���)eT#X	b#��"3k�70s�%�]�2�3W4��ZSaf�Y��J�L�^f�y�+�9_�������Sp�(S����%��A�,/U���̼d.+}��umT	(�L-(S[��225c0�q��L��fy���+V7FK.+[�2��L�HSu
'*n��q�'��9T{F4h�h�Ѥ	"���?Ağ���9a�-\V�>��&+jQ�G]�JXPy�>f%P�#f%P3ǌjfA�9j#*��EVj�3Ŋ"󂱬Qw^�L��qXX�-�͊Umt��Ue2	aE�x^�����l�k��%��zC"l����&�	ۄ��i�	ή�	�{r�cQ����*��CX.MY.EX.OX.IY��`T�R�Պ���h0Qr%��f�k`�%(>�3`A(xfUت�4�I*(<�f��f��5�ܸ��03)�EBH�u�@�O��F�8�� Ј�Em���C����m��=3J�ǝ!��x��W'��q�5<硆��<dR��9I豴'6�E�:��$iC�ss�L���Sf��d��0u,X!	��@�Ȑ�~2@2���q��-Vw�B ��}�q< ,��� p�W��Q $TD*2	���NB�$�bwTlUD��ӿ�_u�W�&P�;^\�K
�Z���٣7�-�x_���"=T���MC%��<��MCƥ!��h�4*X$��i��H�b�F�4(iP,ҠX�A�E1��+>���GR	x�c�`�l��=�I@E$y�ѝ�=XI���Ʀү�Mm'�2�]l������<'�E�:"Ȍp*���m��6sz�l4�4��b�M@e��Di*f,���>���,�u�b3�#��]�b3�׃@l�odO#x#xA&�Fd�L����L�%���r����6����ժ~�n�b�NE$�"�PQI��$TL*6	���O��D�M�^��<~y �4�i ��`��1O�b��"�N�b��"�E�4(iP,ҠX�����S�0:yE�2�`t�Net]��+:�4�2���ɫ�T��+:�Q��Wt*�2B'��T�u/6yE�2*#t�Ne�t�N%/��E'��TF��N^ѩ�����ʨӀN^]��������&��TƱ�M^ѩ��il�N圗s���ݽ��e���ߖ�����!/��~��_o�z3��)y��>^�<�}<J��ɤ�yft�$��$ŭ����^ܧ\��8���uO�k�w���աo�&�6�N�R�r�]E���0��(.�fF:��)%��3#ݵ̌��M.h�����kos�a+a`j�aG7<+ӎo\U������SG��󤜘�B�`˚)�"�bQ�6�s����8�t�H��ry4j7��>�Q��χ�kS]��W���b�O��b���$���U^#,�3@����4:�X�*��� ��-o���8�GH�@L��� F�7�؀��T܊�I�0��kD�7c �� Ƽ7c �ތt|3��q���������U���E~��1ɯ� ��:F�	���k��P�W9x���b��PS	!��o����X�p��n��%�f�yYQ+
��8^�+�xMo���=v�G�@�G�S^���䈺�G����_�ȋ;�Ez����:�H����#��T�s*��G%����YS���jaAUÂ�DAE��"QP�(� ]u���.?萋xE�:�9�IĀj��V#����ڣ�pk��R�<��pf]��!��Х8d�k"k��^�l���e	�~@�1�[؀%�¡C�r���]��]���2�
�ѥ��W|tye�A#�
��H,�.u�mTt�N���:;!�Q�Ur��pXcʙ>*DHt�Q_�ѡ�Jؒ	��bk':�l(�8�YV!���B^�y����Lk�|�A���L�za7�8j��Z���:x��Co��П�<�a�hi�"�a�#D!�F�����4�x_��� �,�� ����QOx�{vp�1��u�� ��wh^�� ���k�{����m��]�龎�?�A��D�M�����"�~يZ�ԏ9I?�E�e�c��3��O��(.�b~��^PO�x(+)OqqiW���"�7u(A5�U�A�?M+A��D��&��>�o+��1�G������k۴��~
�����'�nJ��~�]K!r��z�����o��&�o�&�o��&�oR�&�o��&�o2�&�o��&�or�&�o�&~X�_~\��z��z�?`���bS�U��7���Y�?,��;�:�r��?�m`��_}ܬ��vY�X3��r���.�+���X猒zn�\8���@*��
�R�/V�Y�[�ռӛs����	_���ǩ�7O-m>�At��W�*Ɲ�֛%P�w�͞��|�����+��s-���'/��)f����=���n���|!�a�]vtV,�S�����N˅��3���HG���ʊ΄����3���z� �S0u���\*�_h��!�aR��I���{T����9��&v>?7�RJ�h��āS�[Zbn�].������}X8�9xƗ�2.aQ�~��Q
�`3,�Ѡ����.�aU��B��fX\΍Q|�9,5hf�e���Y��8&a��`3H�/�n�#e�Q�l�:ho/�"� A��}nA������s�\�Ќ/�B�J��l��x����3ۙK}��?�̵ֺV�Ȕ- jl��l���sQ���֬��QY Ķ�l�7L_�IX���ť��:��`//Ƨ���+���X��[Q��e��
���碑�2��,��� ��g��妰��R�ܡD�ʳaD�h\)�^��[��ʩS�a�2�$%4�W ';k=�Mx9auQ��
v���M��t�}��u.��9�*)�4X�J��e��.���.�mcWR��fWR��o_�=aY�4�2�ԂYƭ�Kf��7���G:ܸ�[\�������P���k���+�=�҂}��k����R]���b��&���3�Ԯ���Aq����Iw��P7}ip�æ��).a��بz�	�M0�Z�!�A��agr�9?*7u�zL˲���s\7��1�\6����mQ�(G�+G�X���ɮ�+�k2)�|��+��̭�������\�%X��4<�OQgV׾`u��bX=w�	uD�BYG[��5��P�b��##���0�dt&8u����n���|��8�]f�i�;x�kؐ
���s�W �p$���Пs��KeLcsY���Qg8��!�>��ac�[:
��D�$1��q��d�8��!X����,+�Ol�R��gQz�V4�	<w>G-'�d�hLX��n�- �1{�_�"�����ၡ��v�\�����sh��~���'�'||^-!����������� :���O54>՛_�O��>~����y��a�����5_=7y�}�ԛk��w;��*o6���_~ZU�a<	��Kl��C.�܅�\�C4y�a+U	-=�4!�@A'JU�.���n�s��I9�ֳ��6p���9�!a�~^U-2�kX�Y�ea�j/@�
��!"�B?�۲�~	$ 2��]��_��߃o��q���������A^~����F7�v������������Y�jǻه��o����w �|���\�T�M/>�m�ի�*)�qnKj��%%k@�?�q��^���헖�����YH���|��[�)|��S��?�f��Uwh�����O�>���ک�s�*�j��?�f? o����QЙ&�q�L`�	�M��)�����]H���29v3��9�v���q?�}{B�$��&�X7�����`ʎ��.��br�����zhW��/��.��t&p��:�)��Yk3.W�%��V՛`gko��]��$�����e�͌�;�-�p7��9F|�	��r�^�Sg.�}8��z8t����0�a:�O�XK%�i���͠��<>D�z+�+��q<\a>����<��<(<+�R�^��N��W������[cw7�bvz/�{	=��}w����1���=lH���������VȘ�ލ������1�kF:���Z�:���D�v0�7���^1��xu&��}W~�V����M�!������^����}WL�V���������z��0��no��)��Ș��O����\�ᛙ	<w7y{u�Z��:Gg��&sk��^$�ӭ�VL�s�d?�W����� ���t��lL`-U��"ltO���FRGu�A� ,G�3'�*4e���t�d����R���_�*[1���|���Ç��;��^X�dr'L�yU+���T�t����n/6�K��KW�^V`��~��f�k['�,�z�� B�O`o�ws^X�e/���/���e�ܤ�k@�p�c �[$��S< <o����@�<���}y���0O���^�P�5k�p/�H�	�	���ϋ2�]��-^�K�a�����	����M^)�ý�%|&�O`-|^t�*En�9]��R�&��^�	�b��=ˇ�����z���fV������������?m�O�><=n�����?�r�|��~�PK   #aX׋JW9� m� /   images/0bb515cf-1352-468e-b4e5-fcf5b4434fa7.png���w%��ωm;;��m�8�Ķ��Ķm��Ķm�y���	��ګ��讪O=Ou���"  @��U ���VԿ'��n���ZN  ���D�� |}I�
��g^t=��/;P��'�}>z]"�g�C��8�:�sr7T8���>en��Y�le�U��E�K/���E��ʀ4��@֙���>���gI5�?�#Z�<��
)���G�1���&28~�w�ފ��q�H9�����߽�
9t.��-�Q u���b����w4���Q_0���ۋ3���a)Uƶ�;t)$���}�@I#��a��U���JpA�m����G��x��H��Չ��.�X��˴�}�H��J�k\	�4�˅�@��g;"�Z/68`_�Бƙ����?x�:�T�ax�� ��+,�n�e��o�7&����P��:�"�Ʀ�<��e�-S��īfOd?f�?>��k�\��ێZm���%��2����9)�ض������cR�+N������(v�!��b�R�B"��)��3��c�'�.��[$JR�.Y�,Ԭ�A{��՟�?��YXX~��-��4QQQy��gE�g��\�n��������Jv|{����ҨA� ��z��h��its��>yu}~�v4QI��.?Rz/g9�S��ao�;L�u�D��̶v����p�:6P�q(�ƛ����^�r5T}T�TmG��Ņ���ccV�N� ����]#�.#>�pDzm�6�9c�$s�����9,�W�vh�������1�+W�P�X�lS�Jf�^\srrbH�a�S��FZ:͋�6�]*�,��𢂛-ه��^ G��O�u�� C�I���(b���v�*r,+Lr/1B*@��`����%�!w�����%z�;�tK��)�3#E��P��J8�6}(����jg�c2BR_ځ��e���OuL���3�{��9�]����Q�>�ڏ�cg�2~=�!ZL[�e����;MT9�cU�e�\,JV�p�U���Gy"!��R���h�%^���U�����ܪ����2�7iz|էo���I'X
w_z�t�p��3�b��,��^;p���!�a����߫*�Y� �vQU�F�"�������s �	*��=�Q�o���5�;I�ML�q��}��pZ�ϊsA����q��͓�[cfIs/d���`�i�=*`>R��~��*R׽��
\�u�ܤ�rؐ�d���e]9�������j���Q���2��b�Txʔ�y�+�m�5;���>˶�59󞞝�7��'9�h��Q�}X�:(�a�߱���w_'���Ah�����^����E������d L��$�f�kx���o�=�g�9�RVG��O���і�9dw	���Q�9$�Ne������ko[�D���s��Z�������Q����o;tٶ���e>��c�����7���(�J$�?UG�����L��φ7�?�-�z��X[9�Q����Zn�<]/y����*��4ϝ��{�v�4BV�u���i�3ͅ���1"�iM�p���,�����8V��s1g���{.];h A�� E(N_�H|-����^�aF.1?�W���Q�_�GgF�jt�����g�s� (���O�/�x����U��y�t[�v�c]"��ZϵBD��oO�qMU����������b����}�@+G����[���R['��>eu���[�X֖�Q��p�
�u-K���
��B ����$@�'W�G.��F-��M�1�;�u2�NI�����_�~Z!�R�ڕw��V>U��[ޕe��7С���Z��3�7�2����qԗ����$3B�ڴ	�6�w���"�Ǝ͝/�����)�,/h�f���Rд���^�n�=��X'vx^����}z��C�ef��� ��	�����B���T����������T���� ��}�X��j�l��j�د3���.�?�|i��τ��C,^ZjZnf?�~�R�RE�.Q{�B#\��R�v�yA��3դ�H�y��x"�1����� �X͡Z�8�F9c��Q�jm.xjEr:�}��?�,V��l�^�:��o��O����A`�z���o���������{ &p�0d�q�g 4
 �S�L��PXW����/��Z�ȟ~G��x#��F��-�Jr0!�������i�=���cd���Mv������l�۽"����=����Ky"�GuFėe �.��>�^�1}���g��^�L�9O�p��b�!fļv�����7�$��ċ��5)�mU7��0��� y�X��⹛�S��\��j����E#���������w K� ���8GH��Uw:o�����+/��k�7�_{�7�e��<�k�5�O�n�t���Ў�g4�X԰P�'c�_@gm0y��`�j�d.��n��\�-�<	- �?��_U_�6Q�h���W\Eʮ�Ѝ�`����u���cpwjmhimhh������,+��$�s~o�뭅��<�h8�P?q|Z��G:,I>_������{?����{)~�〶���.E�^
M�R��5*W� �/�.�L
oR@�J��.1�KΎ��Q�4],pd�s��̞Z�=O�]���O]�T�/V��m��ᕧ��� #� +���D�G-����a���}'���J����MTc�k�j�tR�(.5�h��z�viK�^Mk�K�	F�^�����n�/�
��o��
e�8Az����&�SS��I4xۺ��+}�#�x�Kl��hkq<eJ��s�X����{#��4�����a�������|*���I?.U�>���m�L�}u��<o�*z뻚z�W�J!��iq(�N���E���.]i߶��m�)G��<r�:�3o>L,N�+
�M���H�6��4�i@��6�(y��-9a}澷��^Ǿ�:�}�o�M��<���� ƶnWI#��������ѽ#"����]Y<����÷�JӮo8�R���@O�k�s$�-��@n�#㏝��tK6^K����׮��N���x9N��0�zh��<���i��k7�׀���'���������i���Ax�[l�ܾ��KaK��㻘�l�K�a�Z��������ő�6�S��9?Q��3|�Ѣ����^�Ry�w𿽎���y,D~�^k�ׂ�%y�h �/#5)� uQ�G��pg�� ҹ�u�c�$ע ����s��
��e�l���[&���Z'�`̹��aO��xn��2�
�$��m�p�6�[��p��m���`�4�wV���3��A*��H�,&R�?B[nY�G�H^�%��/�p_�v|~s��S�N;̥\�H�|���i��0>^#�0��y���{����a�>���o�x��O��rI���R�ҵ��Y�ޗs�[扼{��@����9�p��\��y�W�G;(�痦r���--j]z<Q�]=�g���/��t� ]�Qh���)��\ 3kC�o`�w�:��ަv���X��p��>�f�c���ݣ"�U���ݺ~��$<�l08�����S��8�wPڅ	��P�/*�{�<�z����>��-7��#�������y��Iڄf��U��핔CF�������zt�͘)�pѰ�r�aG���}��ue�l���#A���k��ǟ����+1����K�I\U��Mʴ",}�q��î��I��u�J����];�H Z���
j�^�M��(-(z�(��qJ%1���F�Z�1�o���β�z�����������t�N�-`�>b�G���z�8�d���[�rS�=Y:x�1��R]-3�e��=7���=C}�&��KՂ-���&e6Ⱦ��F������o�܉ju��P����p�4O����u�#ľ�q(��uu�������j�?���5�:��2���V��.yR8����O�dA�M��i%D++���ӴU7� �B�Jy��AIS�	?��»GsN�6V��,Y����T���E��@�A�b�KMd��]8� ��NM��փ+� }�����k2y㭒w��%�+ ��?6�i�g�u+e��4=ke����:��|�w�/i8��Z�B;5Ԅ���/��htm,�LBh���Pt�g`����ل�O�XN�� "������:Y�	8�p'sd��������ާ|�ǭ����TN���6b�7��5+h�lд�X��t�3u��ˮ�����zS42{�h����:=�[���;Kޡ�[T�D�P��e��;g��Q�����ޞ��ak��S��G�$�1�<-��BN�Z?#Ly�cR�	��#~e���>��<�nC�Ĉ,�ڿb���{�1�A$���L�C%<q���/�p-S��o>Q�L@/� cz�b	|S���<�}2�?x80����qLqQE��6��J�-.Ep�ef�c�^Z�1­v� ��.,�fEG���SRQ��(V��ص���rS���@H��㯚�;��ȗ�o�=۟7�
���w�TS�^�^�1�[�m��йn�$v�A��~oOgy?��>���z��?�ƃ���O��vl�+�(�̜:�[���E��P����6�Tv�콘6�� �>d���4Z��'T���m�Et�)�͔m�"��-U�
�5y�^n�;���%�b���è�c1�A��s����Ļ�~t��$�Ķ�''b�c��#�<�
L3�G&���G�ܦ&�m���ge5�a��{��.ģ�8��Ξ����&�ڔ�o�	���ʁ�Rr
r��h�B}��t#,����|G\��TxQ�!ә\>�mN�޻�/0����rˋx[���运��Z��+�]�+x?��l���_�`��.�#����.N4����[�)W������T__��Ѣr�v�4�>�_U ��`Z*��V�G��j�]�n&	�؀�i=��؅����XO���O�OS��#�F��B���ߘ�k����1�����N��7���/=�%x�!Ō	׮�Wd��Z����b�x��Ń���b�sRH��7,O2��]���Ai��z��	j��rFV������[�y�m:4�,(ʌW\�W$.l�q��h�����j����1HM;ղ���u�Y����4���x>4���D�i&�$xM��}�p{������\���V���U��<yz{{��P^ƾS���nd�pf�4�ٕ�Wșض�;cM@ �����.�G�i���bxS���Ϥ���b�H���3�5�3��C���c�~n@��F]����L�����#��`��:�f����t� ��>�z�Ѷ�fT�3���߳����D���^v�7�O�ET���$��N4��W<��B��"��`����d�3!LB�<j���2/��r�u���TU1����[z���DȾV�gR�c��y�>�2}�Uqh�hzf���{36v�&�*���M��{����x�3
<!$�-�oz���쉹����T.���hzd^_+K����#h�Y\Z�:rխ��A��5��O&5���n����(���BV�"�H���ι����@��G*9�IՐ-0��T��!3��@�K���Ɔc��k��a6ϥ���ii64tfF��|�`��('����E�R�~�V�@�$����.�P� �^�� �r���|f��
�t��pF	w!s���"�La��!
̱ ��3��։<\}�*2I�׷S�P@?��ƃ5��i2	�eL��j0�I�=�y�c7z3�#�m�������a7(��XO��}NI�g l�c7�z��� %z��g?��M_׽�����������EUإ�5�m&��%k�cKn-����=u@�Z�����h>;hM�X���cw������Sh2����I~#������8�c�F��N)�Y	�u������}_��F���Q�����1��.��d�[濆ȥ�TW�).+2��D��Ơ*m����Mz�t�w�+E`��z@�����^୵�t%��� qhf�6�S���~��/=#�D-&Z�o�6�f
�$�J����Ha��:svvW��{��7��,�G����T�r:��@��O��֨� ��hoo��ggI�ni��ԗ��T�������5G��ѵ�];��&P�����d��I��&�OJ ���=[,G ���j�W��g
�������f)USʐF*O~���aCI?�����+�R�ء����һbsXH	K�~��s��'�~�(X����ǟ�䭣��Q�e����)bb\�;rKF�\*������PL
����\jt(/ͩMߐꌪ�xmm����ʵ�����Y�\i��=3۝��w���(7�*���g����zzo��=Ӯ�\�g�$�?N��S��	�
Ӡvg�/��)oI�HK�O��ㇳ�!����Р�Lu�ј����,�A�z�rytpYH�"||�}�D�Q\�l;�&����38�j�FLA��օ���o��J��Y5d�1����֝Z��^��73He��:Id�|���8%�^c��6����5X==�nd+7��W@��j#�dL  �kj����K��1��U������$A�>��1PS�Yr�؀_i���9�>�prJ4��泴�,//����v񰳳������z��t{v���|��|������ �)�#S���/w��NǾ�;e�����.��O��ܱ��h��6�H����EiWVV�+�kڠ��5�6\�h�J�`��-��P
b���c`\ ���EaU�>������u20X�D&5������wوPߗ�n���E=�
�*'��PV&+��,��cy��5��$����oLr2^�p�c�SL����Cc9�4�d��\��"��Y�X-�`�`ݝ���e��5�`�\��)FN^�秧4��Nk��I���)c��8f�{�wN��gS�f_�.��t&_k6Z]���k����}�~5��I�5��o��x�}�6���*�����~>my���	�	�����w��
zL��v�u��Ju��2M��} ,�!��<1�p�$W�lI<~.ݦ�u��᡾N�E��7Z����r{t���:��-jC�������3���x�$��F9��ݱ�2-H{�)|&����'�_Q�]�铰�"}�����"ʐ6�L�7��ͬ p�/��JA(2��([�;N8����KX�Z�͟�����R��`ik������ Z#�US�-e��s��L�u�O'�y=9��uy��od�!�t�C���'�6�5���W�?9���{�T�=)$J�z(tl>S�D��l�*��,?���%�h���w���9D���kW��/N�SW��&v��O1=�T[���}%�X��됦tFJ��	��*���e��Q����q8��ǒ��K��J��J3J[�`xP�����Pv-޲�+��1"=�h��۫o1�+��8����M��,!:�T�FdF�R�fZ� ����$���$�|����/)�gg ��3�$h�Ç��C|s\s}�DT[^�][KO��A�XWT��<��S�VZ��L��RfI��@E
�_���~�|�i�8�h<��?M�Rڵ��t!����X�;����}��Z��՘��-!%��N��62�\�]d�Ĉ2��b������uUlˮ�;��9�����`����=a�=Q c��a2�Է��2�|��$k~�մE����cKH���b�0lm����r���v��֡iCr���`+��+�p1���n��}[�18�٫��x5�#���g}O�����@��8h2���K�{��*@Z7PҒ-���g^%_lL7�R8U��P��ɩZ�SUUY���T��·�bnh��� �1��1���j������~t�t����������s��9���`n��ݮ_�9�O,�0_�([%��@�etϤU���G9��'0T�d���x x·
�TY��Q'��ke#VZ_�D:4����p�	K�	Jj�ߪB��4��=6C�xd�糖��ҵ��S�Q|*:������"��EäЌ�w1gG��h<pB��'�d���5�|Q���� ��f<c5B��٥���Y�ӟ䇎�6�Y�Rя�G\w�H7D1��jԌ>�=f8X/�ɫ)�H`h���W��4p��^<����3��>�4��'$�X�
�I�=�����!�a�~��prj8��m�]	B�'�_/�WY��A�5�X���k�Zj�R�|�p�x���<q�_vxf�l����T��Ṣ.o�awu���dֽ��؀��
P���H���0���7�Ќs�af�Awb�"�W�F�!�_�TX�;�����Q��ܴ���T@��l�c��8o���
&4#T��k�''��^�k"R����v��o�5��K����=O�m˸�[f[Ĉk��waC� �^u��<�4dK̐ҁ�a��K��V�A�d�YҐ �f��zE�a��w_���(%U�a/SS:9P}σ5�t���B_7�a���S`��oi��a����v�íF�`�=��L�98U�����j8������(UO���`F����ܔ�����6����^ƙ��?�O���pd*�v�V���-	W����Q�<'����S`�k�Eg�#�S)��vy
a����d*��P�[��;YJ��h��������"`&&�-���$�$�����ʬ/�����)���@˔8���r�߸uP~�6sfۢi����E+`)�9�@EUB�)������EA��2�ؠ3t��\'�+
;4K����^�Q+@��Rp&U8Y�{��g����P�N���D�����[N� �5��`��S),�p��6�ݾ��R�nB㤲�e!*@�e^5P�t�ImE���k�VU�P��b?��Ĕ�pK�����Pp22�-_]��s�Pv�}H�������i��j��f�<o��3�>w�G|�V�[�Tz�Ζ����/r�X�hi�-䶁�s�OY�Q3�H�!p�vd�KN�Eh,J:K���p�*�E���e@�+�5��'z��I���Ԝ"Y�:�H~�?�$��G\���Jٶ�k�i�81�i�Cl�눞%g!��b3���\�Y��8��'!i�a��f^ϗeh�u`�d�b��إ8I���&:�F���i7��S����G���ΦضI�=Cӌ
�o"[���P��{b��KF��tu4?����5I��V3I�B$��J�[�m�ʒ/a���Q]��g���Uw|��k�_lk����<��[J X��VؖV�Մ�/�)~]�6~�r�Ҥ���)$R�V)�*�5K)�~[pj���T[CdK��Q�����gE���:����38��N�����A�8�@��������M�ӛ7�$��~�*�X ��K����*�=��� ��`=�%V}����/�˅��k�d����X��!�Z}1cHn}BzuN �]-?���߫�Ny�4�́���'��s��
h����хS
Q�Ar�������a��%����D�'Z�$wX��D���%l��kRk�Ă�5���˧�DJ��<Y[��=�tqi%Y*-f�t�Sǳ�L���vz�+��8{��jb{����|2�W=v�@�� .��~-��YZ�|%����*�{-.Gz��j@��~4�^�xQ�_aid��^�cZh�yνz�m�R��W(_���P��ED\S�aeZf"�$��ؘ����jtj�M�D)�]�_�_k��Ӻ5G��U�9��X�q.�6�",�m�9��RG5s@V���,	-��{OǦ����JT�ɰ�qX[�@˂9)7e�u��=��/��Ф���<�+f�e��D��b��7��1z#�8�P��/a��;�f����-��B��zx�-�*��/�K��2K�HG�UI���S�oG��	дb�v�ܿ�߭�\.��4���Ԓ�u��	V�!_Ju����/���T�P�%�ח�m�Ejp�?�	%2&��=�����,�T+�eN��Ѱ��15s�%��$��u��k��6��qgR���dS�͉-\�8��_֫M�3�{/a���؃{įc� ��Z��bu�)�z��������pΎ4R	ڲ8E����{R�T���Fn��RJ�!Frѷ���ّ>�^se�_��`���(�C�.�,�H�j�Q��收-��(��l�#zR���W]���H�$��b���rw �ًb`d+��{v9���\x��%7 �;�MD�GTt���<��1c��V'2 <��[���^�~}��>���	�.}�B�t`�I={dh�����5ur�I�y?��xh��E�{N��� �׃�Amwc2L|W���~\O���]�u͞���>�[��1++m˃t",}��ɭJKu�Q�c��`�~��� ��e M�'�1޿��9B�Beh2uT(ED��D�M��]��5)�%F�E��PT�(M�V)��y6]2Cq��Y/C6|�!U�Q��D�R����$�`
ˀ#L�\t���u
P
ռ$�<ꆈ&� ����0r�:�&G�Ƚ�GAu�=lx���:m�&��F��;�ɜ���?���h���F���QO(�UӉ��T�3�2N����l�A���E�A��r��E�/������Fj�N�!�G#��(�mlU&,<�����e|A��ΡSmPm����CCCc��k�N��-n��6���mmo:�)j�(@��b���8��;�x,���T��.
*?����X��8�Ɉ�f�y|tI�ԝ�@bx��a��0W�w JDy�RS�U�)�:TVZ,7*�����GSKk���hB����o�e�xl���h�Z
���������&^r��*��(���J3��1`�s��3��2bG�6~k��O�L/�N�����WǑ���(�%�s�ah�Y���X����ɡ[BI-�s�#)C��p�`Ӵ`��U~��1!�#E�Fo����7���:���N{6/}�6�,��_��A�x�]��? �e�#wT�S��~��]J�[0��Y&@ń��r��1�HUX�y��t�-ں�4	K4��B��I,v�@?l#v�[��ɧ�vo���c���/	���ߛ]�|���ˎܿ�$<]��+��oZY�|���`��`��w��I1���V�X�a~Dff�X�	h�qUd~ۏh�n����nZ"�n��p���S2Z7��!(YR:	h`�"��QM����w0��B^m�6��0�������C S���@��,g��)��߂R�p�Aj����	I��bn��E��#M�D��8�a���.�'y���o}�lS�����\M��G6��ӑJN(<�js?�-,rW�]t]7q���Hk�:*��%
��G£��x��F*\$���Қ����ҍF�=?$�%a��K��&�S�K����ó�b{�Eb��{M?�d�?*��Ȱ�[���J]��Q�-c��)���6�!C>����_d��)�s2%O|_�ȶ�6��>�W^���.����ɕ��
�?�::s�,h�f���	�_����;PɜQ�T������Vc�#�?d�
n��~q�Ҁ���>q'�9~xJ{����rI�V�1:�	�0��h��O���@���CQ�gOz�/h�g&v���(��6*_�����k���G���
;D<��Y`%�a�uԟ�$~��$�,N�m%�(7Ty9����cd��6욹�.��� ��{�3Y�zA�Sm)�'+l�R��A��Ca;D{#�\��v���v�n�����9��E;t�y3N�s>irtXe��
!��`��O����ڤ�n���ͬk׌{�������B��jǗ �q���d�~��molm���n򬹆n0�*cbrFr�1��ت�#?��"*��N�� 
��g�ڴ�x͸0m���~IHt��tm����;�Ѕ����&���-L�	��r
#�V�c�T�$�ަ'ٜ���Yl���L�¨F/Ɗ��E	�i�pՀ�W������p��U�-�`�	��f����;�5l)��Z	:$�mߣ�ʚ�n��⤠MeA��� �O����'x��|_y0ㆶ?�"��_�X�g��L���v~/F�بC�&NS;c\��M�ѡ��nM]���~*?e�YfA[i
���TUty/,p2��L̿U,Z&��Q7�L�i�y�v/w{�U(�yn׏bSr>~M6��0v�Oύ�ٹym��|���P�R�m�e;q^�n�xk��##��CZ��!U�̏�d��ym�VbD�Ǌn��Y�@�f�[y!��+�A�Y�(��K�O�Y6V��:\����^�4������b��1�7&T���� �a�kb��a�  �C�������5c!��Q5��6�Z�KUG���2n�J������H��wd���KK�[Q��K��\���IB����
�MYW��];`H���N��VٌnW�F�ϴ�jG)�M
��o�.�z���Q�E�ɿ��NN-rO����.X�36��xx�l�tc4�+� Mz�*�Ң��P.�2���Cf]pg�*@��^][+CGk�5��)מGi5_���7������D��#����|^O��K�˾:t���I�2�h^�\H B��5�e;�ec8�j��;)�%�o��0(=R]�p�~W*JJ��;�a�
*�)LX�f��6�KQ�̡�ё&�3������,�&Ҟh�.?q�6�'W�-Lh�:W���b�^=��&�eJ�=�whu�^�4F�m���+�=���P���Ē�x�;=�MN#�~{���s�K_�� �p��S�������ë�]#it��W�z#'�0�z�y�hƯa�K�Q������B̒UU��12�߉.+��tG�Q��\Jk����O]o�8�	��hb<�~�-��9`�n�����}\_U,��uww��Lg��%�O��;�\��R���9k_w�5��.>�?���r��M;�(�e?skԗ���ojU���-?
[����A�����V`Ð̫&b/��ㆂ��� �y��r�x���������D�,ws�0�[-:�#�E���+���~�m���W̲����%�����9+٧yYjh���%\�r7�=Gu(1�1v |����}���|���͌��M +8�h�a:�d ����\�8H�a�d#�W�c��:��u괁����G�y��������`���$���Ѹ�I�jx�X �{9E�_�*�#��V�ͧ99?T�:�0C���ST^�a��@�����l�aBK$5���f�T���c�*��n�jP~��������>mJN���)��M����kX���g�c�$�K�c��"k"\����PT��%�M�8@�����J�LH��]�w d����S�������h422"3q�@*�]������X2
B����K��I�R� ?�7awь,<.n �D�>KbuM�F>t��X�����i6N5���3,�˧���HZ�o��ח��DT��ģ�?Vn\�ɷ�x���!*_�е��X���bn���ϥ�9���Ji� 7tK�����yJZ�]pJp�[V�ײ΄�Ūi��m�v�sۋ��}@�[.�t֢��Bp-y ���%�i'�����&�
�l۵���L��"b�0ǲ���H�2s��譯�~̥��=>���l86'�~�B�֒Y��~�Ty�����Q��[�iI8�!��><L9����Zn���Zq~ni�AO\���"�&����_4�6r9�i��0�u.e�,5wj�����^���+,� �����b%�O�Q@�-2"C�?Ѵ�%�"��d�UӔ�亃����ְ&��<1���G]?���}��sY-e���Cph��)��4�`�7�3��5��D-MHl�e3��b^�B�&�?nW�:d�c�Nð�A� #�F�1�yqj�3=\����2qF��T���Ƣ`���rXcRWQ
�o����M�u�����Z�����h���U�n���TZ�Q�2BD��>+G��|m Ԩ2θ�������Pj�`�e8�>�B����/�
l�4�:��w�(2j�M�!>|S`:i��65-Qu]MLF���ٿX�?Z>��y?͑��j���<b3��Ryt7/�/wFZ���NW%Dm��P9dk�\���AմԘ(�35�K����D6� �_������ �Ta�qa�E3�0y��zX�+��MC���A��2��Sdmr-�3.�����V��ˈ�F�4�˸���NS6$qL6���b ��2��z3c�'�zq6����w�|Y��)z���6 �#��TeI0$͘�S	d���V+�G�������7<k+d�	�.r{&��ύ}u<�MJ�e����ً��4J��40��n��b�,�O'w�Z�u"�Q�k��e"�Y�C�Q�LQ���*�����'��b�sԇ���u!2�8 ��֚��GE�Y�A[�-���<��%��^�-���5%�,�u��8�:������T�|I�����]=&<�9��.�t�x���E����/�d����tY���y7(�y�|H:z�;��0��Q����8�������0�ziJ#��X?�&����T58vR �u���kI=�7��8�V�9��m��Fpx�i(��Ê��k)~yZywB�A�[�K ����u9]�8��ĵ9�Q**ŀ����+$��Gmŷ��a��ʮ�zq��^5�@��� �M&h��-�'�ڐ渰gB
�9��F|D+#S�`�x�u���h\��!�����۽�G�}���
�l��G�B�d�T��_�J`ÉG!���s�'b�v���2��jR�.4jCA�1F�Fǥ�l�˹��˻�?�O���R�k���ڸ|� ��B%F��d(���?�.]K\�V������F���-+@����3Ӓz>��?�|F�+n׵_��5T~h��AiH4��k �#�~�p�Y��v+GWF���`����E[�����	LJ?/�b�*[\S�(e.'�W��N�����n@�(9e���ȇ��ɟ�ʹ38�S>������>�4�`����Y��3v3�X�|`1
]����J&S 0U�W�A����T����D]�^v��M?'e�!:]G�{���u%BE��c�7.	�liF��+bw�i�x��a%�ǶH���7ɩU�8u�.N��P�G�	/�ʴk˜G=QZ�D��N�})$H�ڍ�O`���l�z���o���w� l��3�Sݢ����rMG��󷦯^=>b��Z%��7$��2oY���ǋ����!��[����2���(�Č��D�3���k�������w)�KO7��oe�M�z�ș���p ��>�
8�q`#8M��1V-�ؑ���kw52��`�Q ��i�!9����X�2���h�:2,��o6�C~,���jF˼�x�W�'q���������+L�e��u��C@TvG�E�캹�¦d�Å��2&�c��)�'�	(C����@�B0�s�fc+�F�]
`q��#h�	�tQz�H�cQ�oz~��G�u@�5rs
�7�����F8� ��޺x`Q��	Q�6&�����A(x�Q�"TV���t�? W	��y����P�������	���co��b�xϬ��8���-1� +YBڳ����:%��7h�&#��KI9
�����,�:�r*��X���~�U55���|=��?�PQ�5oT��a*��,tS�^O�*_z�NU��[[D5���ڄ���]"�����O����_as�!�\�8����Q���,��z���k���gM#��[�G8Ð��,�rP�J8�k{��&�&՜?܎����7O�c��&Z���/�Xӽ�	OE�5�xg��KB���+6Ȫ$sg<�Fǌ,�a�7B&68�|j��?؜�0�m�+���5��o�\�h8��\��h��rR�ZF�aE
�e���i��&tg0pF"���e���X��.{?,�ՖOߜx1�P{b�Rj�ⶉ���<U=�<�F9���ʵ��C�1g汄9��C���!�f2���������.��3�����ܘ�5�֡����b��|9������7��+	�K�K��ͬ� ��a�Mu?���`3��;��93��O��:����.:�T ���ό7[2@v�6g�I
����1�e�{v�'�����C�J ���4wi�/��m�A�t��U .��.@ѿ;P��W�RvG���Aw��j����L�[�)��P̆�Ǖ�}Sp��p	g��Aѝ��V����]���+7�3���N�J'��ܜL���r9�+(kO�vR%��_�J�c��˱���,�G�#��+x�CJq�^�edT4u���;J
v8��3�:b'�4�BD�L$��V��"m@�#��3��ೂq�µ�1@`i#�X��&�dn�,gkԂb:ud%�f�I��8�'� &"��$���������K`�\�е#�W��N��,����c�n�'���1�pB�Xa�đ�vv:��ͥ��'�d�Jl�,P檵�c�������~ٿr�S'N<��r�GI@�AM�����}���}�����q���HAk��@�fuuMݼ�@`��x���/��6Ѫ�&nHo/]����=��k�U	����Z.�T�Y���Z@xL�܀p���DV�p��� %�&�/���r�X`P����3�J���� �b?b�d%��i��<���1�f��
��Nʰ���hX�p�o/)�A��g��n�E&1R�I����#tvQ�"p�a�Ę���I%n9��SѶ������bʺ���{��.@�X4�+y#UH�e�-KI�x?=�AZ��C�t(N� }`�~5??O��ׯ���e���ޝ�;

\�B�ײ��( ���E"�H;m)��אkH�l������c��G���i��4�<����)�h�j
eε�彡E%��u�s�օ�/�1�Y���;�B���0>QCe������+�z���n���{?��r��%��P >˷ο����{?���^�y(oR=�ur�!޳���U��0���F�ǌ�@��P�$��ܑ��v������c��Ebg�&�}WI'P�v��fuE
 ���av]D+c��Xa��k��'#��ɬ,W��%V�z5
P$A� ��%�~��NJ�Q!�� JP�8���i�W+J�ju{��W�Hi^�y� 
��^Ŋ:t��p͸�Z����k�������C�eS�1� ���J�(^��R��~L7�Z|D��M<yR`qy�}����ONN�V��q��I�i5���S3sS*ЖH`*FH�,ZPB���z�n6����?S	���/e��������������v��Qja��C�`�W	���iZh��	MU
^�0�A�Bq]��T�v��V����Y!ٰ��
�]1+��)Ԥ3���qB����:u�(!���nG[�37�y��� W)�^����Z�v����c
��8��`�qP�}r�"p6v�}���n/�$�151Y�2Bp��ǌJ���,-Ծ���z��������'��~I��ʩS/?�ګ���^�l���Ҕf����T˫�ݳ�����YW�P2��6L�r�L�r�
i@���	�;�!�oZ����H[1GJ��@�mt☢����F�M�E�#�o�)QsU�Γ�\���Gp����d]�R#%�����r���:r���k7�ŋեK���;IҌ�R�J�����rj�`~���Is�|'�G��� RV�˦����Ib�U�k����'�*ɬ/�l��h4Եk��{����ŗUI_��4pa�3�=���Z�XWs�s��۩��*�1 h/--�ٳG_�����?H��c.\�*����_�<��1B�T��1��hr���,t<�����f}r]����/��F[����5��R�+4�l?�+؁�릱T�/
1���]ؖ�@�.G��v�%��A�ot�5���M 67?Ms41Y��%���5�����N����'6/��gN.�\~l��ǔ����~�W_�����G���!d������b�jM�r�,�0@���8�����=y$Nÿa�2b-x��OL�2f�1 yXu:n�Ӫ�?�
�*�=C��:Fg�놗�֬\jc�t���#�}�U����c��q<�ӗ��Om�F 1;;K��+�?|Z�={^]~�*��0hCW�8q�\W�p�o ����tl�~�i����2ө�>Y,T�δ7���4aj8�6]�%��#7�z�S�Oj}�.LD �T�{Kі��R�p�j�*���$m���:}�c!�xm�̓��9�z�*kK�<aF����7�]��Gc֋���M�x�!��gj���G�F�>M����p0��}o��	!sE�ĥf@�{Y��^{�q�)L�����U�����lߦ}���!�Pq� �� č$%�p�!4�S���4���`���|��y��+�w�U��+_xb�ҥ����߳�r��$�C���j��=���W���0?�o�}cQ�����"�h�x�%G��v�Il��.2stO��@��ZW���:lydl�ϲXY?���iqP� �Κc𱁎�K�%��+U(?ym��5�616�J�K$
�:�^9�N��
ojj�mP��K�.�jn�󯾦�~��7���\R�L짹8~�8�J%T�8E�������mlf�(XZ=;*]!���)u�6豶#�/��f�?��#|.]9�=X9�2.��$én�cYРT֩�� �*�E���u�y��+V��;��uV��b;Ŋz�Ghb��8��bB������M��dB+e(`���8�r;��Q�������f�$�?)���~?�S 0q���MʠK���hI'!�`���O�.�h��ϭ��:������DU!��� �����턶Z����S��2S�2��U�9^�o�/�N=5x��g�x�{>��Џ!9 ��,�W_=���k��O�D��W��p�b�����Uu��-�A�h���F�V�+0��a�ZY Ÿ���$>b���y��Ti��'U�y	�@u�<.�#�y��V�e�T�Ӥ��{ª�{�WD��z��y:����u�1¥H�yr�Ū�W�����	|�x����ՕkW�]t{q�����}�^�yC,�������~�����y���a��~�qLLͤ�m��P��v��*}|W�!�
Z��u�$K����"�T�
-�$We������� =��<�{��������z�he�s4�c�6wZ4��v���zS��EZW��l7Z�6�nK9u�\tX �������ӾeNh~�����t�J��:v�	�{���y^'�T���ky[�9^ı&��ڲ�1Ca��L@s�cS��5�@���-NC���svS@S���G	�-IF�w2�|��|L<	��7�*I-  ��[�� �}ɂ��Was:��C�T?J�젞���wBmP��8��߼u�ߴۭ+��ۉ�V�����? �����_~��+׮�.�nZ��U�8)Q�T7o,����q#����+���k����Z1�IV�E�$*qI>6�v��9=T1�7%��/�U�ޝ�#�d�bT��@�-��<$�e�S�t�`�ۀ5E�U7���իjs}#����Ӧ�3z�8�.�Y�ׯ_U�Ν���may����cF�����qB���)�,&�)yS�L�L����0>	�]J��v�A�"�,>�X��P�ߨT���A�?bU	���*"@(�갂��U��4h�s{�S&[h�B����A�kKX�d��Uy�Մ�N��!�s�=����+��g֪\LW.PaN������5�3(��ӳ�'v���y)r�vZ�p��m��9J���L�J .0hd��?2ߙ54�&<I�s���9Z�۶v$!V@�bYu:�NVq�-��)�%u�O����J������9�|!֪��Z�ۿ����������7�s^I�����~�z�{�z�⥋�W��~���s �J�XmZ1�b}��m��Ŋ���=�hcr���3C�j���&���, PY�
5�𐛘YVFG�$B�H̫L�$ +Cj@4V��gk&1�S���Z�Ea
P��Y��� ��{zfR>rP��;�Jzu����e59>A����Ŀ���w𐪕k�:��~��+���Ϫ7n�<`�� >x�)�cG�y e��U'#����N�����4�uIa@@WmooҸ1�pau��H��zvkjvU�����J:��1�а�'y�Lù�('.��(.�#{ޤ�TK�	z�'i���2��3I�I��X�FV�M� �|��nlQ�����V�:y�� xY	� %�`?�/����W�\S�Oޭ�H ��X,N���w� "����S+���nQ�G�{��ʰ߀(Il�KףO���X�Jc@Ȩ|�=�F�9	��G�4I\�Z���(/�礟Y��{�qm@��E�;9����V�yE�js���q�@j~~N���(^X`�����{p�����ƍW�$o���K@o p�]���C׮^�]}�~�z�A<���R�ysA?n���-ʭ�B�d+4_���4k/�� `��]mD"i~����3���I���2�iljt�i�� �L*1�l/ao���C�\,��12IzERP��䓇2��D�ӎZY\RgϞU�����R����cSj�𤚛�W�z׻h�XaGԚ+l�W�v)������
7"b(U�b�ɸ%/H��[�� ��m���r���2��d1�Y�6|��Vbv��[�ldT�Y���Xh�u���d/�T^A[!�*�����ª��4ԁ}�i��j�k X��D���d�K|��/Lϥ�����5�3�v/B\��Kc�4?�O��d�+���C��o8"��I�uAe� S�|.L�����[�����RK��du��>�0-b��/<�u,5��(f�-7?�ҞLtߦ��a�"�+����6�����HU�E�n1�;-��p��׿�ͯm\���_�ɪo,9 ����v����\��������_@6�����_�Il�nw�W�qJ���iV�L�ri$�C��9�x7���k�a��,|��mF�8O�=}C�b��o2��8#1�ld҇�Aֻ��nb�W�V� ����`<^�f������^��M�E�]߄�3�jf�N��Z�&���R���:�����uR��D 1
���V���N���Z����n4)n���{�� /�)�K�72#�e����D��$�!7��+^e* �IVע�mZ�*x\o�(�~���(L��XAn���04`-�t�Ѣ��!�b-	w-���x��dR<N�<I�'Tl��cY�:YT��6+����@n?X��^��y���Z��Ǿ<j��7��N]�U���@J�#�ZC{Ջ�Xa%�����!�d	����.����֧����Hv{g����Q�P�[��
�i܋����z\'e��8�MN�~V}��5T˫k��{���q:G���#Z��1����VW���g�99�wW�Sr �$I._x���W�]�?����� .jj�-��F[�"5��o7UW߰����=!R@b:�E(�i�-�	�@�JmX��s���4��)]q7y��~']=�V�c�����v�:�T-���պ���Z���cI[2�h���Z��L`��-���G9y���B��9=������f<w����RP� ��ɉTq���7	b۱.�emk�f�����^H�{G���� ��@����<쮞x-�g:- ����ju�9 ^#�Ubr��m�ݢ1�w g8 0B/#jI`*+ 4x1�VbCS��,y4r͹����㒜.�;�to�����o���>������  ��]���K-�@Utg��z� �g���$)���Q^��$�Z,V��ɵ!��	aq������q�_����k@��p�cqU*����Bh�9Bdp&�l�gia�����?�lmm}O/�*�Tr ��G?Z8��K��7}q~b��s�nd�`�i%�'�ەk7)���jB��0z8��1�s*���\���A'�b!�FϚ˹�{.��:q�zsbS��������qS`��*��:��"p��̓\"S�Z���,w�,.,���������QY��Y��JL�'%��>��C���Uo���G���ߟő�O�x��gg��jrQ��=��IzE�������"Ӳ@?�v����ٹJ�R\�X���Ю���(N��E߉8��V��*���PYR0w�UzQ���k�T4,�b�T����H�9XP���Lv�r3����y�a�Yk	�����l9���"��5)	;[k�ԝ( ���#fF�x��14>�}��XCj9�1E�U��	ɠ��t����#:��a�h��\�NCl��.ʹ2�6��j�k��#�G��a#�]�V�wV�!�U,�cF�=v�*Shְ�ܐ��(�\�\�/kI.��F�����|?*�ʤ��8� ���l��z���EO>�������{�~B"9 )��[����W��}�B+ݣ�h�*�cc�4�nC���b��~F���Z+&(r�,<w��A�,��H�6��AV� #�N��Ȏ��j��)s�I9
���2��vd��Ε�����#.p��1}L5��
H{
�Vʈ�p���^�������QO?�4�P��P�p�a��b_:�`���:�>��X0����B)&�"��,���2�f�NމJ�d��wΓ�sB$��x��J�)8����6�̅��Ѻ���p�<$�S%YEl�O�3���$&�Dj�������뵵u���4�(���rH�:ǧ�\K��XppO��9�Έ���wj��6V���'TA��'�RX��}^ E�$�&�cڵ]y�-��Ԕ�q��Eb�M1۬�vz/���b�ڋ,��.� o�$&1��2-�Ě���iy&s���Ҏ��m�9�L�%��Y��G.\x�?NMM������߿��r�r�������Z+��U߾�e]+G�ûze����n�X$�p�;�ZnC!�<w/�jP�n�`�u!���R,{,-�_0�=���g�ʂ�#XG	MQ�9����>Ҫ�Cv����3[T��妠XHsd T�
'wBq��3G�33��\C�0�3ʪ"��r���������}��|�2�mB[T �zc��de�E<�d�@��e�m�(Q�U� "�Ƽ��2���v�$M�lj���'��d��Yq�I�TqW�+i#Y ���^:ҦA�v��Ȍeeb���p1�ae��9���5���` y&�T�wضăF����U�XM�\Q[;M��e��0ԋ	8�HF���N>���)�SlL�ՠG�d	t	��2�vA���%�<r#�Mb����gU�3�@B._��RY_)X��\Z�^-�N�h�x�";d%\���/x�'"+ �p��5��r�^��-���}'�������6u�����_��п�}���z?Ye�w�����������S����S��O�~� ��� ����ŅU���N1.��yT�Ӕ�G��p��:�.�\�B���B/�Rt��#��5ˠh)��q�$Lz��j��~���, ������z��N�w"�s`�!r��XhEi��Ҋ�(F�m�D�@PV6�U�����.�`<B@L���:%.�J��xv�	��+�"�dL��W�QZ�h>��j�W6bXO#��2��Ed\v^NϬ��B��50}����`�[bK6= �3;;G�b��e�6�Q�SJ�=��b�	�#�5��'����m	ЃՖV�(�5x�� �����L8�I�Bο!�\"�`M��]|����$�U�ϸ����S��a�Z���`��j�rM��ջx2�����,`�>/�-JP;�0��x��(ăff���NnG"N�h�������V�\�����.�h �t���Ϝ�U�j�-���O_p%����Ɖ�z��ZY�P;�6SB�"�[B���=S�J��T��S�˔ڑJ���@إ ���Ҏ�������}�1���IؿNns�+c-!���^P`"a��6��L�I�$�7�+g���u�]B�L�|�%&?�]&�:��U�U�k��V��
��ps7܌;�6�pi��j,�����a2���\.��BL +ǰ���N�&�hK2�-+�̥�R��F��/�bX���@����ґ��<�Ă�X��#�Q�#7u���7q_	!@�J�Ȏ���0��������帎���$[��\�#���2�Kqg�B��1窉�������pye�@�^76Umb���l����V"b�.�J
���ia#�l�>��q>J�E��ܾWAr'Y�!��؍�1��8�^���whV(5sQ')�"I+&�IJ��&�qcM�r�T���X�!���B��9���Ӌ�ΐ��p!Eۂ���P; �u=�3n��:���>��o}���/����{��z�;��jo������ׯ��n��p�\��7���^��l�j
�QgᠾC�����(BR2Z9K�a�Q���
J�w=Dry$�#�ll���q�9&@J+H��ʨ�)�P���R�y��`��1\3Pʸ�{]�z)R�J���8��+	8�ʺ~Jf�;Կm��*bAXE����ḻݶj4wH!��p(�C+|�X���+�I�8���@HV�-b��oh,*�Lv�ё8���2��Z�X�S6��2w�+7F����@����IK>�j��<�wx��(~̅��h�wz[Mr��s��}i��;���e+0��*,/�%_�}fv��Ax�֭���H���K�.�L�0�@Q�v`���'��H�x�> �P�>�|:I��s!D��a��r�(,�������1'c���q";��xL,QdA�zK(�b��0�
q�ۢ��R[	�ySQ�z�J
c�� ��_;���7����z��W�����ؒ=�H �R�{��ڽ���[� ~�$(o��8��t]�z�����#���f���W��at��Cyh$ �1"�++�	���I�׮(=��B`���o��A�L#�rJ�Q(��P��4�]���)�O>�-;��zC�l�i� 4��	���{�n�R��X���V�Mւ���f���ٗOէ*��7���MckS��6a�`{U�G6�����x\�^�W�q�U��ۍ:���@n��6ָЦ	�C�!x�� �Z0���0��h�߽��Iqq�Yk�6+kT;�J����RE�#̋b+_���vΏ�j�X8��n!sRB��Ƹ��w�mm+&�*@H���l��5B5.�X׵J���"�,����e�<F��`5"�D�����Օ��e��g踱���qC)gBD	q�e���D��\�!�����ޛ�hv�gb�.�R{u��M�"Ғ(S�<�%�ؚxd[�1���ؘ�3�d�_A��2��x��Ȇlk�vR�(��M6{�j�o���<�{�s��t 	 vS�(VW���r�w}�����3��@�����o�҅� ~݆=I�#[���j3�\�^Ĺ"��50_E�[���95�/�&i��Ǡ�34#cZ͗<Q��pŀ�D��W�Q9���]�f���{�]7*zv�C�5l�LG���Uȋ=�أlbGC����i�{�O������o�������#�<��,T}�)  �^y�[�\�r�_M&�_Y������9s�<�s�v��AN�8h�f���m�ȱ֧���xd-+ǟ��X��Be	���Y�O 7�a��~���� ��me���j��͒9 q>�`�8(% �p�Zǹ�ضַ�X��E����
�����<d�"F@���]��X���Lȩn���O���3$arǰjC�R�b���c��M�D��.�y~EI�r�{:��m���+�s(e"�[�t�5��	M���ãP���NFa:x���(d�F׎�E�w�A!��
伇� r� s`][(�
[{;gx>�u��݉h3���'?�3���Z�*	Z*`5(��nm hB:Jc��)z ���ע%�ļ�~TȆ���<G�ۈg9!DrO�꥜QW��qaE>��!yGs��}r� �qo4��1���Щ��vy݄k�]@M� x]YYu�ն������~f6���/�ŏ����کSO����S@o���'��������_�;�	4�Chks�!�f�7n��7��ĩv�"�� Gљd9�$��2NJ�P=�\(`�[��rCϥ��>��2�q�3)��(�sYB�B �L+^ A�A���0�,��s���w �G]��gϮ�������ս�W
E�/�!��n�ظ,��U焟%58�B�7pt��Z!$h4�fa�qH�ܟo���V�x��R�&��,bq��3��l��I9���|$�𷘋��x�X���| ptBŽ�t혞�c'Y/�٩���$�!�*z9)���
x�-���Pd/0$�	X�v�J$I��W8��y=@���i�z笓����X֡=H�8�r���Yc�7��6��k/����N�[ǎ�T਽��e�Y�c�H�B�mk�
�-g$�E��#��rki6������pkmZs"�b�h�m䟃ˆyM ���}�����|�[7��W���{�+���?~���}�޽{�^Z?�7Vq|<E��^�����$�0�A�:�A`���&�I��Z6�Qj�� ��C���z�.�d(+���pK�8�D��P9o\B��=!��k�����>C`x�U���2|�U���} ��ɪ+��AT�� ���}�jz�E��[�����I������+���^�g�$pPh��G�p����V>N����^�W�:x/����-�#�ץ#gЦ�����c]X����:>>�4/���5�с����H�3��pM��茿KY� �=�y�@���)(��Eĥ+"C�<*\o|�-c����H{)f�	.I��0����!/*�cQ��j�l%��cHQk�i��c%�p�3Yc��-0�r#��o�X�|k!�zI�6��R�S�a]����#O����{QV��m��xk^���{��ꫯ����?�{�鯵L�����{q�{�{闯\���eU?wx�? ����6�Jn�r��G~��?�p�f	���cYc8
�*���%(6S��������T�I�:Kʧ�i�P>!I��,�^UQ[x#+b�����&Pw��a��U�\�[am	a�B�E@��s�rem�b��{�+jܻ�kE��>-P� �P��
a���ZW!T4�l�܌z������ő#q_��5�mA�-){^7p�I���\E@�E��.Cf��.�����^�T��p��"Ͻ)\����8'�̷�wL�&n���1���[#<�8|}&���Fi8��)<h�E���7b^���($Gx��$!�;�`n(Ch��s��G�Б�&�/��At\��7R��	"�����pe/P!��=���-+Tή�ht�SƈJ�4���K��T�mA�s�_F
#�VN*�*X��4��JV-��頌�"Bh;]bE��a�m�P��<���]���S�2k�Bs��`U��Ǽ1��_��W���g�G������x_( p���⥏^�x��z�/�uX���������[�ٍ�Zm���4!�9v�z��|�%��|n��U�I�����s���߅�un�B!!���Ta)5��͌��½BԏX�60�~s�[x槟}����W��[�$��!M�nJ�~����c���;2<[�b���	�&z�y}��5��U��0D8L���� b'�w����F^�w��A~±rL#x�8JIx^��y�=�g'���*���+�г�< �Z)���������g�Y�#Qم����T���51�y���vG���[��A���h�ù�C��):�LU`�Z�
��_�E�YgJ�Q+H���+Vw���iA���K�$�,�F�W�����2F�V�­.�S��;��)E����9u��f
mܡ��yq�7fk� �<�{�1���X�~�"��+�u�{�����q��[o�/�~��{���˷�z��K0::��f��A�7�!��ޡ{�k���;:Ѻc��{GP.h�Ba�7��>��r�
L	2HḺ�R	���Zd#&M$]��J��[�ͬ5�@� �����������8/�<{�瀸��:�VcNC55�DB�A?R��vN�!��	i�����ի#=z�<-H@�1V&���zFc�w4�v���+ڎCy�ک
s e�($�Q�
�7�Y�ڐ�BC��Ă��4�r@H
��cKm��u�%�&���1��8���z8T��߃}@�d;y�}g��x��6�{��*2��=�b�1��+��u�ngk��tñÿQ��#� �ⴂ̚k��;��I`�|➨��u0ף�>;�NA��y�s"�ܶ����ɛg���h��p��I	[;n2
0��sr!l��z   ��9�A-Q��fC(g�ĕ�D�d���Vk�"���Z8ۃ1���5XkB�llځ_�Y_!}�<'��~�l�m�*M6Y/���D��M+�#�q��*	]���F���j�<�~��ӟ_�|���|��=����r��ǿ�տ��{���/�?::�9}���7���� O�C�˦�66�b̥֒���s�"�ڄ�Q�0\ �F�x�B+��=yI��q�[r��ɽܷ(ShI���!�r~cՠ��������_���yo�K���%h��ݾǞ@�� ,@	@0C���2ZL����3[��e����7����nİ�~�sz=\�ŇP���[x&\¶C�L�F�-	Q������I�@�����s���e�h+Y�s<��{{��ZrC�����qߟ���}q\�`�+x�4Hرsa���y�]��Oi]5a<�9��j�������޺s�ϧvB�)|�u� 0~��ɛ0#�_�p/#�t�bBZ�1_�;�I�f��4��f�)�E��؆!e�s�f��ء��UBе`Q�1��C/<�w���)�129��K���&?�b�=`Wĵ�g��om6�6z�~-l�u�ï����otݛ/�sS���߿|�k��_�B�������A����)�d����������`Aв�^
������t�rV�cElf	\�!�m1R
�q����s�?�ʀljC�8SL���;`�*��Q����b�s�&0���d+aC-Q�m ���� �h�F{8x?����.�e9���9Ҿxa���|Ƴ^+��7��'�+#�$�kЏ�49A�I0����@���(��'?�{b�$D�wx�����R
�m	r�y�B^	��p������|0����O((:<�SO=��BsfUc>����V�!O�{�{�R���|a	(�u����=��y�٬��9��5���Psl�~��Y�B!4s���-��'����v}}#&���j���g�����k)�P����W�2r2g2���	O�G|4b���Џ��Y3����i%��pвЈ�&�q@�q��Me�<�0�mO�a�d, ����y�(�{+k��6[O�^(ѡ��sI���w[�)��h>��P��U���'���@�>}�c�=��^�|�[���n�̿�t�=��C���B������Gn޺�/z����l��?��`�~�*CL���d�h`��5(�(ku˴�
�~���y�XZ������دg] v��sH�B�	ީv�@P(
K�2Q7��7��u�0� �QϤ|������"�����w^GgX�d�6e+�0�N,�e/�#r�ř�XK��V(4�J�,�y���=���k��~��<#�B\��k��1!������*�r��ׄw���������x�8��(���<(1y�8���<a��N�ݨ����&�����~l����q�Zd5�~����,�Q���
�e��j��"�n�\��F��\�@m}ɓIy��P�ŻP{9�c�Ke�J��`�7ַ��`�@��s^t��Uk,��6ۛ=3be���WN>K�'k�J�pR(�<c�4�@@:l<B�"yu4Z�f�z!����9���i*AS�e���~��N�/Ѻ�>��������.�o�>���>�
����?�g�_}�[7�P\
峱u�ݼs�]�q���Ãc7�͝zǀJ�N����TiPl��+�~H��
�հ��V��\AI�X�x���~�wy�H)#	<x���h[[�`�A^�b�+�����؟&BT�#"�$�ӣ�����0m����"06���o�#}���W��*;��B?/Ћx�p��E_���V� (S�^�j�+ H��O~�OJ��<+�=M�%��L������y%�%���g
wJ)#�V�P��-o����Ὗ3;�6�;9A���\4,dp ��?�{��2�F���h��'e�fkcm��(X+{wXބqW����&<˨@�NuG	A���[��v�������'�(�~��Ν͌�"s����B��Y(/��*�ȣ��o(4FT����B�
*��"��m
W�S�!��Q��2�<��¥p��?�4�M���A8?���<8�w�E����=��"P\A�L��z�:|�֝;��կ�͋�?yX{=�
護^}������/��Ş��m�W޹��].�yp�IV�Y�z����@�Id9���4�&tB�is�0%P7�qj,�z!�*`q�P(�
(u��'�q?0x[ӵ&%u3e(P�!��n����"�
�i��e����a�!��]�E@�B�A���G�y�@]�RME�����Ĵ��e0<�R a	��ŋ�U�y.�*66͂�����*����pZj���s��C\_��� ��g�9�R�7&����9��+��
{#�����*!����=\�|��fm��*sG�a|W@�$�j����y�� �J2b�!H�n=90��Č����A-W*�nI��ƺaﳼ��ub���C�ݟs���^FB�)ה��@�T�Rґ�4�k�=7�����ͣ)�:Mw�&R!�s���2 �
P�J��T��.���g�S&�
���P�}�Mn
�5���2� ���}A!<�k�,P�����������k������+�!<:�u7��������7~{��>������s�x�gw�ݸy�p��p�ŠWDa��l��nݫ��)��;U��YF��ݣ�g��E�K��-�D5��g	��G]8eU&�fޖ�yl�VT����y9�wU����A�� t+�2����Z"�+l�/jH�衂�/H)���f���>�0n( ( ��F��@D1DQX��EV��q E�j�wlbX�s.���i����XIuy/�>��H��g	BHc>>�����D�*�N)#|A��{Q�P�'tZ� ђ}?g#��@˂|�*���s��h@�.Z{���dL�w��s�J~C)�G��L�f��Y�LH����ޡ�Ͱ����E'P/kpp���!28�]c��X%�9�;DX���	V���G�A*eg��l�V��$M�q:xѐR*��yo
a��(Q���.�t��[�����C�b�U.�QR�A��um��c�T�J^&:4�|%<��B�m/O�E�V����a{���&ۙx><j��*�;]`n�3����o��_}�����>��w�Cv<T
�#�ۋz������" F��n������X�햕CE㽞��5���U�[���̢*��)mr�����G={T�WV�b�jV�J��~Ė�,C��k�����T��ryd�l�:^
A�%���[��0W,f!�  �o���2��&q��ALւMA,k�o(
GfY#����6���	X�W�_�.�b����*����y���4�����6�㈊���Rb8
�pp�� ZPMNJ�1�X���9�Z�o�ϴ��}�SƇ�������#�
�d('o�����2ޏ�P�8oss�mnl���{�����uPx~�*x�^�#d� й7�~Gm�Q��6��"�������>��Nm��ny��q��Rr�Bk���5��"���v���e�]#EU�Sm���̚+��)��k�x��������6BH�3�	^@�vq�ͳd?D\DƮ��ơ��<�����y�����ί���!:*��{��~�������b~������������^�\�Q^�g����2������0�ba7Qs
��n�[�g���A-u��*i<Q�ih�ՙ�Q�;	Y��`.�J)*�d�Kn?�����mWF�����$bJxLf�3�r?��Ll3� @��h96,zDU��qǣ{�C99��7��gm����ڔ��}8&�(J��L����EkZ����d������g��.�g�A��RH.�_���P��� �����t�����0�+ �v�y��u�|ט��ǹ�O��a�ƏX�5�hM��4e@v�����f����sp�O~A��k��!le!�6!+{%�rPD g̦��n��CF<�Bx����ʯ�V�x<i΀����<�)s%�=�4 �:�`�9R2�C��F�2��3��|��|"3 -�=�8il���i�J���p�66��HGa6����a�.�W	���6�I-9p��v��@�ye��H�<8�G�6�V|T�Rћs�z+@����~�+_���/P�����s������_����GM;� ��HH��O���.����q���c�(�l�]� `���(/�F�_&�A�a�JL�}s��}��M� �(G��]��q��5e�)_�\��_ڀ����E8 �un,?���B:��<� BDed���PRQu�3� �=E�ϼ=& ����6��D	�^�Y��r_�Z�\�r��Q*������o�9���Q�P�y��{饗<��B��-q{��`T�����ۧ>�)
D1(opt�)�o���Z`-�+�H���v���|�׶��M�5k^�"Q:�/���5�;>��L0dTCc��:�	�����ۻrM� $�X;f�;
�E�kS'C�#�+K��Aò�Z�1Nh�������'j�?'��������d��f8	S�����T[���?oRx�!�A�Q�=���ҝ�c�>��x?���!������P쌝^{���E��~���3��8�	�:Լ��^�� !W��F�|Qԁ��^���n˪�#4?hc�F7������_}�_<���n�GyhBq��U��ݿ}��_���a���#t��t�m�:�^����9pG��#8��dl�U���c}}-�2b���>F��$�\�tf��r+��s9�3�F���B��s�@��=���|�
���w)>lN,dX�=�ս��-4 �n�X�;맩0����1M�ոi3�ᨸ�I�FA�'&���L�9RI���l�M��Zh�N���Q�0*�+�1PV��P���]��uu8���W[-rh�ȳyT��Α&��ރjDh!��0_h�v��i��c��ԩ-Z�*��ф�㼩g��p#��cy��pT��{@!Ɔb^����Tԉ����:�*�#��<�X�Vݱ����[��)@��gէ��dX�֢�o�g������ĝ�9��:��l��s)� mf���:���ޢ��td����S�au-��V��ZpʹX7~n����\M��!���$@qb� �gn�	G#�)�"ۙ�;A	/�˪�e6�#���q>�A5U[#G;=��F�	a�a���b���P4;;��7���k*���e��}���W͜߭�tV�Y��8��7��׬]���9z1l�e�@*`5�ɹ�΂���k�[��T������/5�G$h%,��������[��9�T�T��눞<�e����x���xXX
t���\|��?;f�֏0����/,ݽ��nwϻ�c�<BU2Vj5�X�x677b�IdN��\��5�X�#�hc�ܪ�-���~Gh2uϐF� |X�-�!���-�����M,�A A����*s�ߐk�[pT.
!t�ńX�\a�y�S��j��=lV4�*Z�宅� T�0��f�D�\�̬�e�T��FB]!�����>	�r�����C�ji�{�9M����������'��ތ�C�}bQ�G��	���?���+�./�X��3;���iv#��rP=+�� �@��;W�1��(Zk���k��o��B�59x���3A�L�:�F��G�tm�\[�ằ�Q�Np�"� ���+�"*�Նu���.͇�	�K
��ЗȠ�<�s��%��e�U,�f��^��e=���f�]X�<�|=�����]�Z*+!H��#���a��+=(p=���7��m�2�f^M��P�	����*ೋ��=�."�)����;~/��2t�y�B�rOJ�����~���Lq�*�7�N'O_;<��|���{k���z{��_��kW������&u5$��ŷ.����O\�I�%X���A�(�߭�b-���EbR(���
��	���wr�MY��YU�=UU�E@�)DU�ϰv����s�+���O輨� ���; ��#Ӛ"��/Ȧ	� �EGU�+���C1`���A�����:!�4���Q��T@^�����	٧?��<x?���	��Fp�~�����ɠ�Tu_�V[ߜ��@P(:t6�B�A�2\����]�dE�j/�aש���ݸ6����G_RȪUR2�b`�$'~=��GFE��թ���f���dY7N�*�2�|��^�o�͉����w!wT�(n��q�f���M���L[��.�)����<��/

�7��� �P?���a�'#$ԅu�͹��rf�!��z��]�؍�H�>�L0g�r�62�oA�MI�����2��<�?w�{��14�R0?B��aƩ�� ��	�?�O��o����>�?�˽���V@����7��t����擏��l���&���wwݭ�w��ǐ�ь$K�Q"����=���'U�guE����MP�6ҁ���7t�)�^e=��-�0U��E�'�:wɚ��ƣ�H���h�e�F�f@k y5R�m#+/u������R��<O��6A5���5�nĄ,����q�ٺ�1�P�
=���Ql�����~��g	:�{"������AAA���F��[G^x)���k�?��v�� dŌM��qd�FN
���SOy/�����[�ϙ+�=�i�J�?�c�(#�\�F|v [@y�)�4��H���kyS>�)��7�`|a=�E�m��g���5K�y�~���f����8v*I|zڍyZxN�O�<��Ru]�:G�d�;kD��-��G4܂@�ΙW�q��=��6f#W-��l���v�I��2�_R&�8W{J(�6� ˰�O�P�|gt�m$Gl����>��S	�?9<Ҟ?����ϗ��/����;�@+ /dμ���ux��i?�g0y`@���x�.�}��}F� J��Z\����пs/�]u���;��#��"-�f(�^p����?52f>a>!�.*@�`MC�&*���U��E<�YPX!�#vc��f͏��^5����9x>S���*��A �^G,ˋP�ڡ�'4GS�E����p
���<�2xw++C�/r�`��A���,s��f�1(9|Ƅ��:��7� p _8��s�y�*tE��Eb������5�����]w��[\7�rSs/��@~�PԊ�ZY[e�!>��3��1n���N���/��>��/�x��F�zI���6x疭�r�^0W�$h~t�*�b,��D���}�u1�aP��O����G��ax��w�m�(��2��`����{zz/�l���A�Ϧq�����K�:���M�n�l^��l<�g�6��|����/�J�@@���f�����F����|�D
cx�������W!T6�25Ay� ֘*����
נ�$�G��,�^9������������wo}��_���T\�w>`������������]}�7��� ��|��cl{|��mo9����(p�e%H`�<VR>��ϕ��-�u�U�8�yNl ��*�d���藺W�0�LBrR�v^��f�U�P�b�r���ǄLAD!
��6��}K�IB�����jO����,���U�+Y�R�6��f]��R�،����?�^�uC	/
�>sƼ(�|px&�R�"��̈́w��G~
Jޕrj$z�������C��1G䒲�Z���r��a�t=(i(/xrPvPF�I�3�C�s�g�� �'t�u~~	Λ3P�wM(�m��2�dv���Ⰲ�T�"oǔ\�����jn �N�RkD{��\��<���܋��72�"�i����H�B|Z���HI��D+a��$iEyS��~#`�_��l��rD����������{������`��P�I�+J~�s[����B-0��h���sz;KzƲ(N������˿�̇_ j����*��h�����ߟϦ+�rmA�s�a�ݺu�+���XC~/�p�]B�d"|�4���تIX�H�j�7q��"�ac��t6I�<�w�R\ytOE'V����r��g�V��g�n�˭1��p��v&dS1^]��%�x"v��
tc�Q"��,�R6@Ah���0��9ۀ).�8�~�,�L��0�`�@�)�\A}�ӟ��	�7�����a�Z�;�hP�yU�4�I)Ձ��B.(.�p�R�l���0��sS��~�VB�8*�^�ց�����e���}̩�\.�U�)�ϩ�	�Tp
�����é����`�h�EO.�eh �o�ִ#��gUXCxGe���(
e�l@��Rul��B|s�Zb�a
�:�Λil-.�/�/��"�Ըmj=>'ƛu_���kw�@�A!𴍜�J��F(�7�oRd�i�x��2�i(� ��,vIa�۴��f���kj�=C��` 2O�?����1��2�ZMh�;��eJ��hI�{��=�^U���f�y�՗�ӛo����sfۆR\��η��W���ٳgv�c� @Μ9�N��굛no����E�W�Y�#���x���:�/T��r�m�Yd�hs���>��d1%u��b�QGv����`�\�U���=cNFт��'!�}
��B.R@-[bC������X��q����H�Ye)
!u�Ѹ>�wy�yN-k Ud�&���Q��"B��(xB��<��jSh�rR��U�г���	��e�:ˡ�T^����#�sA��9Eۣ�V�c���Y"�YP|B�Z@<	�'�U�i����+O&x_8Dv=u��ة���Cf��Bv>OȚK*Σ�k�<��S�B���F��Ca/���q�G�C�c
��L|�]^r�L��w�a����l��ܪ�~��bþ�B�P4j���$��0VP@|�ʔEb���D&O2�q-B�R��]�롃,B�E�		�r4��ë6�8k�o��o�so�����?��+����x<p
�Ol����/���k�+��f��r���x��y�:�栟G�E�]l�Z�Ql��C�䡟��D9(���Fm��I���Q���SN�ELd�+Y�!dĐ=.�K�e4��Ѐ����".z,R�֦SS<\�u
%�}#k���a�I)��OY��B;X��Ɉ�AzZы�a�C�Fw�`�� c����$٪�q��Y��9n:�
v:�~u-nb/R"�BoJ��P�v�'�]��!i�� ����a<GB[9�������_�UCDʅi���PB�T ����q�1/�����8��7�p}16h�p-��o[n�#\�ǖ�
��
R�\Z���t�( &�q��5��� �!�y�!�<,D�-��O��.���9t��>��g w^>��HR����أA�D��*C���9W3��r\�߬F��l�F�ת�5j򀎃�R�������Ya Sv(�M}��y�Bѻ�8�Aj���Q���dt�1B���hB�~y�Rf4���ޟ�LF��K_�������x{� 	��r���o^z��<:9��_ [/�Ta}轁����5/��<$F!�4��J-��:�*FlIs��O�G�G
9-�6)�"u����/X��E����uO�	���JX�f���4m^���!D��	�1��`�F��mB�c�aN6�)C����>h��R�@�Cc�pTBh[)�e/R��B�$R�a�Uč���}�w�KƂ�b�����2:��������T�UK��IA�F9���Q����/Y�8p�����)H苡]�1�o�Z�sh42σ��K�a��,��u��3��9���6���!*29��!���^����'����4�� l[���a�U�	���"b3���1z��"��|�qa���c�Du�xq��Ӻ�����\ʙ幹�����姍�������k���hoo�ZX�9EC%sk߰⍍gnܸ�;�7_z�A$<P
�뮬|�+/?{tt�����Qxy�ꇇ'tWa�[((�CF��[�U��za���[�sA���K\ZyB���=7�3H*�)��i��cq?sL��� (C��[��(u�M��1yE(�������0ʧ�ET�����3����9��Y:��׆�k�P �+�����/9�BVy�\�*<�[����Qw���s@(��B>oR�F�CBy
[�%��Mփ�JJ��s'RK#�\,��E\�t)�R�M|J��?q\C5E*Pe>/�������!�'a&/J�G��Liu���b�D޶2�����0~��o
B�0�T�aU�w�m���9h����.�����|�B�[T��z��M��QN�n0G/�C3�>_R���Y�l O�\$C�h8�i�+�g�Pj����uV�o���N���i�Ċ.,�k�+R�l�
~n���	���;ƾ���G�`� o�h;�ι"F[���Swowߏ�m������Ɨ�w�_�����7�W~� H����R@�.�}�6��>���h4u[���n�
ŁS
qK�	�R0�Ń0A.��"Y���u?�Hd^�����M�&�+)�$�e]�"�P��.��,yRp��i��Fc��!9���Z:�ڎE�H�
"kmXK8v��2�BG�#�8,����b	��{�����O^`b�V�+W`14O�)	cy2�yv8dm�j� �'�yE�!M�����uy�Fy�]��a��2!#��cV߄ހ��-l��h|5�o$m�r^d�j����5q�D�d
��aeͫ�֢�_�K`��ȏ�i�=�[Z�%� � ,>�݁4�;�51
�K�~7��@kG�C�e`[�0�U�h�p@Y�xun��|%�[��I\X��׼O[ļ��oyg���|�pn"�M�_�f����d�[����[�h͗��kz�`1g^mc��%�6F���{��W����ow���*��F�9�>?_��?���3'Ǉ�z��qP�0�����o���=���y���I��dȄ/6-\�x��]�>�a*�Q��}B4��N�RԦ�	ϔO|~guUՏ��װ��� ���X�W�`e5ZO�L�K� saW^d�.�a+w}r��5��Bj�C*aX�](J�a�5C�p���bs��_Y�Rd��x�;�=D���x�t�&sZ���WxG9�v�
��9r�<�"�rkI1��|�c�/�f�F�&uAŹ��1e﯍
�Rԗ��.G_�`��ji\$��@��e�홳ɠ����!�E �ND��q$�X~�}
B|���.̓A�Csg�f�64���ͬo� *0�.mC�rW���8�6&h���P4�[�XEb}�r4�*Ư��J�s��`� �Sh+2��dp�5uRR�ч^�u�-�2g��'l��L�Lh�VAy�~.�'�T/X�}�l���m�ń�uh(��Ϳ�Q�ų��JRSp�� ��-�8���Sn��f�g!������������}��.��x �_ ťK�=v��w~�m���{�m=����SN�p��q�Yhʥ?�htcs��?m��ѧ{�y4���c�$�����;.%R����k��r,^���J8T���hY�
�H�K@ͧ�x=	b,Z��1�f?�S��{:nN�ɸw�?Kp�>bo�ktKJF!
��"��K-�uH����u?R�P��.�~����'�(�ÔO�r��*B����Y���mM�z��$�6�>�B�J5Us
M�c�_���D��'�x�>Hd�ќ���ދ ���r�w�����6N]�,M��.�l�2���:2��B����U��X>�gq' M��������V\]$eH�f���v�|к�Z=����VNS�"���T����Ѹ��c�3�,����0�Ԕ5�"zx�jԞK����*��z[nЧ&w9�%_OѠ��B��s��""7'-Ɂ�NF6Y��+I�����-����|�o~cw��ݝ���x �իWO��/~~<:������M9�$؁�}�ndw���
�6��↥A�fT\Pe��X�@����N�.��]��-��,�z�+t�����\@�S/�?*ޓ�d���SEV5��^�Λ���0��� 
+(D�,JR��Gҽ{Y� �Z%X��>bR
�&*K����@��9G�n��X���6x �6�g$\du��2<���\������,se��/�=@��5�� L�j��9*\4
��&q��g��8� ��P�s�Z�'��v���SjM��b�K�9�[.a)�h�wua퉣̌�E� C�d��x�{H��y�HmMI�����ȡ8r�H�*�?��*s�T�#'��5�4υ9)���ۂ!��o�7<�uh��	z�2U�&~x�񸥲�3YM@ �X��:�j��G����:�o�9X���Hsm?���_��d˯�@;��#�$O쑀�d��s�s�He���������x����s?���/�3���q���n߽�_x9�d��*����᷻{��M`�v��#](��fneN�Se
���R�+O/!���\ ��Y����(�e*�t��
2}0s�B,ܕ���-8Y��) �5����d�!��#�b�x��P�v�����.Mى����L憄3y�Z2hǍ��S�́�LuSV$H��xRRq���Ƒ���(mX1�D�ٿ�׆L�|aت%�a�"��YH�$?�+��c�H�s�.���v������t��z�)2�s �z�l*�]DQ�$zz!�u�wzN�<��I�kM�9�.0q z�\���PC�"��.E���ޜ���`�ʉJ����(����i0��mT(<\�o�BpRB�����7H�f����Z`��� 9�<�x�M�ο�#3�
��<�F��kR�*�!�_��4B�M|���<PP�"��X�Cw��\&Ȩ2.��a�ya逮�vɋ����1jUmA@���!�vg�4C����U������+���O._�|�Ah��W@�����?��O~�x����.O�C^%}�`�.��V��e�"K�Ġ�s�{�z��a��+�
����VZ�W�'3�!�\*��Y̶�h
�&�{��� E�7�5s�Q�g�!�G6�}�6�~�YD������{A� 5����ȟ�+K�[Q爂���0X�+K\eS,���cZ��{��l��ܩ-4��\@�u-�JB�7�ψ��g@CQ��)؜α	�{N4#�~���pu���.�b�'f�i4:����	4��SP��,��L��,�у܂Y�ɐ�53��Á2��3��.9t�\��u����G�PyO��ƺ����O�/��~�S�r������iR>(a�M�9��'�����uV�������x̺��5�N��E��y�0��\�q=�ƨ1������ �ax�=��` 5���"�ѷ�Z4h�����|�#+���Ϭ�z�Tl5��J0�|����7`������c���ݾ���2N ڹ{ �m���Ҡ���f���!9���!��,�Ysw��s<Ú����o�U4|��G��T[�a�?1�-1��I�u��ag5VP�a�2��P�ZZg�X��Th!:�,� %v��_�C�e��P}e���w��H߅"�����ݼu��:g]{��������;wv���7/]��W��L�9� ����?�����?^4�� y�����߾�筶1-���E(�\�k����J/XC �\���+S57�Ճ#�3\��� ,��#B-\�Û �B�qZJ�m�)�7Ƃ�0Z�ޒ�DK��^@	�V��S&�o�A�\i?��̙) k�	�~�/w��E{��u�e�#���S��Y
ϣ��,9��]��ss}-z:�1w(y��P�E�tX��9�v���p_A[�Ɨ����M��ޢp���kT@���ϓa���~��x�u�NM?z����~�=����7�t���o~��������潠@y�	�5m�g;��_�Ia|!4Q��<��+�V����rm2m�'4��'~  �\�y��p�a�6�N�ޱ�!|[&k����Yy��=P�0f5Y
��!��5^��LX�8T3lȉ�)r�Z�`�a0p���E�0��"PrQ�T�>�|.r��fi�h�8c��-�I��1�u��{�]97�i)�5D2Pw�Ƕ�s@�)\Cɂ|��e�8�"+�>��M��qlnnl�ǣ�������ozE׽�����y���.}~:�|�(�M&a++JCB��Ћ&)m Ŕ%��[_���K�b�yWǤm^?��h�)!���	«�3T�[��IN��R�hX�@�K�f0O��~'�c/��PJ�L�W����Z��}��m�a��H�=�@��K����CP��n���B�[��[+��T�KHB�1,#����<M�S!���m��Ce&��6�a���M~<����}�{��^֊����._������C�	1��R��~޸�&�.gy�}�ӟr_�җ��}�y��sv�?�(��Ã=����r��ƄЯ*�#�	E.�A��)4̕��#�����~�̓0�q�/9���0r(^|��44nB悆�L�$/lk���=���'Ԩy. �T
�\�h�>	���ϛ��5�����:t�ĂWݵ�A=I�p??�~�������Ő���y�����Z$V�N�&m&������#�!n��[h(���Ӵ���=(&��T��έy_����VP�M}$+���q�� E���֪�����XT�-c�ߦ<���Ͻ��7�ڟ�3������o����~�m��$��V� �c̘�M� u�9c�2�Y,�sh�p TSv�ZK0��RwYB]�u^�	��]���[b��0��Tu#y͊Bf�v˯�g�Pm1'b=lN�`!'��\�ʅ+j	}��Cq��'�Y�|�Ԑ��Z��5E(k\��T�a�KHC�h��С���,W�RFy^���ݴm�q�U.��\��F��W_u��^�ͭ�9fW/�Cυ�M/��9�6�����I6r��/��;���/��e�{!urMm��dU7�dR���N'X�yi�k�w��a�2x08�f5&F���_r � (j�ז)������g_KHP�-L����V��prS`��w)c-�ή���K&zOS����LA��3+�Y�!��fc����zb5�_�97c�	��u۔q_�Ò!��1X>�i��"gM�p�I���7��B��&s���+�7\�l��1]����s;�+�}��e�{���/��7:�=��3��{�x�*�k�~���?���h��Ţ�tl\�m=�w��������>y�9�e�g�-BM.�6
%�����e���b�[FU�>��DdC�S�9*>l��Y�R��Jd�
5�m
M�B1f-\
�:������ٞ�+4h���N���+�D�=�	X�i��������j�T�1�@�`e�h{�a
��QG�(?
E���^�֑H (,�#���8�]�����e�T+�-�3�48eH�r��r�����g�z��������u��G|������Ez�Bu�ϟug����w.�S^�ܹu�Ȥ�=�Զ\ϫ�Y*���-�E/�	������;���X�C�/xZ�;�Ħx&�-ٟB�%ק��1,���9iܘ~=�
9��t�3�����[FB�BW A�
�1�,��������XI�6�Dk9Y�-�b� U���W���t���<iV�*�|�@�2��C˘�Ftbm��L
�8��?�q!xh���\�\�[���_ x(�8.Cn�Fl
�rf�{��C�mumōOTD
���q�`�m�Z��}���J�J{8\;s��_���������=ھ�=�����<����?Q�1f_�ҨI���u�{ǌ�"�VpP	��K�Y�V�ő�^�#G��7A})��
֭�Ң���B�T�Dϝ[DR��J � R�Y1[{ވ~��7,$�ݠ�R^��E�gh�p��nG�yH��j�K�FEak���Yֱ&$��E�<�?$_5�!!���b�T�Q��[�W�Нꩄ.�'6)>k�-k��?�
���{&����#�<��k��7�|��A��C��Cȥ�'G�������_��U��>�>��ϻC��\VS%�dȵ)Qd9�Ma9����OU3�.އ���Y���a}���{��
�q�O�sa �#C�{�%c��I����(��7����	�e�C? "��r�PT���!�Aa��gϿ�yʊ�gfD�P�Q��i�.�r�C/��W��̓T�_ݣyd��yc踜>�c^�Z�|x��j�e�ɏ-I2����������7��P���_ZHr��ᎎ[�bu��c�VWח��W��� y�W^�����������yO* ��7���?��_����eT=�ݻ��О;F�u��O��9��$j�$!8��V2�-���qe�d��EZ�8�n�wKp�==Czњ�3e�`�،3�.
P-v�&������A��J��f�p.��@�
��S^��g�ío��A���<��Fa`�}�>���A�l޽�4 %���&(����ڰ-|�����ܴ�e���& %�D@����b�X��j:s;ރY��u�.=�����poϽ��~��\�Zo_~Ǎ����_x�?{KӞ��!�ӧNi٬9zK�j/���E$��K��
á&�j� ���s,��[]Y���f��������z�Jf<��zD�U����K*��9���a�'(w��K˥	���Fާuc9��mM����N���I�;F�
1�g��0��BxX���Aj�����(�M6P��擿�tD�g��f���G���HL��\z�&���S�B-�+��}�4):bF�r_"��t���PMV�ʐ�nA#���XY1��@8��-��%�P��x<�2ٙNǟ�p��'�;�,ރD��It��KO{��s���Ċ������{��g�5��-��f�'��5���o&r�<�+�&$0��qEa���`�aq�(n�`�S�0�^EAJTR���h�&�#�WV��=�^e9��msm3zM8,�* �`�+� ��m|���<���A&x(4��-|֋�.x�e��[!�uw�孹�3P�oY�:Gϭ���p䖦ޝ�|�Y��(�0h�F�g0NPP8H�
Y�����o��f��	�A�,���
Ɔ���G���iB�/_~˭���u����P���u1hfǰ�"��јs]���<{�����#&�S+�%&��	�N��F������1��iCX���@#�h�X� #ڜ[;�as(`�6��X���G���R^hMϮK��x~5*�se�����Ph��54N���
�rgr>a��7
U�}6�ż!��'90���b�?��(ߩ��: ]#ϫ���,��+�ܙ�uu0T�����X��=�O�]!�`�l��y�K��ŋ��v��=���l���~�K��'�S��h�������@%Ӓ~�����1Q��Y_���ZQ�Zm}n��by��+*��	�����T>t���JN�7�|�鹉���?���܌��
,?YĄ������6��P>�x�tC�M��9�)���\R,�N��F�2� ����>��2p���
�d����m�
�.������0Z��J�("�����%�dU/Z��iJ k�B�C�&宿<G*?�'���^���x<%�ی9�?�lH��wۧ6����1wӏ?�`mc=*�<D�f!�#�,�.��4w
1EhrՏ��C5�<��*�E��hHx>�kxրX�]�l���bؒ5�z�0['��<��0�B����4�ԿI�>y�Z�C1�����WK��ğ7D)wb}��0��!�C^74���P����P5���C�2-BB��
ԍ������1/�d����^vQ��0
R>Z9�%����5��Ĩ����*��X� �3#r=�y�8���.[[��L,c͠q��O�u��7�~�O�����q��[�ܹu�^0�3[G"ē��7��g���u�q|��GL�j�͋tTJ"�ڂ�C��@���Y㦔�Q�������V|h�w˒�4�h2ޫyi��9���)�J��J����p�X@P<xo|GF�@�̡Q��Q�Q �N��Ue [ț�B���D�Y0��k� ��dXM�,	zZo}�T�Y��37������7	_�>$@rOPy5��'�TV.qr�`��T?%�}�kܠ�5�W��2q���p>�Ưhu�-����>�u�S!lZ��<GN_t?��,�<,��؄�2J%�ZD�`�8�m�8������dN����b�l�Q�~ȝ��{�V=������1$^A��O2��,I,�9��%"
�Z�s?���B���xY4����^v�G���-q��!dF��� ��7�5��sXOle^��	#Fϖ?k� �GW�4G|���k��K�戊��m3�ш8��Qfre�{����s��/_�|��{��=��vw/n}����~�?\���L'�w���g�
�Q��qS�ȷ���rPku��P���!��)'��>��$��,�P�`5F���0���Ef���Ժ�"�Yf��\��oT�A�W��3�d�ֲ�B�F�/%���wI@y �O*͋�������H7W�QY
�`Ⱦ�E���[��bm!!�N�9q�@\:4!t|x�jL�|��e%�$��������C@����?o2&��B�C
m|x>q<I_���3gܭ�7��i�1t�����D��V��f���x2'q$�K,����3��=�d��X�LAr����R�8rrKr��g��$�RQغ��TH:�Z����'x��nȢn����j����*��A���f@��tfL�B�S�3�������pĥ��`I�v?>nc��#[F�:��.���XN�7Q҉��}P�,�� ���5�Z�1%�����q���/f�J�W�hÚM��6>�JvA���v}��pѦZBy�]i�6��ZΜ,N����b��07��8��k�4��\����n�|q?S@�w��˷Oݽs�W��|�圍����6�a䫀:�)�}ۢ*9	ti�.V��8���UJx��fb
֚%D�F�.�_�o
 �����hP2﹓[GyHI�,Yya8�t�A� ��MyLQQt]�D�-�Z�Ux&�(��b<X���:�AJ�l|�o�9���H�f���Qp�q����ͅ,C��t|a�֖�Ҳ�Ś�C�*C����n��&�^�7v�y�'���^�w�С�d�z��g(�N��/`IX	븜�ՍM��uʽ��Ew����q���,��h�J�*L��֔�4�^�x:�;8�\q8rP<u�+rT���6�����Pg���֨����u"�F���p�h�,����y�&��\!�92��V�-B�����_�T�85߳�T_���	򂺐�W6�L�S^�tC�\&=�ʫ�5���w`��𢋜t���8_1���ދr�Ld�8$Ob̥�	�3̍P�e�v�c�Q�j��P�[^o>��o}�����ϝ;w��#�{Fuݛ�?��>[��玏�0`LzccS�G8�+E�r��J�CI�YgӬ�O6�8��;�P]���mV��]f�4NT�v%�L�C����_�\�@܂�Y9/�6t�k!�d�
)4�Ń��t�@�%�$�b������'��˘;@����+!�
I������R(	yX�ma���@2`ؠ��s���6u�đ{3�Wy;yL��S��F��<�+Ⱥ�0�:��^��k����"  @߿P`���Ϝv�?r�k�a���bKww�ј��Fh�N�9��
��{|25���Z������O%y e�ʓ��k�zM��ad��57J9[�[�Up�;^�ĵn���bJ|nm��錞���J`���n�6��e��ύ�}0�
y�Q����h͐������B�~k_�Gљ�^�P�7��LNF1Z���9��\�pͥ�Z�Fp<�D&�����-�L�����`���: B�n(&���Ay,cHI��\YR 	�-����]��6�{~H^T�Â�[��N�z�!�v�,�-,�Ct��v$�ս�u����޹z�7._~�;��?S@��/�w�^��������\	�/����	�����6s�e%���"!f&����La)�n��5���j�SU���r�G�!��O�	ލBr�����"���W��:XLHv�C`�?0CP`c���V��,+YdM�F�L�J���~<��)�T��I�K]�qm�����:�*�s~����FBc�Ï���7yaBOI�AA慺�W@�A��x!�*���F���	�"��h���B�0kee��x��w���P0Z������d�p���f�]ya�GE����Orq^M��ʐ88��.η,Z	�*ښ���ld�
�Gb�F_ƍ��Y_b����y9�"Ҽ310�/�Ҍ@%)�B���;�c&��FE��S�����)�q8�V�X��1��H'�Y@���	2�71ܬu��k�La>��s�՚��F	oN9_?&����1��,�R�y�SرY�~l�.��H����B��/y���3* {O�)l�qx�N�>M8��l��t�{{?��K?����5���{�	����������ǽ�9���M���h� ��n�&�Dף��)��z��'�]��2OA���䁨`2�&�|{K	�읖�]�dU�7-�<7�gS<Y�[�<��G�~��R���W��B3�]���3��I�H�-�S�V3�@
D$ˢ�^V���H��Wɪm���<������`5�u?y�D��C�
Wa��KP�,�A"+_�,����]��O؆���`r�y��_�vŝ9�cφ���N�w�+�|�u�qj��92���qz�nz�A��R�X�cU� ψwE[�b�� \z�A��<�
�޼�����p~��� VN
C��!�ٜφ���߂��$xs4#e��-�c��E0�Z^U�|��������ێk]��[ڿ1,x�S���g�Wŗ�9att�ҩT<�K��M!�����2��w��L��@��[�q�_/ �M	�nP<	���}zߠe���˥�;JE�2�6���,��LSA�J/Μ���ߎ���#�Ϯ~�ƭk_� *w箺���P@7n�عp�'�/��Yo�������MZ�h`Ȯ}?�%)7,wS���M�!{Xa]�_/X���n(-m*	��zwE�e����s�dUE�Zذ�Q1J�e%�<G����S¡���X`�ZZ<*��H�`�cϩ2!���ڳ�?M���$�!�B-�O�y*B��kk<�9�6��yf=T��P�c���/b�;E�	~��)���)a���B�-�B�<d�#�H�rR�/	9�
�Օ�O�՜��W&�Ϟuׯ�ܝ{�q���� �蹓���{/h��N�r<�z%P���:::p�ն7�� RK0��a�e?��*���3+ѭPj��Z�Ct2�Ɣ��Q���9Υ|8Պ ��7���B~OJ_�ע��ٹU/D�؂p<4O?ᘜ�֩s���o[o/֖����s��w�0!Z�#�=D���:�Ζȭ�ɠ�q���a}c5�jЁ ����ェؠ�0uׅR�zCk����~Gp�.�h��U8�VC�y���a)���/�II�c�����
T��Z��������=�����^PScT���ۼu��G_}�����Q��y�
��?���l�|�k����w{�X_�x��z+���;�xzE�Mg& ���*���x�5��������Q]���T'�H�:M)t���h¥#����F��NV-��?!d��
�ɱ�8`���O�Ů�桽�!�T��J{f�"4��K�Ҙ���5*����ǳP����0M��zkP���A�u�[��p_'\㳹�8�B���t�M��� ���!�8 �n�	{�03��z���3�k�C��.C.���W�z�A��|�X��M���>�{��F�q1��������bn���瘞���Y�wo�,�!��]ַO�5/`1�'�#����
�ɠ��s�p����`m��=�`���gK�hK
��v�4R�Hj��G����A�����p�c4>��,�7�W�qF{zE+&�y�K��ʐ�����eU����� Q�S��\w�mwB�Z`��Z5�(;�t���������
�v���}�:���~.P�Ƽ�?X��@�0GV��M�ԍ�Y,�Q�
4,��N��a)�tJ�~Qyc��q`��'֧	�6B�i��B���Z�����ؒ���I���:��K�z�@����1�'��%ЂX�;�Fn�ށ;{n�wD��^��[�[�]�t�����E��:I�O]u��������F���Ȗ�*;
4$�No�Yd�#�d���M��?����Yv�sx$7A��Q��u#^E��^T"e�Bi�0�T�s?����k=�>�=���y�z  �x�Ʊ�X!���A�W�bĬgX�\����fT�`-a3��Z'M�!��[�v_�d��TD�M�Q�h[**��G����!ϏV��$2���v&!��{�[�њR�*�YSώ�wwI���5B��>��me�̍''Dqap�(�,��!wL#b���R�� �Ki	&��1��\�2����Q���!��.�,S�%se���z,�C���4�0�B�!x#kÄ]�z:�-���TO��hD�c��!�^6�k`�)$N�"1h��rAW(L��$�E��6�~p��-�th���vt��5��MԀ[�X�ܕ�VK�̅r�4)l�:6�!�w��+a)�*���ު*����m��Q��	l�=ݸ���#+�b^���RV.by�*x���X�o��b�7+g��v�6/ܽ{������s���[w����*6�)���|,�v���Z9[_?�����d�q?�@���lq$�n^�X��,Q[��
E�u�@��*�\�!�y��5�=G*lÁ�AX����<JZ��ǖ����L@���fX�9[��=L�8�
�>�Z�1�O��Ÿ=�|c��9E�٢0V?�`�j��6O�k��@HX8��Z����1�E/��8@����[�h�NRP8�D<���(�&m[���H��+}H�0�`�	�,��#��c�n(!�x����[��o�n%#�|��G�Д6X�`���� �%�Kg�����`E�y��rR��ւ���'HB�i��߻g���(���)G�Rh���M�+[k���`���T1��2��8U6>�U�o�sN󖞅P��5�CH��R.��Kr�Vs>��GK.��-:�yk���m��h�-��F��J8<�փdZ�RY��,Zc�8�i���rh�p�&�s#���v퇮ߺ��;w~r��ُ����SU@~0z����3�m}~0X=urr, ��4:9��P�;-�ʙ�=���-)�<���������,��,AKeM(?	M)��:[�Y�y�s�x�h��0�%oBH#�ac�LSz��\L滤������/�XWP�k�ZR+���s��!�ХGXKE��8^�$kY�֘���6䢴����%�J(e�,��2��e�R����m^�~'!�d
B�&���.(���/�>_B&�D��!��1����w�&;�?��a��2��ח��8r/0���yD#�5���sD���N�<b|v��N��-�~������G��s%�3h�:$*�@�3�<�����\���l0�:�k�G�9�]D*���hC���K{D�B4ʫ2��:^+7&�=��`��E�E�o�U@Z2)���[�+��B��ot==_^�VVɘ��p}e$���K�y���n��+�X�������O0r�^]�۽���7o~�_����nݺx�ڕ+���U�Z����O�Vx�d1J��w�;����\��� ��u�-۠�f]%�{A8�	S~�1����,9[�M=d(�6QM� �0hh�6�� ��g�<�(�Ur��g�sb�8/�@�E�iJ�>��Ⱥ��W7ӷ�j���W4�N��߹s��b�.r0���ҟy��H�8��7
g�2`��k�ԶqѨ���(y}���ډ��$rcٻJ@��$y��]i�7R���QS\OI򭭍0��BƳ�5�q}�9@���<�ϒ|�ݯ���#o�p,�x0��Νc�9�HT�M֖k�pP f��r"��Qx�����YD�a �*�T &��SP�,�>�����rt|<�ڿ��5	t�q;�w�n��F�A�x̹�s�|���܃�����g��yҬ~��Qk�(,lK�bc��ʅ�_��� ?4�\����f��!�.l��<yaSt���/{�����!�f�p���.���JUm���i�O�hT��A~���-W�u�&�E9ll0Ih\x��IƋ��#7��a�Y����a�Yk7�#7G��Ͽ���'a�~J�OU����-/ >��)��x��޽玏F���f����
��=�/���^��Z��*�JnmZ�����q�[U�|)�E�ı�[�8�
BJ�,�y����T5�~5��a��r�A^����p��˫�gKĕd;p�5J@F�.g��͎Ff�'@���tDO�§L-�u-�)fyS�9�U,�wt�!'�/�����Q��֝�1�u����.��ss��~H� Ŕ`�AF}�5з����F읣�A@O�9vf�y}�ݶ�;�oH(��*h	�\h�л��(,���v�=3<��fR����x�oy�r2�h9��
l�hXV�q�]A��1�CyI���x<2�E�r�z��˗/{a<�s@Q�YX�hZ�s*/:�ei�hE���d��ŷ��n�¼\=��Eޛ�X�%�}���]b˭���fw�t�@�����D|�@|D�  (	b$#����ke�Y�gD�������c~��"eVIO"�.��Ŗ�>3;�$�oY�'XS���v�v��]���1���x����H&������o.ZsN��qI�{GD��e5��26�,�0X#1��2kQX���xk�Z��?��a{1}�'�}�w?����c��ߛ�裏���_��N&ҏ&��R�\y�˥ ��������$���}�d˳��.o"ӛ�A�v4�B�xc+ދ����򩤅�壍��\f��1�M�!돱�((\�(t��@� ��%�-Jۚ��m�ĀH$`J9-\1�\��h~�ۏӯ~����������ۚ"jK+o�$�-]�͌�u��o���{	a��I X y�]iC��/ϼ?�{�>�0e��ܚP򤻶�`�\hA�����lWb��`��$@.r�ն��xy�AK�j��#�����7ƛ�|�����'��ϱ7_;Z��AP��s��|�E.��h���Y=�d�?��o�C.B�4\�!�x��ӣWY�Mc�����<"�_�sG�_y�Ww�*�P۽���A�3֋f���o1���=xU����$b5.:#hH��{�������'.\�y�mzm���uCQ��g);��k�J3�;����$P��U�Zc-e�S�����sU���e��r�T�㐓O3Z9\�`|����:I����C)�!ϭӾe+�y���9	*B��$�1z��e�A�����/L,/]ה�G���f}����W�z� ������'�&��^߼��`��%��ŽG�7Ţ�s�����������ǨG�8]�E�4�ǠpJ�� �豎!=)�SAnՄ]Q8��M!@?�vY��K66�=5�C�"��F�v�i �x*D�]�a�*��ѽha
'�������_� �w/s�ۤ�鳮()2
t����Y܌��)T�| 1�����!ǘ�k制��\ �Z�z��a��^����l%N�C��r�ڡY�Ѕ!_��w�U�9���tȄ�	_]�*�����X����y<���_��������~�{G���u���g>�iN��.bu	b=�������)��A=�
�M.~�5����~?y��������7*xrE�0׬�-����=�y�`&�Ӱ8H�����C#d�xY-g<�����L)+��+�z�f�Z�����21\�4���}��SOe��>�1>�����Ȝ�>=v����(��5؞�*�0bl\Lc�G����������x�~��M=~������O&+�,<Y��6e�+����M��M�G֩4�c6M����a=+�*�V��Y�n���W<f�s�-����
^vk���VI��o���a�	b�����;|RKޠxj�K߄�T��1YsF��sk���7�IȜzR,�W�������$8z��0m9�W	�68O��7/�-�u�L�"!$�Jy�	]�O<c����"��S,ƒ�s}8���6�S+-�����iL	K�!������HL�	��.�0��۴�$P���k�J���C��\f��$̭�b-Co�U�n�v��i���M���tn�i�A�p���cuoj�#�|�u�a����:n:$��G���%���5/E�����k���\�1��FYKqk}H����7z���z���O�r�J���)m�*",�n[ͯ�P�F.�&����A��ͯ��W/Jk�Erc�U�S�͢��D��xQ�-7׷��5�k���������Z��
_s��..�8ÀuTi���~�φfc^���<�f��X�*=�t��_�}��q���{3ߟ)ͭ	�\E{����������
.�!��i��v{9���R5�Ϧ���_�>xߍ�������fsyy���?���������-����&�������ia��M#��#��zW��G�Sb	hA{�҃u�,71����;�z,ض{39��G�T�*2����5�=q�K��O�6
������q�}�u���$
m<r��ɣ�碪7e�j� S���wE�p{���N�sm�cN�#��_fJ3�Xjx����ҳ��O�V.FIbųC9IyX���˷�2@�/i,B�y���*���a��Y��i�1�,H�C�*�f���Ϸ(qJ5Q����|͹�0)���ύ�ujM<��;��������x�+G���%�
sP�^SsC��ŃVN�!�8K9WL���viBQc�؊q�>��I>�Ɓ����K�1"<5�Ӿ���aR*F��_��,�T���nvے���KHۓ�.r��<��>G��U.�Pc�@�SHD���j�E[��:�nf"QnO���ϻ��w���繜�39qK?��pgR���o���������(��O?����O��ɼy���
���K�٠/|24�P�ʅ h���M^�aQ�cLsj�?P�vv�RY��ӯI��c�7����Dg�ʵ)�	� OA֮�܇>D���:��3G���t7�]�����=Lg��Q;N���G�Y�R�_�%����0��ʇck�	���Mʹ�u�uE��Z*~*�f��AG.���LM<,D�	�*�t�6ڢ�^�Ķx7$�"�"��$\ͭ�l�#�z]iւ��*;yd��Q\5�v-)��}Y�2Z��R�mY��s�Z���9�dD31f��@>����р!���~I���uoA��ܯ_oM9����{�!#N��(�ݜsB��<R���-4�@�C����sJ4f)!��� �<���O��i�_���`�&l���������B\���Tz}cq���ғ��A�6CD��'[���*�Gٚˊ�4KyZ��o[geN����&�.e�=�4�((V�ch
�H���U��E�uv#P���R�6)#/n�1�R���©"hL^��_ܸ܀�"M��ow�ŸZX!�t5��O>�ˏ��Ǐ�z��sJ��E}��gnn���i����p��7�~m/�-�{|c�L���N����M1UrRPHX����TCVTiΦ�{����r��p��r.,t$0� 2���5���Y�%��C��܀�0���l�'[��⥄wR�Q
�;e:iÓn�o���y�� �_�g�Fk\�G�D*�I@����Ր��������?��"Eq�=�7�����F�!Lar�G�ْG���B؃�z.�����1���ʍN?�ӕ�Qr(���}��ݭ{xx��ڕ�*&�)��t�¬��X��ϊb���bo�P�����ŝD�l�W�t�k�b���u��j���׮+���:�;��E����ysLƑ���zR[	&�=�,�U�e��il��*U���dߋ@�`�/��0�6&ήݸrH�3gM�`{��ؤ`���󽕩r�� 	�3��\E7Z@ZrN�q��8cT����1՘�ӘA�TN���Z�m.=�VK�G|�����/�����~9A߹��/.���������4hZA�%o�͊��M��r5�����XZm��9�c�o]���7�}���&d֣$���2�~\�bW6�C�&r���L�^�l���~>��(�J�@� d4�Z��ux��fV��6T���r��Q�D���W�g���� ��,�?�}t�U�HQee�zpu[���h,č�6��c�|�ͱ#g�-so!���kԱD���sV���yŜ'���qp�<db^^�� �ΩP�Q�^I���6z߈� �1����8v�{�����ڼ� �w��?y��噍�8z�Wk؊��
�����*_e��k$�׻2���P�ā��zd��ֻ'yElyf��;w/-`�Ҿ��p����AV��:mVV�[绺sQ,sZ�s]����q}�5B�ֹ7�a����0yœ�*��bZ_�P��7��wVí$"ge�v+V�Q$uX�dgz�ː��ʽ�$�U�ƙpC�WH;\wۙǋ�,HY1F/�{��H���`�{N�=�cI�����[��CV��H���1Q��d��t@0*��k6fS?{]G4Du}F@J�jR����2�lQ��<8xۉ��l�{�����藿��{��>i�G�w���?����O���)�w���J���%q�-TbO���B����X&����EEK%��с�s
�ai�Fs�0Ϯ�a4��X9��<�n����<e������U����1�}�D6?��ˊ�6�6fia��v���GZIb)�A�dS
g���x��-~�ZϚۆ�D��5>�� A���ٹ�3l�I�S�������<��w��g�
��pdo��&,��/��q�����N�u�~k��~�o��^��=ː�9a��M��4TK7��jLT/���;1��,.q;{y���,�Z��onF��x�V���-)�P;�A���sRCϔՕ�*c�@�ti�y0|Sj/���E�z�ׯ�(�XE]�u�ބ�)C���Y�2Ҕ^�{�:t��'�C�"n����s|p}vQX�Z':��I��q����:��K�4��q���u��Q;oӶ<s��}�]l���s:0X�Wm؏9�c�)���cSzn�����3N�U�P��d.m6?x�������:}�-��s��_�⃛뛿1�]�D��\M�N�+��p��!�!�A�@>H^��
�<�VU7���b?����0Ò@���i�V���_/Ƃ��K�#��p���J�?[�Q�e�w��0�D�=�Z���W��XJWP�+X�eLjk�3&����V��%>����ϝ���H]VɍC�'h�Tg����,�y�cޜX�2��;��9�ړ�#A�9ì��!�֕�M��~/:��#��`B]�4�dK1���^�Uu�龇\W�s>������y�>Q����sՌl�7�b���saP0�xBxIZN����ݚEo%�Z��q�*Ϫ�l��ͨ��������NOl��My�JC]xy����r|N�,:�78<�R��ݖ{#��gx���\������5jP�hP،��BI�u���<bU�o�m�,��|���E{�8g�ѐ��a֥�+LYN������˴YU⋘h��v鵘������AjSҭS��G�82��%�7慌���Y�%䇏7{�F�S|oV��;�[3ZD��8/PugE���M��w��盞���gO�tR@�s��Y��ӻ������n��q3�߭��(���P�JhS 8ef�"��1Z]���cy�a�6�nU��W�����؃3Crй1���uᑌ��OBh��x�#ͼ��xr 9L��:�7	�1
P�\�)���6��Z����'��<���u���,�{չǣ,��s/ҙr���
I�Q���V�ni� `�Ѷ���QZ�cf%�>��,-{�|��\S	=l6�r��n�x>��J:��B\^���U8Ȱ�����f.��4��Kx��i��t��aR�ZgRޓ�+h-�Ma]9E�lR^k~(�E�%��Vñ/�
��İ�u�����`5����P��>�q�^�Rw*�M1r(��1��<���xgR����^���5�)��L��������g�v���O���O�g'*<��R
x�s*�}"BN����>t�~��q��L��؉���+bg�V5C��ue$��v�+޲���	U!b.�x�ۚ�����Cì�&�����VƯ')c��D�R��ȉ��|��d�ѽåǂ����n����K�R����b�?����	N�8}��w����/]M���c��7�Z�c��_�x��>a��L����d�M"X<V���*"訞�S*.k�bp!�X�{&�貆U7��d)�c�]�X3���&|Hp�3[F-qs ]y������h�X 6���'Ԍc��$d��C`�;�� �RtB�r�K�V�65&�Z�v���[e��|W��5�;O��Xo�)��f%�Mv�@ڌ-�@���C-����U]Q��b;
<+��R�[y>cS��$_�!�exW)���S���(voӆ�'�x?����[�ݫ{��e��+t�Mλ�	�Zv>�C���	�.�V�g+�ո�<'Yұ�[{�aSűƣg�[n����0���������f��%����rx܃M�ف�����*���ZF�w���簌W�5���[�VR���X��*{K�A0AIZ%�I�
�ա�Aҥ�-���^�Y����*���	ǳ�3S>�1�"u��RU&������n������/Ɲ�7��1�T`�8ݟ�Ї~���w��w�)ޏQ֯kb��]tӾ�s�^������"]$�"�i���~<XGԺ^��D�k�F���<Lky�
ڷ�g���^�� %�Zdj��M90�2G�y.�ULL���S������e~�t����S����/�5ڸ�W�y��������������9O�VT@���4�?|����~��G��O�ӗ�;:�S��ѯ�m��N��V��*ʊ�us�A?x0���{,8�.�����x�b-jRgpG�@�@�hx�t��])�*�A��-We{)/��Xl2$�{�x��o��k@��M�?�M�7�v�EbX�Xb1�D
¬�n�-���MVu\�� s�}t>$HWrE#e��A,K��UX��{E
�'2���@���3±�T`���jR�X(�<#p)���_�}��D�ASfX��ܧ�J�{���Y"�ژ9���6
bj^޽S�<��l�I��YZ�Ͻ�Y �,���)��=&�θ�d}G�Hr}v�Y�2�*˯���c��J�7��W/M�j�u�\7@�X�:���+�K�bJ�N����M����׏�}��z>U�Pw��j>+�EY��7k�`p��U�5��f��#�~^�xfcFI*���˻Q�����/mt��0&�ݹ;�'��XR�c��s5~U+ÿھJ�~ڣO5Ѻ`ol�p��,wh'������yv��I*UD���yo.��,RT&d9K���KK�P�D�����;�q�z��?�>��z����?����ߘ��&�x�e+ˋ�0X�oTyzQi���y<�O��UWn�Zm[k�}���a�p��x
�e��3��&Sq8��3��L�\d6��1+TY��M&����@��&�B�6Ҹ������!�mn���[��m)t P��!��})�ǃqjg�	�C%y16%�I�/�}���9�Q�~g�����(i*@Db��wa���+�5�~]2�3�x8�8����0z�$�T��g%7ޭ3��F���rZ�@��D����"�%P[� ���7d$L��#{'E���U�aEbA���x,��ys���3�ܫ�>�G���<�&ޓ'��5��^���dC�7+}��M�._c�C���?N�s-���X�#�$A�C97�ѽ+�AϢ
	�"P�C����=���*k]s�1
%�?OLo�v�(on�h5�ͭ�%�`���|�9	�;�Ylfe���S��VFh��V�y�k�X�������<���Y��������њ&z"uo4r�˖z��Ň��|r����;S@��ӫ���s�Z�s{{�"��Њn����O) �b6��G���mPV$w5W�)���Z\�2l�`k"�p��p�U�^W��
���H>tvҢl<�)� ��d�Y��Q��rnѩ�qE8�-s
��}�M�)�TW��3��'���
�x���]�a��P�l�����)�e���G�GT�釠���^� �v[a�<Fz�<}g�������g���~D�a;�%��Y���[�iKg�An���Af�Z1?���2��}]�Ӹ����������K^���w�}����|<WE�\FT���Y�C����q����_����/����9U�ȔL6�hx��C��#��Fg�X�rU��Q�V������P���4@����r�uϼ��m]�I�mk�(�D����c�<�N�ढ़|M���A�9�����h���ٷtf6�hN��d4���U�~���R�f�O�ZswUUFP��Յ�y�����,���}��'�g?��o��O���
��w�}~g�?�Ѵ�`�s���m��呟�8�)τ|Y�ڌR:�)�R���q�T�Y���x\����P���+���:���	g���QΞYA�n��d_��&V,9yh�#S�|�s��mN �Z?�l7����I�IVt����y
���Z�^��B?�}`�=Q��J�O֣%��2:���Ϧ0Ȧ�V`H�Ձ��Ƴ�У�-��Pb��[�7Q��\6(	�F�\Ȃ�0\�"X?���nd�	�eL�6Y[�)��O`�=��BT �[�$n[<�W�#!�vx(K���b�2�x��=�{��޸/���EZv�a �Ȓm;g����j���e������9"�轆�r-�<,�p��a��*=���)�9A���%�ݣ��ղ��T&L7G,^fh�$��+�U�^��j-�=g��p7�ϊ��N�Ǜ�%lZ�xR(��Sb��c����\ꏮiMY�≥���yC��t~6ɸkK`^�W�ڙ�%�%_!���l\�R��RBM�n��cX �P��(5�^</�[��������m:�J���+���w�����W��5}�I���D��G�������L�p��r/�����id�SI��h�
�g@U����Z�c�W4I1��m\�Z��%�¾
<[xC�F�,.;���G���\!ծ����f��嶴Z����������3�E�2��(��O�e��|3c�DƝ�.�
�+{x.%�m]!��!����>p�l���*��*8�����9U]CƋ�BVτ��c�����sS��
�3o��J�2����L�	�J�r���:p�{�eW��xe���� ��o��hz��e�U��^@Z�WlO���4L�]�{��^-���K �1.��v�V��:�m��!WD�{��ߔf�d�U��֔��-�8`�I0�3��y��2���j���|���̕�Y�:V��⽹�V;���1(�o[W��o$��&=�1��9�<��`�=�,�aR���Z�	Ap֝��w�>�J�u��~�G��(*�?
�O��_>���xx�PV��>/_��^"�����⵺qZ5릶K���*�,�.��������%ţ��(��,k�w�FQ�lJ�ƋO*�t�}3Z��S���ӼZ���6i_cMO�Ʀo/Y�!�� ��n�!��o�p_���e#p����C�Yघ�æ�\���T����<�����P���uD��"�Hk��ފ<�T箯��g1���Mm-+~(��sl��u����/.j#���xl��x�8Fg���n_�1V��4[�gS��}�n1�&�X����T��Z-�u�30��yQZ:�x���q+gqI���U�X�HJ�E�1�޼��3A��D��X���*@�s��a�9XǶ�[gG�k��
2���b��0���io�7Bm����
Zb� uI���1'�J��d�m���e�h@�O���U:��Ch-y�����V�ǮCw�����k�l�����R�}���ۭ�y...Ӌ��*�6�wV�y���6r���6��������>J���(��?��x}s�'辂�.Pv6x��J�_jVx­�ꭠ���S���RGoi[N��!��tļ%�h�(V?�	��g�:����O��$���#2�t�O=*���i��AQ^�L��ED ���;����`��g��ښ�#�K�q�+���k�=��E`��(MR��9�L��荠��[�g
�gq�׾(9,R�����q5(f�*��e�L$f���/�5�$Q̕~H�d�#�S��={3��vh�-�'��Tb<N�{��<}6��gDn�[����=_�s�bc����s{o��-����X�U��&��R������S@p��
��fl1��Y݊�{��ޗ�&/G�y'��t6K�F����s�u*�[�n]X�.��b0J��R=Z�'��q���T���}S�q\/�	�Eư�J��t��2M3�~��sj�m.�w�֨p����<M���Y��u��_���2����i>ܦ�||'
���/�ܼz���׫sc��&A���t$o'��lDmϔ����߷@!��c�/lo�� �����M����\�ci�y���Lppݶ�%��0ꋠ�3�痫���p�<b�=}�Ą�Ƅ�>����Y�l�:��٦���d�����7��E��Y[*���e�ϐ�{Q$�i�H�(��������嬘T*(H�X����B�����ʂ�Y��P�;1Q7%�!�|�t��Թի8'��])]�_��T���\Cۋ�/��i$B`��x��F�[������S(\Z
��QE�9/���w�K'=|��֚ -� ���<�_<-�{Z�<�k����v�X���<����e��������ܣ�䭴�vUNG�� E�QB�*��z����n���ׯ��x�d�W�0d��^\��q��`(1Ɛm����Ƴ�4��d�&����O������gk1?1Bŷ`Z^Q��q�G�yf`�B���-��rʑ�C,R�	����3/ŭ�����t��UZuM6�l/���G�>���/�lz��}����f���������`~�eW��܆ ���ذQ1`�� ��b�� �&*-�&X��Y�,huC�!.�GTkO!�ƊW�\S���5�,RHQ$,B�ű�J���E�ť�����s�Q)Gk�jQAF���})	mH�Ƹ3>q��d��
�%����1�=�H;戴u	�����߬)��,1�=��7Cl���|�SD�����wF�n�' ҃  ��IDAT��Ld�m����ě
�r�~�cz��E�G� p(��|Dq�8+�q�T �ef��9�ݶ������������� ,K���CQ��P�~�����ϼͤ�I������:5^��2m��%��g�d��/�]7�=9=Ͼ�[�v�3�1�����7�7��;�������������"�Bȓ��w��h�����$/4yA��;8޺Z���_?y��c��؏������v����ݭ�3ǖ%~����ií #@ܿԦ�d�����3�aq�鷵^o<�˅]o���"��N)���C�ݑ6���dӛ��-��\�@� ��^_�,�v���K�΂�#���h�l���,�U��ϱ�s-���@`�(`k�]*dbsAWm�����q�PQt��c���b�w�ɯ�3���벩x�no�XV�%�%ۭ�Yl%*I�P�0��NՁM�,�b,XEk��=�X�ꧢ��A�z'O+E-��ި_�z�8%I�%��=H<6�T	c�2�4@�V��eo}eq�Ƃ�c�Y�""@c�"isp��zP�����8k<R��ݮ�C>�< �k����rJA���7;,�R��p>X��^	��l&|p�i" ���N{MP����t����apCQ�<�hkR����(� ��y*�ol��&�WT�i�v޶¼R@�4l�6�f��_�~11��'��u�sJ^�V��_�XU��B�M6�hħ���ddg��Y�h?��/~����ߦ�|�u���닗/^��i�_���L[�}��%@H�7�Z&gN�8�3M���AoG����=�k�����9�����C��ՙi.�sR�,�6���-b�n}��P�~�ݬ�6V(��!ƛ��XE��,b@�{\Rj��DF>�05a�TE��+�XɏL�H{�zmm;�P
9Cď��<�<�h8 Px�f��ڪ���s���5=���~��l�p����Ͼ��]��H�/k|��ERYjc�V�ڴ��-�7� �F�G���|s]��ax7V�m�������v�+A��x�nl5��@u-1��!ݻw�� )o�״�#�{����4���J(C#E�~���<݀�����)���>���?�4s}�k��t�]{���r��]O��o�KG�ڼ����h��E[�kڪ���M��2L�d��X��2DRMֵx\�7�n'lV���~�ۏ��g�}�o����ߤ�x�u��W_޻y��m�\�'��%�d,���T�ͪ�*E���Ն�n�uEL���5���1�g���l��^Sk��sO�=	ϟ������Q��\��0��7���g�g q���sc�¸��������,4c
.Ί����h(!�&�?�ˉ^E��K�2g#��w�C���Q���}AJ T�"X=W�uB�')�ok�qy�u����g��X)�x^�&���TƟձ3I:Z~�΂dZ��!��͕�V�
�wR�1���uk�\�}��`�EH�r�֛�\�g��-���S�;�Z093�����>�{[�0Ţ����؛	(�uJ�M�a��fc�-��������)%D��q�7������O���o�h���Ky-MBt��d*���0�Y{��}�>0e���:]޹J��y`1F��0
-�U*�T#��13�����ZF�����B�R>�lH&��1"AN�����`M�*S�7�4�̎#F^֥+*(j����^m3#�'�t0���Ԯ֫�/>�䯩w��ҿ�
h|��������ogc�D��Ǫ�Mȴ��Qxpo�����z8*8�@�YC��Y���ܳ�K�����'�	+����1��)ni��y�$���:/
��0��ǣ�+��_��,�]�!��Y`�/pz`�X5K�m�1�f�
��3�l��gFu�W`5M�����X�/�����Όǘ{���t�]e'���Vo����(��jY�C�F��(���Q�״5ɺEq��y2o��'z����¾B� �F/>�q��|�oxgg�=���=��a�A�@A�Xx�C%b���ƽ	dmƲ?T[���s��GC�}|t�K��{o���<~��j�4mϱ�J"��sE�U��[�h�I�����c��5�<�+��b9�?�hJ��	��SK�%��W��m�����=4����>Z�Iq8?���e���Y�����/��[>ު���^>y��?].����+rBh�U083^�6,\�� �C�����'ߊ�v��i��3�2�Q�Mz�?w�u�� *�r?��P<#<:M,�b.RN�h��-�ꎣD���:�~:���6o�cް�1r�����Y�MS�+�EhXu��ҕEI��(`i�u�7��bA�iQ�:o״3�e���^<k�1)��;f�g��F'���׃�X���EIX伦�����j��}�}�H3��t���6��B����C�/k���u��&"G�8J�Ϲ�lgLEV�ڇs�������D�ԩ��V���M܇�&��N}��
�cQ�lD8k�64����h��/�������H
����3�vY��Q�7�t�U8]�S�Tb@� �k�}_y�m�Ϩ���yb���ݏ�`쩁����O1Tr�Gձ��bh���⾧��\�^Ϸ��V�^:��-�>�Wj�we�U��`F��{suu���G�ܞ�*���gϟ��v�8�
�J��߮�V���
��6������%6t�C8���0��d.0�rel&ϔ��R����G]`L���Ya4�R1Ј��+t��_��q����B�r\��M#*4V�6a��£AX`9�80��S ���r��x�R��bKxW������ɕ⴨X�h'��!&�Y���J3ZOKy�
�5�6�c��E[�n�e赺��m�u����n�rA&\�6��d��M��Y�(�+�ʕ��E*k�#T�����Te]�>�&�)��}�.L��ꂷ!8�թ�2Ul���RK������4H~��4����1�j���T�a݉aec?���,D�fMi=q�T(�qݧ*/����u�6�D+����8�'c��Ó�Y/�軺���d�$T�91��_	R*ܹ,(s�k�v��i,Q�7L�ߩY���5���Ƒ�cA P0���]���83�^h����7	T.�֦�E j�F3�H�����}﫯>�����g��۬�V��?>;��w���Z���(��y���=	�~�p�5y�>K��]���n:�sG��$���kA�1M�"�g���`u
������V�Ce��#�T�����2ݯ��6v�����+!���ʕ=��bu��DW<��;�gE�o�>��}���o�#����{�����s�1����zu�yKS��I����S��ɳ�,�!�z�(���]��Fbk^^���H�G6��\�*���	$&��x��GVnj����={.%Ǚ �ވ��m}��ej�w2*��$$$t.Μ!*a��ޚj/�(pDo=z�g�\�0��<�b�Ӑ�^;�-%���U���v+��R=/5�S��lM��L��/�E�g}u�eY�Z��f��6��.�$:��B�&R��gt�^�	#u�=wo[���<�i�o^�Z��'_��P�����+����D���16�}�o<1s����S<�ٓ�ID�*Y���Y?��q��ɛ���b�	�OXev�D�	�Ӟ?�Ɖ�%�
�*����M:����˅�������[5\���i�fj_���^tow�����k��:�Յ�w���:�,K�ݝr��&e��޴w7^�r�r~�z6��'m��sP���v�u娰�.ˌ��|�4�9\����}_�fu��2��>��FG��J������Й��j�Ǝ�Am;�v1����s�K~���0�����0�bn<Mo�xk
h�������0ߟܦ�[��E:��ɸo瘵�#c�eaP01~Q��p�8tV�݅���p�^b ��GO!�bc���,k���\z���M���95��-
E��-������cZb?��:�9��k@O:"��3�����_�rl BB�آgZ�� �qU��Β7�J3'߇<$�qČ�'cϕ�7uMm�a�� ���z�����lj�7��T����!�C�\N���ͺ���ZΕ-x��m|���y��j�Y��>�:U�Y;z�F�����{��s\^�ᱲj�.@��ɨ\��a�6{ό;����Ar'���)̳M�ӑ�WI�D�"�X�}Y�>��IT�m�%��FӴ^�;�RbC��+�T�g6(SH.7�F.�ax*|&�x*�Ħ	dW<sZ���J�5&C�ڕ6�4��f�yF'Q�P�s�����YZ�,�%�ζԘ�0�E�6֮&��2@�b�/���6D�We+A�f�w�HP�<�?��/W��������p��'���i�(�ֵ}�'(췱��7w�' \����n��@R ����8��\+Ϛ�{+��᧰�����z��J�K���Y��D�4��jDa��=dկ�P�r�
m&J� 3���D�?�zU�<��=�]��g8��%y9q�!����;��q�RLXӌ�����h^��B�*��
a��Lig6B+1���E�EB[F�=�����9�2e�w�챒b�!��ok_�֜�SȄ���a�DH�j�}�{�䩱%�ߡcg��U�`uk�/5�/ g3�^ã�=S�tJ��ogr63BF	�HBy/������֕d���~��L�|���n��5{2�#��k�:�7f�qy�(EK��� �#&�s��<�[pb��U�c7�/���,������V��k%�m�&<��¦�ڱ���uD�Q�_��=Y��&���r���Z�8W՟L���5~���O�jB�[S@�^}y���˟,�Ņ�!�j�ñ._ܝ	�6��-�N�h�9e�I����7��+k��d�~;��6%^B2n�oS�e��0q��B�a�K���^\��P̶!2�nE�V���q����i�/��Oumu��Y`�D�-�
͏bY���Qj�Vc�%�f<|�(`��1��(�&$�����4��s��X�܃	�ܸ����gda/�It�.3�(:Y��	�h�Ul>(�/�;aa}���e�Oи2��g1g:rp�h` x�9f@��ygz�6L3�(1��":�un����(�{@���~������\\��￲���%a�{D6���}���TMHv#�Q�_�����ؑ�
�!OK^�~���e,F���FÁg���0������j�2ʳ��k�o[�ʌ�SD��W�;x�Tա4��u�U���_må�
K���6�[�IUj�[fh����In?|��ك�����^�x�Y.��M�Ye'-��^�1{;����U#���c�\=�Ek�&����°O�s+�]d���ç@m^	�Brٍ�p��s(y�o�zo,&��6�<ZiN&�T�X�4��1Og��M�ܪ΋��?X�4Pûd|9'^J#B5O��M����(p��>���X��h"��y��9�RFX̧P�k�Y	�W���+�Z��Y�����C�<*3�>��/�1�$%LVM!p����Ĭl�+Q˽�q����!{J�$'H0�/ڜM��7�g�"�egyG�g��������J+)�����!T(��S���1d-[�����=����XŞRP��a�a�R{��y�~#�e�w!�==�b~K��ZL��p��p�!��]���Us�N�0�ъ�.K!T�e���\�ׅ�Aq����_X~����w�	k���N��7ӽ��y����r\�?y\��^�/�xo!9׳����8��7��3�ѡ�}Z��b�>e]6c�0��r+2}�==��<ߣk�e0
�f&W�l
�z����}����JH}k
��?��\/��b62�"��Z�:V�E����2sm@W8h�z�`�7�X-�S8��	����3B�Adb��bM�©�ò������I���`y��X،׏Vi�¸��{�'���É��A[-�)m-���@Ny���ֆ6���ԟ���+q��3�X(K轖���>��J8����ܐ8�X��T�ٗ2Q�[�}�L�`|��<У	�&t5�����>ͳ4�b,� X�-�qO���g�B�A^7�ƄR;f���1;�OI�:ί.��5�y��^����څ��qD�'k�J|�5��=:�Y�*�k��`�qb���qJ���7å[�y�\X,��A���g_���+mEh!��q~�I�hGD5L�wYY�v�v��?����(�\^b�aD{�ؼ[UT6�)��"�WR���ITl)0w_�;t�{���O'�������V�4�?�'�����ݻ�ݺ�ۨ��<eN�.�umk��<N��9��i��'�I>�7RsIv����6z��_Wfe�Y�E�g���ʋ�+��6�h�"��gC�������)�)���2��yN�(��cG���a�c�Zx;�(�|Ƙ� 8	<s]�}vq^�'�	|h���q�+ω�½� ��2+Y��P���~L��F;5�߱w�7��x�]�T{�ƅ��YU��UU�>��&W��W�����Vc�(��s���M;� ��BaL*�3�ws0$%2��^U�p�q
�+�X:[zO��mK�#����f��?tV_&Y�E 
���4Ʊ��?��W/\�h+��.ǰ�{��<?.dɳ>(�{�=��Z�����;I��x�(́ y~�/�'h�k�&�uc����>7�e���E���+��kdp2�E�Gg�"��n0�
=z%��)����䳉�������:��?%gu��|w���ӧOiA�Ə����A9�no~8m�;c���1')��xS�My
�`�<���</�9��7�}/�n��j��H�� q
�ٙ��F�ޕ�X�x(�o|�,X�4`Š�&� $�Q-�Z�'Zس�ɖre�u%S���g� ��|�t]�{�N@�q��Ү��b��ma�3�(�F�)��+��5�!�|ed{�k܇���#�*~+J���(�X^S;��y#]�[�WJgAߟ�TB�!z�>�sL�������Ѳu���l� ���J��¾���!F��g��B� �W�s�u:���g��\܅u��z4�����������-���%��4J�Ҽ?f㣮�MG��ʍ�>k�����#ڀ��BA%¼�`��P�82>R��w���[f��[���`�,lG|�i^��u�Ōbo�=g�	rc���މ�k�|0E\�Z5G������ۛ����?kH�[9�$(V}߼7��0z�[,�����}�d��Y|�-�C�}Q���$\�v��/*7�9ߥ�<��x/����L��ٹťtx[�M�s ��j�m��+s�H5����<�Y6:/&�fz.���z�JO��5ILe�1N�+6�xT��I�k�8)趩�a��%v
�zѿzeקZcB30��4�ߠz{>I*��S+#/HZ��hqUL��i.r{�d���#Hm��Ob���7��	 ��K����4˹!�@6�{=���̓�u�����Ef�1@>�dV�QԇC��<L�AZ���z;(�=��4�۽w��
��r���`Ijl��u�Y8�X�࠹"!��k�=	�ĄPQ!x\�>���]���<\��^�Ί�{�ܽ�N�^Z���c���*=��Y���Y�XJBF�a��}�Nz��+�����E^�t��_� mM�=G�LdK�O�_�!�O��A1ǅ=���[{�(�)l]O��������	�%4���Ҭ/}�p^h�¤��G��ɐ1ڹ-�ɝ��l=w��`NHU
���f�6������F�~+
h��崠~0	�͢��-�r��z[�!���Fv!>g��m3SB6�����ɧG�UЅm?�G>�+XV��_g1S��U��XK��_ara��&��j&c<
�&\/2Ģ���k,��4Ҝ㽔\�,؄R���.�>cN�?��\��LR�Y�xc�ߨ�pzMJ2>�~�hu�P��<�K=�@6��:�N��;�ǞF�;�,Kʕ�3)"y��Aez���[�?���p�1�Pb?�G������=���T��H��5	����Y�#��Wo�}�➔�+%�#W�5�8��6a��O*��ϰN�S*S�|(k����}yyU� h����-�����>���zNq?18�9,�!��,�ٺ5�cufr������h�28C�5���j����m�k��@򘏩7Cv��2�i𱳴��X�.�(-}��5,���cד�Z��x�ٳ��[:ފ��~��4��i��N�CP����)AJI}CS��~�-�(�"kΏ!,�>`6H�d��	%F�H�]�Ʉ�K�d���OƳ/�=V��%�S��ME���D����I5�(�Y�̍��A5��Z\@�X�</^�������)#:�F)�>����e��b�h�@�.n��TJn$D�U��1Gɾ�$#:P5������{wKf|! ��џs<�dU��\b)��!?Fy�P�M��63 ��$�������)x��"��ƥ���y�zLaޚ#ΉY�+�ZT����]t+gr�*W�θ;��G[��?�����w�( �SC�X�B��U�w�
ﳌQ;Z=�UZ��Y$o[0Z�;�z}4�A=o]zRm2oHl9���,7��7�񩲅n��䋐p܃�#{d������͆���7�ӜR���� �c�؁��g���>�)|3�c�:��ANcw4�)�O��̚���ڠ��d�t~Zt_.7�<�:~��t����ݟ��g��Q��(�/^]M��4+#	���iQ8�<�E��b)0\��~~��[�1>dd���u�@��.v�s�7v�鱚���2~�kS��Ʈ"���C�c��)4�K^W�U��q�tJd`������ <g<�8�V����_*Y��-�>������:��,�_�0u ��jk�W��1��=��Oy���f��ua��E�.o�;��Q�I��vMI���\�i�LJL���62��!���@77�%U�v�����u�Z*pJۖ�8�?�����¤���hF�;��w�����&��I.b��jb�>+�e^-��o��{�z��=��ރ��=2���~lס� ,�g�/��L��}=��-O�`=�Y�#�F \�ҁI�'z:���>N��z��&�^Ǳi+��L�&&ڷ�ֳ�ٺ�36�R�*f�)�F�9h�2(����e.���O�{5�T�gzm���gO�pKm���
H-��ſ����xozȮ��L0-�e����e��C�@�;�[N�0/�3���x-��"�������3��$�0FT�2\`�ҔE��cG��4��Rv�h��4�C��oBlj,ʢ삻�����M�g�qmL��z����F��c0}�%p�Q������AqQ2�r��t~�%�H��ŇnjlK3�cb� =���Ql����ri��e@7�m|���ed�0�fM�5�6����tD"��ޗ�:��S篩���k���������8:�˩@u9� /�Ii&�5V�9��Z`������x�(��v�!���X<f:tV(x���k6Ve��@e@�@��LalW�s�v�k�03x�q��������4�&�9=�*
X�e��|��!��\M�;$ۋ��]{�}ɇ�$Tw���,�O{Hތb:V��(��0P[2#0��-aܝ�����#e�g->�'c�5�������)|���77ۋ���>�:�.��\@7r%�c�-J��k�lnn�ߟ��[a½q4�����O^�b0Z�,	zX]���ٕoqZ��h����רV�Y���hD�ZͶ��{H�쳺E�%97���[�s����&��t�C.R��&����,��"Ѐ�B�����(}N��r6�����Xv�P����
��^I�����xP(>y.�k<��(��t}�"tO�n�H�5)�'!�@{w^6�b3f9�C��,�:mc�X�u�5��3s��־}/xoq-I���{���8D�-��ߋc�;{)�vJN��<ɋr�(8�WӘ��($��	��i�	/��7��=c>�v��f�)�zW� �٣3�z[�@�#����/���:tK�����P����#�b+��	�mVJ�F��BJi*���K$# ʓ�g#et�ɼ{���V���^�X�k�݄J��*���°R��^R�To^��g����`��_}��[A���I'�����`z������2��0j�4���Y�Y�Ε�7vx?P�Y���5�Y?w�ͼ\Jy9@p��L5 �&
�I�w(eQ�� M�����x�t��q;�bXpq��J2p���9��M!�XTQ\L&�B,^��� �Q@Z����Mn4��a֢[�C�3��OhZ�8�{㚌3�q��d	c�ZO�Y>��Ξe_��P{��i�k������m�Ӻ�!4��_�ź�6VE������\
&�LO-�n�*��!�q�����z^�<��{�dQ���5��UZ]5[o�����
z�Ӻ'b��4TD�����$[�p:�c��Oc=cgЛ6�ޕx]7�L��;Zܚ�N�_)P�/5�#&���6Q��eǮxx�z��O�#�e��ҭ5�0�\Ѧ��#h�y���׍߼/ښ`ʘEy��J�\v�w(�=4�3c|4�ǌ��!<G?��x���_N������&��o\Myu<�?�tc���&�GH_d����
�[`c�]Z�զƕ�J=N��G�W7��k�zt{������f����+���g1,�����`�xS��ʦyiI����u�
�0�J٩���`^{��&�΄w�p� J�F�@x^z]�Rˠ�0E�8\QcB���鷄����~��׶�ټPt�y�����A 4�Z���V�L!�I���5j�Q����%Pk^�Yz��Ȃ��m�,���F��57��
#��-s�4QSGo�-;뭂�,���(B�-�*P��BN�rB%gt��J��Z��E����~2Q�պ@�Ժ����ÙP�z�t��Kߏ"�`b1��#�D�H�'p��ymݽ/���I�/�#[��P�!�6Y�Y��ֶ;C%$�׹� �LOT�U����~f� Oz�� �4�5�Rňb�s4k� P]G��~�=Zjg��o�D�]���P���_/�o��D�q����\��bƘpOܩ¢)�W�]�I�_S��#��W���n��W�_=~+EI߸�n_�MV���v�^){~z�E.j�:��������v���-�ބ�z��"���}j���L����>iF�?�,n������_�؞&b��MH/���U]uk�)Y�MW��4'���Mi~��������!��-�����V�����,L	���x����l�N^�1w��%3�7 ׵.�+UTj	��1z9�L�i�5����X�
{>�]�$�f�
|���*��w,�`-D�,8�デ��`�1��n�3�T���cR����<_�0%��?�+({kf�f��X�����S���a�0�,�C��P�zxu��!U�PrU���c�)%!����cn-p��C�{����棭A��1�?�����y�$pK[9L�XI��)%=����v��7��:����\f��\QX�4�kt�JKd��G��-�ɠ������>PN3u�#gL9�kZ�굥`����i=ޙ��.��[5�i�m�W��A��޽�~���X��c�hl�ҸL��y� i�
NM8`u�e�I5�������x�;�B�;CT>Gs�>=J<-���KO�6u�r$@�����Ç���?�{�8�b��#��g��K���3�&��܍�h:����ɢ;9��=t��r�x���p�]X����?��
G�V�QU)�3�l[��"Z_���R=���4��:��]d��q�QJ<)�dzm\xux��ܧI�{����ٴ�vΰ��:^Wk+Djm���0}��������X/�U���ݙ�ͷB�~�
h��i`����\)t6��Xc[�~L�N���ڄ]�#�C���d��z16�u��%�ܢ ���s��>�V�5�Ę���pW>5N��җ�bq#�U߼��K<��6s�������ZZ좩U"�-B���ׁgA��`�q(�"b��r�ճ� cb�`Frs G`M�#���`�����Y�r����Q:a�,�?�J��}�j�E5�°�'�G�<6X�:��V�ρr�K����󲤌��DgPO��LJiS<;�����ꗽy��;���-y��L�>�u�f��HBa�PyF ���5q�fwJl=f�[/홏��/�/K�<�_h��ܳ>�������|�*�G�\�6����m9{�i�R�8.K<J�DkM����%�i��R�[�(Ց�'ed�/lL�%;����C :�tt��a��iFh��Y����ɑ�1���R�2J���$�T��W����s����8o�is	2/�3�u����X�k�/�󮲵�n��z��
5Vϋ�$bˠ�r��}��G�������7����n��?�Ǘ�C�O¸�v��Z��E�M;�E2@�S���kLA�P����,:9`��>�����Ea���g��6��v"��`�@�!��_���ׂ���-�s�մ���bL!�	L��+��c�-��s ��
�:b�
����$��0�����C��6c����i:AB��t@����:�M9����� ����t���6��jVQHH�눵f�����58c����+״�d���\�^�y�Bd`�4�P�2p6v)�։�������-N��C����J��9fP���S�Îy�I�:7ċyd*�A�.�hb.�U௸ƅ~�/_]�s�p㝆�2'�%Bo�0Ԫ ���	p�6�	������(74�qg?}*�]؛&���	o�����O�Z�QƸ�%�j&�! F�S�u2V��͉VM��z��7Ԁ�L������'ߟ��`��U@)��r������	�l���]nhr?a���gօ�|�p�[�(���zDq`9�`]D����j��� ��k�-k�5z�\�
��:�wk�q�l�#����(��(ۨ���ꅑ��ɄF:	
��c$A} :<��Lz]Gq6-J�\"�sXّA%%5��:�����N�}��9m5NN��a�M���2�&��c!_���L7��H
VC.����{��0�BT�o������.� 4�����r�:�t �G�{�pj<�\�r`-ǓCyxax�\�z}&����c^Y����\�١�� X�X��DE��ڄ(������4�\#�Wy<yzx�*Z�#���s��~)�`�,����Fߕ���?x��b�����앸��.��uߺ/Y����{Z��D%�Q�W�g0B�Y̷�*!)���3Q�;rC�v7vYC���r|}_��ï�<ި���w��nvw�}�����u�x&)�ET1���̮��(��cG�Y��2�Z������>���F�#'+҃��R#*z0n�Đ�0��f�62�>Fgi-�j��a�]�����Y�18���[e����t�*�9��x�"DQ1�P�Y��?1 �7)p&JƳ�%E�S�L/D�<|��`���x�Vl�..-��`.u�hH��6���pqŞ9?h�Aa�(�3=z�(�;��c|����ECqa�Kh�Vخ�����ȒW\IH�� X��0>�x��\]��o{�\�� �l�����4�c쳭GǶv��s )5�EhfO��|��~�{��6	�?&f��6���'tF�g�Yօ�������ܸ��5�"Ik����n�6�x\�쮼F��Ə��:�y�2����N�sZgSR��m�!"�ƕl�J*c&a��J޺����{��%e�(��k��r�k�:W�n@��;T�-�mWH�+U�{����*u�hΟ<y2�|}�U@���������A�L0����R|�+m��i�yN��ǃ��,�8u_P��J���l*$BBQ�E��{x\�`&^k����:��8(bMr����"i�x��)�x�����!�ӊ�V���B�ѓ��	���Ǧ��b���{�zNJ�`>6��2֑ͥ(��߻����z5�9(�D�)Z�q�u���;��Q���k�K�	���F� ������'�dKK�u��T��s;��i��Wu�X�9G�~#Vo�*��{6(j�I��ʸ�l-�bW���(�؄�4^K�D:3��!�~�{O��^#�х�z��Ӳ���Ҷ�O/���J�׋u��{I?��(���*����ǻ�1Ͱ��M����H��6(�`{.rU�d%��,KՇe�|�ӊ��H-��k��j�"=�/Q�PЛ+'�lw�'O{�^�=}�����n��������AV]dv�at�ƒD�ˈuk���.Ag�ʸA��$�x�){?sE��}�`ąYi���1 ��:�"1a��
��Q��5�6wR�x�'n
�ɂÊ�7�~��A_�����y���n��V\,f� o�d�g<<&��wA]�R�eǼ �1�@hK�M��8ཛྷ�~a��j}�V%WYXk�s�q$c�m|�d]+ -a�1��m7͊F��mE�ZB���h�3��'�� ��0{s�~ύg��1h}�q,g�V�F�,�7d���z�l����}2_e�T �-�n#�kU���wJ����F(�^2�V��b6禧J��bW���{F���am��-A��>�{�&Z�cf��s�ODEx�G�D�x�:�������܉G4耵�6���L.���	���>�φ��QƱ�>&�p-(k����ɼ����x�q_�-�EQgM�$�.�|����Q4Y���;=��9��䘃�:�0��,��F\�>.1��a�9�Z��?''ֶ�b�uY��3�9F�V��'n�ƀ >���j�l#��8q��P��AQ�أ5��ej��iâ���DA!ύj�()�0�p�0���̕C�5N�
�
0(��=ڸϽ�nQ+����g^��q�ubk�WLG�K���Og�M����}�u1��"���k�'8�6�c%��ƈ=� i������m���t��&^R��[,�C��֨~�눋鈕�Y�*���8�\8�j�(C����Ũ�~/7��?��p�� ����;����vu}y0�ه>b��4�2c���IA���@Hn��g�Ϗ���o��1\ަ&��ݙ\:1����ݭ��A��yϥ����̤t�h��9e�/I�Zl�n���oTM��;��W���I�V�e-�������[�ÍB8�1�a�6A�,$��\�\�ӏ�g���zf�h��H�D�� �^G����;Ц����kV}���.�`ᮗM�����a�b��{P�Yd��9�(��c�E�8�u�T�`��xM�w3# �������+QI��9�J,�zX�Pݧ[�i&Xm�]�@�_M��tϫ幽���������o	����C��a�R��!����Y�ӏ��rA@?�яl?~<yI/gީ�C^�Ww�e�gc�C�ޅ��]gϱn�\8r�����(zg��3�A
��p�6���3�|q-Ǡ411�ݡ@V(�/�iJW�y]跞���,w��qTS@H3O��7�E�A@��k����偲Ɨ��R\T��k��'���D�g�PYC*���"�ݍ)�ݮO%q3��|L���}��!#�L��'f�a�ϼ�a��������D����>d/F/^�� �[YѪ&+��2�<�oٚok�39�D)&�Cm�̪��3u�az1=�g�^��d�7����o&�_.&?wu�i}�C����Z�,R7M�d��N퓮#Z&��ܺ��`�i܄Ϝ�>���KZ�ZlcQh:̢�傗�{C����g�k|~<��\���6&�
�9�V8O#6@�H����L�>51�0�bѥG�q�$%b��D[�����u-Տs/�r���A��,�`���1X�X��s(q	 �3� t�������'���|z������ZP)	�?�0�#�Y��ν�e̱�5k6�e���g��ҦZ�����3]��XR1�x>�f����b�Po���/z�Q�G���K"! Q��W�z�۠`#|������M���(>�����C���G��@�@��(F��w�\�\�<k[�� ሐ��{����Dm5i�8�p!��g!��7$��NC��Q��yk�7�w�����2����*���b������ȶߥC��S��H��D��R�|NoqYM�[js�3�ma �/�_,�v��|�l��`���R��W�.��8/�B�x��Ʃ���Xdp�-��f>6l�b�o����0��P���ݬ�[S+q�|g��}�xn ʺY����᱆]��2�}-�S�"@os���SbZY@�}�׉��zf�O�������w��]���O�o~�[SF��Vˍy @�M�鋸�h����g_Lh�������-++���u��頇���ke��h-¸9TW=[�W#p�h0��Ϙ���y����bQ��h(�z=��'�7��)�\$�B:����,sDU�
{�����*���C�
f��S3x&����Ez}��^{�:W̠ qb���[g|5��X{�{��8EcT�@"���!7~k�'����L�Ϙ!1���C��R.U�	5Iەة!=ņ|e,mO����Ȃ�$�&@�A���t�n���ş���/��O������*���8���)���AՕϲk�m�އbt]i�������t !�XfM}��B�����E1�Dl��@m5�3���V�-��P�@1��<g�u8T�NYpcmo�}�U�[��
���J����)���Ygx8�!Xb.��<���Z�F�:��7�P�_G�Zti)*���Y��F@K� �$9P��Ycn�����˟��_���/�H�w�� :���;��穙'�EKjo$��N^S�e�>��SD���,��^�n0�Z΍�֕`J&�����Gx��D�B��b<���O4Ƹ����J��v��c>ʓ�I���O�`��=x
A?��{íL��L`b��ò0UQ��X�|�Z�y֘���)P�9��g��-��h�-�̟�)߉|�o�x$�b��57��s�4�s<�e��0�q���(c"BTPcM�����Y,V����i4�5�\��Dui�a�B@��̃X��y��̖!1�8����EW!�+^�&\5��K�g�;=��ѝ�S��Ԇ䱶��������b-#�y�}A���-6��W�=�~P^�c�*"W�e7'y��:���>��s�Sh#zC:H�D���%yz�NV:�1�G����@��v02f���S���/�GXOkIJ��?�y�ꫯ쳂d����q�����V�΄�j����B��'�|6yCL���Z%���J��T�&���ӎ m
�3��M'����v�]4�z��^�{(W^dh,�ܱ֣����p����W��T���U�x�+�̹�A�*
@(d <ּ����ܮʠ�c(?��B��b4� ��_5ě�g�_�)�����r��Va�1Y{k�a�p����L0��l�|�G�?�
���3�Q�f��X/x�s;��D@�b\q����~����x�Y���Ja��Fc.�S&5��6�úI-LkL3�UHF8�4>��Ν�֏�c�pbQ�-���D�a�	d3b���m��ɞ�n`EE�h�]X��� ���V�w��-�����b��9>��8Gd'EjkT�ܣ�"�5Ǡ�U?f\�u6�X�h��7��%"��1+qB��5��H� Da�	����/~���o�`��~��y��=��p�^^��F��������1����o�
�߻����$e8}5\*������<%�YL�G�ϓ�g) �����ߧs&�3q;}��抠N}�`��@��f��xO�@��'�o	����B8�b�^y���AwT�-����0<uD|n�imVC&4f�y�*yo(���VÙq;EWN�@ivO�����2)��d���<�LU����lm�~��=�V;w'O���v�r��E;i*)��X,��EK����֢��n��F��bHc���@+B�t�c�..�x�>ll�T��+U�C�q�²�~618��f��馈����J�DEj���9��m羟Ǡ6뚫��G��-�| ��.؅���D�A�G��`A�������Ra�nf����X �8�>�� X`�)��XM9h9��]XY�?������υ�zU*:0>x���{n1��;��1;^�>+���L�����_��w��0v��2�Wg&p��Bٚ��˽�x^��3��w������p-���k��pp
w:���h��Y�g��T������� +0�:H!���ȱn�P @4l�'��O~��#��������K�����a��PI"�XB�4xb���v��:�Rbo=9���f#��,�9ȗ�b����/���s^2+ʭ1���^SJ��XP<G<���C�E�wl{�E�����u���y+�)pQ-�!����A��:�~�(�� ��䐙Q��J���ڈ�K��b��y����Y�iz�{;�;{^�hb
����u��A�@��{Q|}�2`Ú���w�Y{������s��c����Q���4m�����Y`�(�^��",��cI�����֮}Q���@�1}a���X/ưN�1,b) }Fυ�$!wu��>w��+�f��C�{�w֗I���3kS��o���{�_]���+"��Lwr��5��RYB� ��?���HFB� ��b�A�;#[�UE�\���ͼ�y�Ngz�� ���o�q�	�[�bg�s�!b��k��Y���,�ϞW�|����s�ѓZy\�7���LcX>�{Q�A`sI�}��5cE�H���Vq��5=����ZX�Ӽ �Ț��_dz���j��XKB�DWB�3C�{ģ�C?+	�H�$��kU�������}�v��.�D��cJU���z��W�n����u�f~�0��X��`�ʒs��JM��0ǜb1_�����#��u�)�Qx��&��)ȗkw��^�����'�W�}>���|-�Ew{��Q8mk���$lR])1�A�ܵ���yx����J�����*�ۡ�ڂ؀����	<��v�������WX���3vޒ����>p�J�,�+�5�5[ӆ�k���|��V�c�36х��@TUc4����X#�^bW��_�!TyU���ZK`=�q��ҹ,F5L�����]�/��P�j�5����՜����>���� Fs��%���ə�;ν�����Y-�0�ң �j}Y������E?��RЀ�	jR2�ؘ,BD7l�����5TA>Z�'O���N�ӝ[7�e
8�L{{�#�e�F_|�� �N&y���h��zsC��9[̳!-[�ʙ_c�U���
���{o��q�h�_�H6[�])d	�-M`��"g(���ԚQXV�IC�й����Ws����NNc�����T�a~�oޱ\��CO.�H���Q����á���͛A�o���s`�P�"+�ܲ8؛f��td&�!��e�,�}�g}�r�{��
.-�D�S���I�M��zֶs�v����j�\���G?�ޝT����©��)����(h��-뙔���PY�������֓t9�E`��Ŗ�oР�_����3���+@Mש������n��m���wte3�1�td��8r��6`z����5�S7�F.pX��&jԲx=���Ū(�
ܦ�H(n's��#�o����հch�i��qP��OЕ�S��x�n��5��Ճ��;�NטK,Ah+V�|�7���{!G`��D��ͽ�N�뾣aV�v7
z@sE���������!�^�j�l*+GZ4��~Ęod�|X/}n`�7�������['��[����:O�p7��֢�Ÿ�J1�͞a_ZSDH8_D^��){�����>]��E�ډHb�5u ��ɽ�O����L��RE�Y~��uS]�ۻ/S��&�{�P��=��\�����<s���������m+~aA�^ry�>Ծֵ��g�`����� K��U2���Ӹ>��3��g���r�,׳�����>=���p������
���Z m/^��9�#3/&0�P�����b�B�ޯhQ즳��k�CI�������7U�n��|l�jp���hĤ�������
��
?�c�i!3�i��:����F��Na�s7�i~�L{�����@&,�BЃ����9
.*/f��bN�,� �&���8ͱ�� D8�gF{2��kh���� �ҭ?�V������g?��%W
ZRġ Z#
�ͧ.���]CG��~������ѽ�#w�����C5���dzn|M��@�k�{F�5��"|� �.�:��A"$dȳѠR4MB� �@Q�p�e�OP���p��|=�����~IY�*���Ñu�"s��h|��(ԕ/�'y�5��<t��ƛ}���|�o��z��)�+�����$(�ж�~�P�p�:v�� ׅ����D���~&W�pv��\�o3�0#_��T�(����P�GLV��q�u�,�&�g�^3M�錯T�}/1Ř(���9��L�����Ȱ�|�F����LI������e������٢�����X)A��:h�0�>G'�x��0�i3:��:��=Bw<[R�� L����U.���y�G�;	hQBH�o]-�Ȯh��@X�@O�`��JD�\��%a�ĵ�k�z֦��
]E"<3���F�KSN���}XE�����3�yQ�E�g ��E��l��� �U��g�[)
"�ߊ�#wg�)|ȅ�̠-��+(���(,�����cV
��́8U
�JUtw�]�;�瀵�JE�OM�i'�u%��"����g-����c���������z[�����0��O�䏏R����&8����;A>)���:E^�E�`9^<X	��7I�\�[ZՑ��M�ʻ�΄�+8<s|8�K"j�0���Kc�ˉZ�1��^�3,�ޓ�׽���z?�Nf%�n3h��8\�LC��(�v��xx`Z$���H���`�X��wt�u�I��Ɖ����ZT �̈u��X�H��XufE=<�B�����$�M���7��>}b��,���w;�2&sݝ�h����ۭk������g�fˎ/?���G7,s?Bo�'BN��Ys�}�b(�l^Z�����uZW�|Q�Zh�;�����-U`������K`�}�
�A�(�k���! X�q�՝;'�5w=��[ �q^�H]%�{�|����ڎk�´�����X�*�b�}��Y�=*^���X�-<$)'=�O|.Α����o����D�Tqo���\g��)���v I�d���T)A)�>;+���,r$�N��U��a,v$�B�י����|��ad�>0M|,�\<3iW0W,��B¹.V �P��GfՕ�D?2k���F�i�����hʣy�4��*L*V���EH��x&s���ʺF\���\�%xZa}hD`Q�?&@J)I4*	���8_~�i���*Wk'��5��yS��T,�-�1���t�\�"�״rE֟ϔ��q����~Ĩ�2�{�?�������
%�5���� �yh�5e�f%�(
�KJ���:�$Qy�H��J�8��:�g�Ӿ+�5�|��[��ٜSk���G�w�2��<;
�2�QٍJv��T^Us�t]�-#�<���\�uU��%���y�]|kP�����Q�6U����q�m�LU�����p�6���J{���js���seog����s
�Leh�McD�f�\�6g�mn;�u�sݝȅ��o�ss�{�"�a³��U�K�/4��*�bF;9z��=�T0F�3`2���YO�0�����ef����V�^�T�Q�8����L�/�ĺ�9��ơ�=��\�G��X���3bT��������G�����?12u�`�ym6{�����ktϥ��O�U����X���|��;�����;j©RH��*1�����V �q���́ @I�u�p�C���|�����k�)���M��`��U�5�Ѿ�d�v���QQb��7
?�������lάE�w��r�3<�kQᛉB9""Xx��[�b�F��?q��>އ�����J�o��`q�<fη��b3�h%0�,%$4�;(Ex����Ua�����,'�� ��P���wg��n�������Q����-�0&T�o7����|z9#3��_P�&�5��e�"C��M��iD�@�Q�F�8d���>-����o��G yXm��F�g<v���u��#6Ï���uJ��6��h�vttkn�K���?tG	�(<J��q�a�OܧUF+�5A��}� �ϊU��d�/�+t &	Y@���*D�͓'٪��u����G�<
�8w��R+M�����#A�n�B��Fx� ��n��-F�A��ϱRM�V�����Js>��$�Y�a��ڧ�wԦ��-_�+�<�B��J�ʩR�w|LX���m�g�5��"�ٯK����%8����B)t��<+@q�����}�mC���n\���L�_~���1���Cy����8�a���o� ��W���yEX)>\$��лwn�v�X9�ɖ���=L,,z2��B��:����mէT�T	XK��$�F�ݡ3"�#�Gc�_^+�)9�DР�z��M��",Ǐ^���ԷH���@��D��a�0R4I�3���d�#�`lDY�a6! �r8�<���TW+4���@Z�+}�i�y���g�u[J��0q@sMJ��O��`X��կ�Q)�ޛ�{���v�=�\4(5������{�U���}�H��dPJ����a-�V�Q��t�܈.dX]���U�������M3�fo�TU������X�����O��)*Q0BYi�E��뚣|�\�B���	�u��9z.o�����nګ�$�r�L�ϛ���2U6b���rm>g{rrd�AE���`�y���(dQ��p�'�p�ZV�Z/E�g��D* �����[�I��)�#�z;Z�}*����?�����k)�g�k߳H�E�x��
�����!�֜4����M6��v����4٩6�^�y���5B,����S� ���0�@����h�FfN�1���-�%	�P�������?���c�B�����!$�iD&-�hmF��m�t3�Q��c�q?�)�F�,�`���
���~��G�U�@����yf�(q������.UbX�����w	r�*���e_�&��(��g&���h}���Qj� e��,�*ЙAiM�i����!ٸ�й��%��Az��¢1����,��OE������w��F��Ê�o����Y��� ��g�0'���`XQ�%�p_�MB��Ju��
�uV׋֛%���Y)�F?m������uQ�<8S���|��;r�Z�7�q�R+��y�L�֒�hb�2b�N�h�(�C�'-���̳Es�&7oS�b��Rg��u0U(d���� �ن)sz�b�H�6�z�[���FS|���4=�]E�7��D m�R���3�U>��#�|��`w*>�,�eXJ����i�$P�N��	���H�(�8�>���%2��f7�E�N�0�"1�E1�>/�~"�C��QՐ����ީ~��ߘ���t��-Né+j�t,Ԇw�]��;o�:����6�o�4M��`9�ϋn*�A�H�x��"�.�N�Y������$K|�P�����`5f&Q�a����0���T�N4jJ��E�)�qo~�rlU܏:8 ΢~_lD(��:�[ڽ���
Pa��[�q�
�B��oU�s]�l�Ŋ�x||îʡ��xf�Yx�^��3ګԣ�\��j5�X4V�E�M�΅Iݧ,�pI�pe�SW�[�J#������.����x��BO�E�"���a�B�]��*#B�X�;��\�V0�qT�tᦿ�U�%A�B��!8�'�9� YT���OaдThBE�֊͵�ϡ0V��դ�@�#� �J�6[��h=��5����b9s�X�������	>"�H#hF�����*m&|����ZY��Bi��Z-׊V k���� �����eOs6�f����7m�S+Y�'s���1��D���?���E�����9��j���ƈ��:%S_����7�%�?�]�lՔ8hkk
�^�����G���r���6,�t1�DofK$��uA*tnH�ՙ��L�8?1{B��g�	��y�`=|o1`��{rr�9D�˘��yĩ���}�u����$�˲O|�Ogs��EQL�{���.%�W W#R��5^�xehx������r�\Y�(A=�k\��pu`�x�ߙu@�͢�{��)Ծ��Wy�_���>�ݥ�I`�3�>/-��ۿ���yK;����@�-0�W���A�Id����!ڥ�ш "�͆s�\���u�)��N���<]�+�~8��0&�:F� �!��Gs�5��c�3���iD�&j�S���na��m��O^SkI��y�yʲ&�F�!~	��<�k��7߲�,!u�y�I&�8�f4��ݧ�V	z������Қ���_���oL���$A���[��w�}�J�D�
k6���DNh +$Ht���0����CD���U�����@q�lD:�.2�(�i�(P#���;�j�͊����u�J�P����_	���Z�K���{�����a�ג�!g��so�w~~�?=A�3Y8u���zd��V���:�g���m.Y�Q�~�6���M�2e=M*D!;�Q�����-�o�$�����Hi�w�p&ҹ0���AIv[,NF�h6[^��Je��U;����m�ml��)�����!�Y	��/Zy3I�͇�Gy]�5L��:8L6u��/m}T�22���C����X0,��VP��)�P��P�����s��S$�.����B�F�rd���D��3ɧt�e>9����3X#�v��̶�ͭ��i������>,-h��?4�G�����=����U�:�`݀�hw XZF�bmr�������yi��Q�c� Z�Ѻ�ZUQ�`?��Y�X�#**ъ�bu�*�#�9Ѫm��<<W(!|^�iL~��
~�[\ ���A �%��s��"��ɟ!v6�i��H��/��[��'��,�^�+}�y��
���a��\�3�sh������7����7�����5B�%,wi}ߛT��r]].�t��chkʈY�*j�铴χAO�K�W����*�W����lx�'m�u K��$�fl��&,����A�bӌ��,�X�	�0�eH��p�r�X`J���*E�.�I�)�y��(�6<������{Ƶ��A��1'ָ@��zx0,��ъ��)s����e%:P������ꍇo4����M�ĩ�Z�J*����ѳ͓Eq���,�7L�h=$|����zl�ѝ����S�L�Yh�L����zhF3��(I��_��R�'�@8���.��'Bd0m�6ZD3BŢڍ��V�3{ՉnT�V���uT:��r[f+�(,����3��>�VU�OP�Ia��Ǩ]�S�˰v�X�ϵ�����ލ	&�.�w܃�[����$r'��n�ł�Ո�Y��Q�1��<�ko�<�+�T IiV
Z�vt6���H?,�w�ܼ��j��l��\n7�AK��b�l>�5I[�qT�/ &�_�^��W�RI(pA�}N?`n2;ߧ�%:+7�Z�<���g��/!g#Z��h���"<�}wߍ�V�|4�'�&�Y	���0n^G�E1��\�>�0�>1X ~'Bh���b��d��S��s!�g>0�B����ɡ�/�H���E�٣O�?Y����<��`���1��/b��d	zY9��������ۮ#U���XC1W��J� <�j�"�r�υ5t_Q4���)ZA�dȫ�t�SK��`1�U߃�F���B��d����Ĉ�Ș�޻����2��C<'�Őq�f�=X��r_��귭Y���a�/=�0`�|r��&�ϳ�'�t�Sb��3G/0H>?��pk�1_*J�}��fu�x)��Y!�k�-��J� bKKx�.�W;s)�"&u-X�oS��y7i� l����ft||k�h�m������<�~HZ� İgr�V�{e�_W~�;�>z�:�q��s�~����z��IP����m��k�a�7j���&aB��]���т7��n�һ��-�@�eUQFH���6AC�%�����z��?Y���3KƠ���/�7��1�o���Yӭ�T���[#^�[��{��!*��ȇ<�V��B���{���Yr Rr�t�t,0�J��FH!�6B�jG��́(0��c���RJ���].��,����tt슃E0)TzVUT�X�/M�Y)������Ϫ'O��dh�n>�o{�d�I���z�=�xD֝�o��<���H�U�ۯ�+K@�Gݹ����m=zd׻y��b�k��mD�ηnmz?�y�#�\����]��k��\�-\W�r������>��6[��V�Y�O+e����	�G�#=e�b�Z����3�}V�PR\�s���<J��5��J��݋�0�SRY�WYay���pd�����j2J�%���;��rf�j��;����u+�D����� p��"��^��pe�|�d�X��!�(�3kPg�Y'k&����XΗ�FV�����'������ ��\�QT�]�"��ݾ�1�
�+@�y��>,D�ϚNg^,�z�h�D�F]}��KkU|��m�tE��$�eܬ��q�������v#���G��NJ���A�5+sb��/�h*���~e�ay�T�qN�Ne��4/z�S�ƾ�#,�@An�{+k1Z*����A�i�'����G�$Tv�+k�=���n��)݁Y2����4}2X?-�w�R54�آ���g���,s3�zy�����ze�eZܥ�j*�"-��/��H8џ4k%��[O־��7t1��7k��$x���\�5�Mls��8�+�:A��J��8�}LԂ㹠{)v��z[c���k轓���'J�'��$�Ͼ*���~��9�J�+s����)�LF���8�Zյ��~�X�@\�ޠ'&�k	�O��,�}��O�|>C��<,U��by��5���Ui#n�?#�wa�RӤ��È^}���ZE�֡/�?��<o��W��ʔ����|�־�"i�ߵ�<a�p�6+��[u�z6�@�o�T��]/PW˗�.����<6��	��Lt7��c>����Y�w-2uܹ�kmM�W�g��p����Zz[է��QO<=A��|v��r/�{��|��n[��x��ۀg�(�5�Yn2��@�IL���TՁD���*�):��ר�@�h��StJG�A�ʣ��:�Z��eX
��9���Ai�S��.�$�u��M�x������m������g���z����/�xd�KU#�7�3�F�p�@������⑰������6�>g�k�%��+�����>`�%2����#g�fFП�I��D�F,ʚ��B�^yZ!���Qu~y��� 0&F�q�� T{�v"]@+���w�e�L���3�Ї9?r�1�~G�Eq:��m�E`��f��.rB<kl��k/a$�hL�㹈V��_W��`���B����5_����c@1�*l����b����I�{6�uM=��$O��W*����M�lZ��4R_�@�m�5qd�J��7� L��uH�Ƅۡ�����w�jt�F���ǡp����κ��B��q��z��(��p�׮+a����~-�[X��2[)h�\O#�t?1&J�Xp���D����X��&$�1?%2�-�3���Ou >3U"Њ��:FM�h.�Q9�[S^�D]��H4_���׹�s8(
O�{���bN؍��cc��QU�����.?��OL $a2���Y����g/���m�N����v��B����HX#_�e9#��s�E�d��#�1Q���0�󋍵��Ei�k��4�p�͸�:
� Ti���,��Dk7C���	��1��*���=M}��5{��3�}�KC�¹1Ā����WзY�ɷ��Ӫc�K��A�__;��|R�i������Ol�(s����5�xo�}��K$�_�D�:T��u3۴�o��X����t����ٹ�H���7�x��{�V>t0,��U��-j��&�4.A_[9L~X�w9��%2�����v³g��m�_�v���pz[F�U�ޏ��0T�΀2��]��͓d98��lJaM0o4L��rxTM1�֊��6��Ē�	ߏ�ebP�7V�J���Axa�p��5ڔ�9�?�5�O���X3tXI�seo����	���֓�oV��/�Eu{(�gf>��7���4ՙ�Yɸ�~W����V�E�-p �6Z#��Ȃ�\z=:	 =?ES���~<��?�g"��%P�A@
�Yk�*A���b%�Q&Arq���N�3�e��B	!�N��R*��#l5e��)�!�����D���A |�{��}#M!2映�yk�m�M֌���ʯ+(�0�\����:)��ܞ}�$�#����Z����+�ۙܕ��:���<�7�F4����YJ��)	M*�d�gX3�=����Pě���j\���SZ1�z��������SfU�
c��ɱ���F���8�#�7�D9��v.LJ��)�ଃ�g.���>Ga�N`�aL;��[r��YH0v݃R9�,m��P�`1"��<c A����>Qp�9�>�hS����;�`��nL���o���?������f\5����0�_�'o _,� T��b(�}��z �`��Eu$�`�a-~���6Iÿy�V^���{Ͼ/a�{��g���d�M^��uWq]�4X?�h5�^S%�g�3�A�9�kr�Abٰ���Dy!�MA܃(@�@X}�7tnBv[z^���c`��������Y/�.s�gb{l���O�5M����sp(_%���(��$\S��:��}	���:)k�k���j,�x��x_jj�T��³��)��u횉����>��H��U��6�6�nLHy�x�n8S�^�V��������,b{��H��:9a�Jf8���N�qy�|/=��ػޜ��sҡ�ӛ��M��"]�b��y��<�h-=�	_�愔�%5Kɫ8�7��i��Bؘ{֠<����I֪��N�/��jd����w�0�ш�������nmik��ٸ.��><{��%������jK���\�ESD��蓏��>�}x��i���g��z��� `��˩�=��������i._?���w�N�7��>�_��X?�;�#)J�-\��Vj>�����������)*:�`牉os� �z7��?M�Y��yB+1��}�^P�`ċUAT�p�(�si�j��!���~5hSL����p��k�X�'���nS����o������2���G2L:}�@L1����}��6�5#��Qj��X DwA<G����9���'��Z�����sכ]>C�w��S�d=9oޅ������{�V�+���w�Ƀ��E���4o��R�#���I;��E1�'R?����s�����Ơq+�m���dU���㯱6��D3)&�TU֞���j�h�vHR�[�Bݛ�tr���Qr��d`����P�^`��W�X{��hc�)�Qd�8������[`�դ��@n��	���G@5�b�h�Ѻ�9��軮M�͏������{����,��έ����k ���sZ�>� ��¬�wTSܦ����FX{�N,�.�F,ZeG$�eMO�������g_g�x�J0����}h6zP=�u��!������9��* �T�3@��3��k������ܢe�A�)��JX3/��8KD���܌��	��'U! �qE��Uy�O�Q��F:�Jc7�r�Y�t~�$�ZnWk��w���Y�G������\�������p��q;��·�k1�y�f8�����*z����쩿V�� {[�����>$`�!��g󝐈��6��w�^m�	�kd#�V�Ê-�X������"N����e���S8�*k�f�[��<��f�@����Z�Ä���^�y1-u���G�ź�����p����X=���52ZxS���V�P�h^�V�tA�U4��g���F���B�^��8��?�m��@�A�f�������(xd���i����uJMQh�����[`Mt0c% �	��Fa���P�g�����]��`�X�w���<%�ns!̛7�};����	
>/�Eߑ�f�4]$�,��vF�sj�N�&F���=�=/�.�"N�V�/��|Y����e� h��
��f�B��I�{D���
�)X� �Ư'K��,���A������)t)Ht}����A�ă��~����6E/���3 p-�[�K�����L@�!�-f� W�>7��������b���}6��q��xŉ�ۃ������~����@P��'
u��0�¡�R�0j׍�ɫqN:}/jq0��H�7�ir��nY#jX0�)v�vݽ��1��G0YQ���Yw�p��v��3��<0��9Q;���4����}�0Y��5�x�s��>�9Da5Lkm�ԙ���% 5�h���Y�_,%�U-�*�S�$�-Y�ȳ�������`* � ��@C/u�
}m6�6 Њ�L�]����y_�--�nb�6�*}�F$f	֩���p߹����#�5r� h�9B1`���PPJ�������D+�seRRm*��M�*��(@4|D���+u��3O}��!)hp���Z��v���8H�َ��iA����0�D^�7��rư�@Zʼt׍;�1�����h�F�cF ��z=��W��89�8^� j�[������y�1F�C�J�i�
s�5�§U]�-�������͗0}��W�]����mwեpæ�t�"�����ב�Zn���jr��ʐca�l�G�0ꊄ4��e���)P#��Ou�H�Wr{}���V	�]ͽ��*%L�����)�c�6�B���>���O��f�'� ��,�����p}O�A��uXx��<zП�_QL����7���y],��7P�`�8M-VE��J���%�'����j[�K\�8:���9
]��*\ZK-Ue���Ջ�dC�04,E4���*b�A�Bz���y(�M�J|_�_�Ba-fne�v��ƴa���J��*�ν��#�boY~iS��U#&��?�궭e3˰)ъ.,ǵ��$����>���UH����d� �ot�jH��@��+m}�ܙ�+���:�bk�k]��YS��E��R�Xf�֙�b}E�D�ܭ}2�5%z����*0���6h������e��%0Ԧ���{~dg�����?���o� 6g�Z��fmoSpK�@��W���,�������t��N^S��e����FHE_��JJ���B�y}	�� �)!h4䨃aF'��m�_�N��-��)�����鹅�޺uc�ы�x�ւ�G���v���Ȭ��0�Gh�� 0C�x��z\72Ғ�Q�'�ˇ�c=�̱`��_w6�k#��z����ϧD���1q�d��ڪ�%f,�l>˖��TR���Rm-�#�?�a�@P8f���1! ��w�8b�v�!�u	3FC�=kf)ZoiBXI�b^�Y�V���Dr!�Ɋ� �?��byh�)yE`/.[*���`�h]�
�O�d�zOn�8�ZTI+Iup��
��$���v��*���)���2o�������ݹ%���Zq_��*��-Q�9��Y�I�yK A��#|��G^ǽ��L�U�9���u� ^�x�h��ۣ��g�$/ �h���٬`�QÌ&/���H�2�{��l�>`8��f��5��-R�c�\]��p��'i=y?^�g>�	���3����P�Ƨ6�U��R[l��0K��%�(h��q�>���=~zN�u�(���dØo}/XG*��Y�tߒ���)=Dz��y����{���\��׬�]�sE��ȅAª��eRz�*_��bc�\��Q%�``&��Y<�U��=��\�Gϭ)Zi��}'+jЩU�\
@Z����pFc"��q?�*����D=��^�[r�d=ɱҠ �3�Jp$D��+����	�� U�t�Y���}"��py!��U���m�N�Ң��d�u#�׬��ꠢ�QT�b$��î�*���uV���q�@��Fʇ�q�q��R���S�EQy���|b��G��N��ym8���@�Q .@ѿ�l�����o<b8�nx��;�w��Y��ǫ������o_t>�����i#��!�CQ0�b�F+��6��4ݭ�t�"�⵺	�,g�r�Tۈ�|)�|��3�6�)� ���eE�Zo&���.�a=3$����b�,Q�4�E�d0`F�&��o��}|�H�hFf�D<�87���m�ô�O �cm\�_�}��_ -�Zvb�h��Ǥz�Lx��9�����6ͧ+����zt4�cM����KEo\�umі�/0i�����;
�|2������{�#�gA.�/2]A��'��Ն�P�)�sr�@L�ư�3ܘ�19>R��k��Y�a��,��)4�:#`��v-��/��CTIX%�K�Ҭ��T�@�`���[���~�)��B�4k��iܸ�:��8߱���%
6��~�j}~��KO�W4^q?��Z�Ά�9�5;5�����=]��XY��JB^��5����h�q52Da�����q&�5�5
c���|dM(:��{רa^|7b���AS_y��6����X,#]e��ɇXl0��)B\�xq:�{�)��"|�xi��';̍9��َ���z���E'~�p_������Q���O��'�d�9ܼ��6��"\ϸ:�Q�+�ܚs�¤����6�~f?gR8"É�ژ�����>}7��q��%
l�?�V�샯Yɯˠ@b��ڵ׻*���r�`@�N���Â.���}h��C+�/&Բ�Q�$�7BY�H���Ps��MI���؀�@��K�7A�M3��,ށF�E��wAo�nrЁ��|�dށRt�Z�vD{"���}g�y�:O���I�kz�YsSn�;��TR��]����X?�y�F�i�z�8�����zZ��1���r��ԡ�U��7U�֘2ds�*�/fh޴j��W�SsE�^��I~��m���d��KL�uHb���6�`�I�۹f	4�s�<��y��\�8����Y�~�xqT;�3O��F&�+ �B�XX�ѡ�@�ս���>����^������%�h �8gY�����F�i�@"0v�S44���v,X���L�P#LE(i����P+Z�[P��"`��m֎�_�c�M���*��$��/�O���hMq����Kk_�NkHx/(ace�8�o3�r�d=V�7��($�+�����0�;�HB�5T�����?-�7}_�J�JH����سw�9��C#B���Y����^�V��fm�z�!�,�Ԓ��,���@i��«�lW�s��m)7�-����N�2��[^N���S��,(��z'�Ƴ���V�	�&�p��2��r��X�k����{�~trr4p���~�k8�5�A����A3��N���z]�mr�{
�эc���>��,�g�Ff�x%?���zk����~]�<��fg&pv�{
����Q��g��;8X�t�L%���0��a��Gg|��P�^Ci���A��J?ԛwngT��$SZ���p=a���6�<��5�E�P-1�[�#WG��p��BQf�zf��5p��a��C<U�����O�1���ZԔq���B���y&�G����e`�j�b��݉�Lr��<�C��+��l��Z�˗v}J�8��gm�⢴F��"D�9����oܵ��Ģ��v��3������Va�	�1z�Jq�)�k%�����4��s\���ݜQ�rI�×E�"�3Pyt0SLP��E�9s��V^��(%А|G�X3%-�Y�zoU���~E+�����k����)�s�sU�QU�֮�'����������+esϙ"4�����J A1�߮����{���`�3��J������Ur�-��ֳ�P�A9�,�l��e��w��jA�C�6�̋�Xg����涗k|^�+�Е��ME.Nϋ-#/1�iY�hAYR��:�*@����ڮ����{R}m!q{��t�������0�E��q|��;���UˋW.��]�=b���K�w-�����ȑ?��7�l�O��*'��[IE��3;�ge�t�|]�+��΂}jc�Gi�\�&�L�P1���L9�a��څ�5��Wi���>n�s]N򣓫5�4`�ѿ����s"d�B��0G�_ཨq����Lp%�rɈǊ�s���ⷢ�?ɬ�e_5x>�v�T�I#BB$T� ��qk�ᓇ5o
,<�m�u�����������L�2�����9@��s�t��Y�4���� zS2|����L�<K���E�gWK%�vY)�=����t�^��4�ىk����Ҕ��!#����E�c�;����?F�xD��d]�s�y���W�l\>'V��^㇩6�Gx�&}FM���X
qqe8�Nv�1�j,��6��!��6s�Za�g/�s�ѝ;w������v�����ɦeZqn]�7�'����c��S��"����Ӥ��-B�4jWU���S(�F��v�%!͉��6[�6�]rc?�������v�)xB���Z:�xKx��p茑�JU�.�/	��D�fu̜y����	c��́�1��%:��-2�)t����CX*�!gU�B%�MmZ]���p�n
��(��SC����g�oL�:�T�V�|t�����JѺ��Rx���|h�Mn��>Gp k�Ş0O�1B��Ҷ{�OuF>K��#!6UF�3�ˀnMň�(`�>4�O��>+!������E����
�Y�!��_�~�Y��x5��ǪQhں�w�GHو�a�/�Fu]�8�}Q�����/uPv�ʭ�}��ٿL߲A�&)`�6����JbiT����~U�M�Cq���߻w�7�x�z��5X@���j��`f^Z���C�о���3���C��ITc���\ckh����|�0�q����ܬ��%J���֔pa�.�0"�S10W[1u,�D5��U����	��a���D�qO�%��B�)
.�1� H A4՜!�2��P�U)�d{���S��Q���ȾBOA�Ɉ�A1bM�0�b�׏�pH�֋q>��&:����"j�1�$�V�
FT tsӌi�9_K�������!�D�CC76�IQR%~�����&b�	�� ��ų�d�@���:�m�M�
��a���0h �{�K�D	�2��@�9�1���Zl������4$���¤u��x]���s����t��"���"��@I5^��z��g)Ѻ��v���t@�z�u�l�^��������r����s"s4�X��O�`��Ng5��*E5�r��0�֡8�~R#%7�B�2#v�r��R�Z�k��R҂���+�`S) �n�5a�mWz���(MB]7iZ�u�J�~��(��G�,<C}1OBge�)CxyQ��b�`p�N�ժ4?���ȢdE`�D���� Ѩ֛��yg�jv@kJ��s�"�-ÂcW#�}�;��(�:KBu�C�c�J�[���:C���¢+���\���7�c�i����"3�	����/F�M��b��ڶ���rV���AW�4���g}��#��g�g<k� Pj�LT��ܓ����!4����uέs����LI�v�y��8��,Yl�[���{�[�oլ��s�v��]�N��|��#d�U��ꚦTٯ�9�Jp�|�#tAQԤ�ݷYy����\C+�s�~�?�/@ﻮ�/��[?�\ �������zڵ��Zi��Ʉ槔�(ڑbm�g�u����u�!7b|{ML�.զ�k�EH�7�bJhoe���p���QT9�g�.��ܯ�N[�L&�AT��]n����-��i,�b�W�.��-�:�-?kri�%#��UѺ��X>1ڏ��A�y��G��5�zP��8�YO���i�>�܏`1!�5b8xԦ#Ì�M�!�!j�b�Q�gK���Od�b��gS����5F�X��������#�?d=� �Q!y�hU�z��*���;��A�R��gJ� �UVB�G�S�s�{���!s��6��I,=����D���F F[�u~�>ջ����oܡ/my�&!�Jߐ �����D���Fi�i�KNe��#�a��D�"��=۷���gw��}�%x�\ i�ܹ}:�ϟ�7�ݰ�3�8E ��E�SK�f�R��nkd��B��WY�������R�x��GL��E�t���03=IQ���T���@���<���\��k���F`�`��5�Θh��"K<�|�xZ��s���vű
��'�G���u���\MI�b���D>2Z�"L���"�l���|���s/2��}�d��6�_XѱN)�-��}-��|fʒa�d��5� *�5����S �J�S� ��:̅��W�z$Z)&�j`m�P�5G\|�kRY��E�G+�y���H����Z5��g<4�():�����^���oRC��� �E^3�B��L,����H��e~�;w�ez�gq�%Z�+������Y�4YE�bMF?e����P�O��b ������}�Qp�"��2��j�w�})�� |@F�i�V�yJyN�|2Pp�=.�l%
�q5�/�;(5�
<o���������7�|�'�j�t���F��փ�6;��䶘͓v��K�E ����ٛfH�@��>�+Ӝ�q�j����W׆(���p�y:8�hm�4�����ꫯF�
hsh�Q��/1֨���_Z��I@^�ہ�"�KKE�[#��d��0�B�;�cb�8݃���L���q}�����\ݷ(����E��#���"1�y�!F�o�#�?<�=��͈�X��N;����@�!���Pa��Ӥb�X��Eķ<]���i$���_��;���@/��~�(lu����5�L�3�^��}u��t�!�/����m�U����9����zO���Z/EU>|�0W��Z|���ܫ��X�+,��9_��sA/(,��|,���ۺ��G�J-�`-F冠��y���r��x�w���+�E �}��ݼY|3l�R���)�IVbx�������<L��'\�*L���肦�=cm); �j����,�,�d��%�.�#k<"'�4��#/G��;w(����~y��`AKL^W��_Z�0����e���櫯�@ݹ};� ۑ5CFa�Q0��p[�/��>=-�$��M�t8�|���jβ���(��ܭA��������\��$�E���'8�Sha�C�K� �2�)W|�\�Jఎ�F�p�tDk����Gߏ�
0s�Ƞe���`{�kX��&��/~�/�J�W{���	k�1��s��T�Hg���y�xXs�uy�;�7c�E� �s�oY �Q�X�.n�~U���>��H:eMt/	͙�u?�F�y/t_�H0=�������W毑���9�R�o�Y)��e&@�C�\[��ј�[�f墼C���*U�p�f>�Qa��F^�yfBv8wA"�I)�@���������ŝ��>~!��E ?XmW�ŗ�Y|���"sx�,�Q�*�mر\m�̒�<���Gv�f㨶h��ոVY��`]�!�9�+�e�O�YLU<��-�����L/DρA����С�����(kja��!�d��X�'�Q������ �D�\x-�_߁Q8+Մ�%,��u,Z?��i�D�>�2̒�ՠ�r\��]֍��!��B��׏45�΋��(�>$^c_�/�G|������X*�����/�s�/i����f&,>�s�J�]���s���:pm�s�+6��ڠ�#�魷޲�g%�u��	FE �k��h̲���D�4i�����k����ً����ʊ�q_����a�b�o]`�X�^�a��-і:�HM�C�Zh���h`MF8а������p�$�����7����F�ƽ�d�\�wf2��W���=�D1����t]q^���o^%���Y�����*��}D�ӈ���Mfjj(e�4��~�,��1P�aڲ|�:[��F���h����EB1*��CT:�C��jh�Ƌ��<Xd؈�ӈpS����65h�E�����#�PO�WF�	?^������#gs�o��ZT���;����\!��;{/���G��\�#S��(����5e����>�����9E8ڍ�C��д!�2@t�<����Ww$���b������`��蛀�F�׆���^lrG�	"�T�D�~��:�g��L��u�ϑFd�MU�����(�:2�YJ�o˼Aj8?v�,j��ڑ��Rbp3	���_y�Fӗ�I��}8>7�_ǵ
%ٻ�\�?�u�&Q	N��vPП߿u�e���k@~���������g/6�d�����OTg����r%~p��l,M8�1��Ku�[���͵b��8>�k0i�;=;�5%\�ܙY��"��|�2�ǌ�=W��(!C���a���h�e7#ͅ��R� ���?e��*aL5r��x5���;�BG��u'4�hy����<�$����{�:�OW�aN:�7�âe�ĵ`����_M��2�!�/=gSl?*?Q��(�)|Ƶb�@\o�C��Ѳ9+QT�(w{o��(:�e���%t"ĽD@��O,�}6�Ѐ��A�w�~�T@��8 ˨��ѽ���4�2��~9X<z�H���=��wӣ
�.�wƳ�����d�M�Ѿu���Q�v�e��<m�(��L���-��%Fӌ�`�:E S���%�1�˦�V������W�i�4,D�?���׏>���a6�D^թ�)�������Q%qYub�N�;���ð�})�k�t�^�+xY�^�y��L#(���Q��c��O�Zy�['�����˵ՙ;9YV�D*��`z���	�u���<X�f��a�=m�<�c=��j	�ڛ�U����i�9�a���D��{}�����p���[ϪC:��8��=g��j�:f���2C�Z�Ͻ���u����Bf�ȖWw�J��p��0���-S>�`�p4
��{A0��`�po�>�*΢s����#�U�IhFK�b�b`��������E�6&I��26V5�"�Y�4y=t�w��X(��=v�,j��4�8$<�i�y1��zM���bY}��Չ۫f�.]�*p��L�ys�b�՞èg����*}�L��$$]A�~c���S�j�`^gMF���IM	h$HP
�����ÃG��|���_ׅ����n���%�uU'⭒Oe�:�6�s�Dl�f���B���T��-�z��Ԇ�j�CԨ5"��Z�� ���+��MES�����թ��/f��͜��L�u6_\��#�˚P�!&�Zi��R��ϳV���G_>$��2����g�62��1*G�FnE%�q��T0��h��aLa�	cu�M�+��4M��\�i�Vb|�Ã]
D�k�x�R�,ZF�k�'||'�a:e.�FX�6��
��(��[�*�)�*&���F2��zF<W�ω2�g�� ׉���y���0>c̳kC%�,khk�ZP���V�:"@� h�����o���]�)�>FL�~K����������`�"�B0
�H�S��ϗ`�A���H�H��o�����=��y���?<�����ֳ��y��_�u{�grΆ?�(�r����G��{Y�0��ł��T�*c7��;�Ƥ�m�c9���9���6�B��'];��R81'm�zO�'����f�S���!*	�&z�h�w4\i8���"���{"�٨G�c�]��"S�Z%��F�z�ף�뇷1A�L��"C�Y ``6�I��Vd��`1O�����d��D˅�N�!Z�H�'AL�J�P�0Q��;2�H_�=W��x?b��1��.��y�(0�#1?+�ӗ�X4����퓯����(�&׏�?���3�%

��'� �_��3Vs'�t@s��q����u��K(�XV��=G�:��[���"5��)�KװW��H�u��g�Q�y�-]����*S��Ŭ�伓�£cl�� �ȸ�O7�?�N���ߺ{�?��?��@�ݸq�/�>�O���ENk攘��ˉa��Jy��Uƚ4׍8h�sx��ޜ9{b��&�$�/��u4]xV6���@�;1 B?cC/40r�&%-��kiDgĠ�%�'��5WU���D�Z+Z��`�ZHf���P1��rH���8���vc��Ys�Ͳ�Ht��"+>�R��5ph�{`�������(�٫�{�B$�\\��L?��̉ߣ�c�
���5���N��B��U�F�A��a��jܴV�fu8��7����wI�mF̙�}Vi {���Q��z��u�9#S�Qw��5֐�V$���������-枋(����,�l#+Qg��v�c�u��y�@��CV�W�u2�]�����^ؚ��ǘ�c^5�ud�p�� �c0K�+��[�%��)'��]{�����7õa������������曯�\.������z�<�\�|	#_ܗg�՝{�-`���^d��8m�~iR�J��U��HC(L�i��5��~b��\\Vm����p�~���p���YE꙱��>A� X��m�vx��S���gG�Uv0+�zL�[V���!�5�ǺT�HOzqn=��A+zqzfڑUR^��O8|J��26���<���(;�|
&0OϹ��5����pM�E�'�&A�Xp����kr8�vtpl̀�;:�a�g�=ZӺ�͂�����m�;o4�HM�F�:䧧��7�X�
��͸�Iy�|OJ
B�@ 	*/��ql��
���X�W�CJ�K������FI~�5�Y��LV{�u"a��Xz�������8 �d��1����������K4�	����>=�%���y/.O���}��X��hQ.����IrX_���-�^t3��Γ�h��ڗY��:���B�	�b��6Yo֖��}�U�2D�gMA�=��/:\Z����WI�cU0έN�^��h�k���T���'@�(��pU��}�2b�I-!��;�ˍU���(�w��L� �3�۹���wIIt��Zfv�=
���0n�E�;
�&!9Ns(�QPٹRE�a_���˔x~hg��˳�ݻ��~��O��8^� �x�w��e��O���*Z�kf���ф�V�������_�EJ�㞚�1��@[~_gF
�&�1��r�l��x��@��Jr�R/��8T�V���A���mi�L.T�vٍ!"�E�i���ߘ�����8I�#BUv��簃"�t?��|7�T�|"T��zp��\>}�Ԅ�ɭ��(9���p�-��N�������z�eXh��l}��v!9N�(��8��0ZB�k���<�ǅG�%q��>�&�$��R")�7Z��Y���~a�f�51�C�(�{3^#�R�����r�#��V���OMݹ}����gs��X�9|�ɣ��OcC�}��;Mܭ��`妺xV`8A]��vd��ڭ);��|�-2h"Z �t�Y$(G��0��G+�󦿩��}�!l�>P�bЏ����ǲS%�H�a����`�.�>�:��7!Qyd�%����u�aT�c�t���5N&�P��u?QI�G@�
�0���V��M�/�߿�Z��U ݾ}s}tt�d�ެ��M4Jj�c�g�>K�NPS��8��e��fa\Ng���b��,��3�R�ό(3�Ŷ����"��<���9��<G�4�{���q�&iL���	��&�n� �X�#$K�v�ĥ�UW �0�ޯg�*Ϊ��o+�B��q#fm�7�u���`��{@ʠ^��{��7MI�����K�:��Vgi]��}���"$��b�d����DFJ�軺F��9Î#MD��ԩ͵��+N` ����;<�¬��b@B�߲&:y~��J���D��'Z7�	h(����Drg��^��UO?���%���ް_��iZ�������zx�N��ޱ�S�w?�^�vՂZ��<�r�%�t��!.g����R���v�p��A�_�b�wS�y��N�ޣ��Hz��};��tm���M~�^�S�{S��i����M��X�)�4�-�f��u�6SBQ�l}���M�m��b���A�[�-��?����]tr���Ν{�x����?D��(��1����FL��z���ט:q�} �Ǖ|�A���+L�v�h31��(�U8Fq���hS�"�/V�*@,�O=r�	Nm]��bf5.�X,JW<��k j�Z�(2ƚ�� i�0,�&��.+F�F��ƭ7��o<���g�V�9���&�to	$���8^>n0�5x�y?�� ǩ�m����rr�kD�_�g�U�3���G��)-�KU4
�?����O�[�U�7ZxXC1�&
W^C��/�Y����h�@|̇`�Áv����j�>������Ձ�*O�xtܳƤO�of�I���?����������c@�V�niHН�n��GqVAp��l��;����v��v��λ��H�����{� :}&&��}����1��	KHkBu����7zNo���L�LE٫�%�r�"���'i��P:@�"�F�$�Lo��4�cݤ�	�6���E��
�7����������_���?�݅���=���Ͼ���'��]��C��������`�����8��}�lT�s6Aj��G� b��g�kp�#�sB][���{7���K�a)Eã��E��X�{դu+��R�#:�5<���Fe��2�䀏4��l}�fhƘ
���c������k�����=���O��(�7�?�~���J�?����}���]��\�>&�RM6�t|��g0\,�����sӀ�{
����=� m��0�C)���(�+Bs|�aȣQ�n��a'>���\c�����*����M�0�s�y�쩵�s�z�7��`��_�u�d�+�B�K���{dp����
ꕇ3�����7!s6�Ӂ9�,�)���e��Ԁ����ϋ����B!��=�d�7�V�(9gEy#�k)ZG�i|HX�D��6�,TJ�A	{v�7�\�ٸ7�s��P&ὬYTv�zG���)��{��֐�g9�(������������k�U �����_������||2,���p'0 ������H0�a�.�+�sj�2��7Վ-�-T~�nTJ���c-c\U!j,˺t��5Y�ߟ={V�{���~��`��I�u"�m´.2��z/�@�'��P���cڛ0�a?h�,�헿��}�����i�%E�x���?��?���?��?������|� ��$�2ZV�����/�ʚs��BԀ��u0!��
�z�Υ��W�6�54�q.���Y)���&�y3���E��4���K����<��x�y��?�~u���A�=�~���>�����\l�0O��"?�Wܷ�y���~�;Փo�U��O}��Դm��U:kV�x��m�Uw);
l�}V�s��_fޔF|�0c`�=��h�$&��B#D��}|��.4W�^��Y=��	E�UE�Ζ��$����gP�b��mƽį�M#[#O��r��B��g�&�k����������E���k@�{yx����r}9<�Ic����阬4�s� M�����ò��v8����C|�:���p�+�FM�M���$���׆�m�Gk�����inr�����P����b �Le�h[,&��jK�iR���1��\���Qr�C���c�Ƹ�&�3�-�ŏf��V� ؛�����_�޼��;��˗i]��|�8GJݺ�/�>����V?,#�/���/���A���{#�����[�u!�8��
�_���>,��a��`8q����!��r��o�46��:͖�����pM�ڰ���	V�?=�]�3{����G���3��է�~Z=z��z��E����~�u��� =�����:yn�)>�@a�7az:(7n��g�{�S>�B�DS��g�5*&�p����E�7@J��1H�:��U���s�Έ�$�Y��(�׊�ט/�ֿ�0��*�?u����OX��g<��g��h��O��3V���c�7���(��kQ�dP{v���_>���� ������=hP�|x�0Q�+NDpv�ω��2E���Ņ���skă_G���.I�z�6�Vrՙ؎H�P�g�C4�{��5qb�����}�O>��4u��lLx팉{��2^[�����<"�0�v"�d-q�&���ώg�HV�����4�	�ӿN��k�|�I���}��TV�|G�����AhKp˗��K�&[���xt��)�Z�	��y�D%�=�k6�!�-j�V}"�׉�Z�q�cRa�O��[��"�ʼ�P������Zy�w�y�����?���g?5ea;���鹅��7���o�%/9cq�������8��|ǅ�g����~�Y��ѱѤܯ�O]k;��0��r#�%�RϠyn��YU�XA$Ѐ�@@j�&]NQp8?�#ܛ��!��t�'�J�ΔjE���E�z�>h�j�©2��!�Hk(Y�\s���Z
d���"���	U6]�}���o�Տ���k�] c��o���������w"�{�Smf�ɍ##t�S6�˼0Ҝ<x`X��5��0^�lɗ�����%�41S��tڴ�j�����gM+�]��`tPC^���4�/ά����^�%��g�eA�u�"D���T�M�j\OL��h����莚��6%�A���*�^zAF�v4����g�L_��W�m>��}��t@�1l�զ���lX߿������}���x��]{~�_[��4��İ[��U�J80u������b���`��p���D�{>E�F`�0y�ͽ� }q��ak�ᔏ�'*2�]�-ae��!Iy*HQV�n���'VC�>����7���E:Z�M�5���|3�Yd]/A�������=	��P�:G&�ЗJP�0���8�!�?��s�o�H,΋~O�u�@�@e}'F�B�1�:Fb�h���K��&��@XZ|W�]�J����G�7�}�_�|�RA;F�
��*�Q���b�-4�G��6������ZLk�~��ٗ?���u=��_�x���@��_<�-?J�sJ�2�8D��o�F�hXE�����:�F�[�F�󈊶���3_���f�/3��`j�	���"z9�-GgV���{��g�3-�wI������Ц���5+Ӧ��U�rHk��7<�^,V�����å��g?���V�A���p��A%_УO?��%!�g�54?>����A�#�P!�=�uAOp��C�U�u���q�x>�lt�# cpT��'4�a֠�F	#�Fc�߇���,Q��k�k�o����_V_|���ǟT��j��B�T�j`�JR��(9R�����url~	��?��zgP������ŋg���Rr˞5u`m�Aǀ��G�t?ѝ�ۃ��g�"��6������� $�4+^emXW^ӹ�P~FG���P�R߅Q�s�i������3�h#���"Br>R���\�?�X��O��t�X��$gw������������۰�����;[�z��ᡕ�s�C��@%j������h4'�}^ڱ���%�и�*��1nQ�T��j�	�M��M	q��9[l�Ao-�R���S(&A��^d��ri>��vv��%{�t����҆;B-��������1PAh���ߺU:��m��F�btii�?d�5�w��޳�޾ck��<~��U����쾊F�6i�6/<�\9Bj�e�$��V� �1�Ah?K�,�!L2j��$O �0$���烏CǼ�H��p¦����^�(�ݸ�#����FgE�0�"aŘpj�Ժ�h��9t����l9���c�?��z:h�BTIz��[E�'_�"8�}�e��<���@���j��{���AOϟ>�����X�AV�B���E;i�V6YوLR֒���N����m6���b`�P�Y�T�8��*-7��$���Ơ��*��9�V���.�9z�(�D.bEe�g@�I�g�s*��?�$��(^���UXo�����;��<x���-�ߊ z��''G?���t��Vg��X^a>z�B�EI�*���ͻ���"��J
6�2����}�4ڒJ�К@A�,�`9�o66�D5)$Ra���,¶h�f���@�	�2-�1��.'�(FmE��(Q�����i�g:8���Z�'_}m>�w|�����4=A*rk��<{��n��ڭ���kI8i������S62ਁ�}"�k����h�8Z�hEE����È~���o����(�Z5b���S݌�+��G�aC���zا��bl��|<Ϟ{`�Ф��*�����ʄ�, �!X��Y�I//#�m�̴���sCa�Zя�Tg� ����(P-����z��fY۴��Y.Z��F�
��haFX��UI����7�O������E�f��^y�[�y���<Q�AR������|1�������~�����'��������������a����{��/!�Y�{E�Ű雽5�C:�	�V:�S�=�٪�&�*�����i�;\��}'kP�w��������@\�:�E�jF���F��*��]Y>��`��:`��϶#��jI%':Nz~� �,'��#+���i��Z ���Kϩ��=���ž�z���9����ܢ����o�=��wM�����\	̋�y��v+�N�>Wu�����FK��<�F(@�O�i#�{!+U�5\�/F�vt�� ����6�J޳�O�[����<��*�g��_��IGH	�^�yb�ž��`1��~��`SY������1ŧ�����WY�7����[�J��v����(+EQ����Q{w��,A,�Y�Gɲ����ÒYs��aN~�"w����D�S��0�9iEI�>Kjo`�ߥ�~ݦ����j%Ȉ�)�y���zDe&��}Ys�4,�1��n����'~��O������aA�����'���G����lX��0����g \Љh��5�O�Qj��ϳz܍sb�\��AÍf+��Û4�z�\���������*xb��M��&�@�zAѼΖGS����!<4�QD[���p�>w��]�?=M0飿�u������oTO�����/���?�o�2NC!���t]=���4EWݿs�zqv�{'�zB��`����Y-��c�pp/E�Q�(:�5����#���sd�� �E?
	|\S:��e��z��a?�5�`�"Ø�y���aG��3N-��>���m��poW�%K1i}����`�2�����Y!�PT+Nʖ*��j��Y���a���V0�?C���Y�I�����?�}���ū�R�4>c0�Vg���P,��A�Y�Lt_�"���G|���"�î��~E��?���dU֢D�]m�*�~ ?��8��z>
�$����/�z�����k�~�oE i�����
:�i�n���nW�k��9���x4�*��c7�]�5��0H?Ҏ4�/��J�HL[��}2��>���i�	�p��*3"�K�P:��9�!h�1����u"tTڄ�����g�g�A	m>�N�G��'�����0M7@Q���?�>��_��+���k��%�'j��~,�UBF>"E��p��58�"]�K��/�V7mF�f�>�#�X_��;Z0�e��]�S���뱀h�Aa�����0"��h�#h&�H�"���-0H#Z��s`�*�n����\�<��{�ۮ�Nl�s�Xs���q�hQ� K�,���"��YC�1`�Ǡ� �S #A�� n ��ĉ�n�h���v�-7d9-�e���e��8H��z5�����[k��^�H���{�&�U���s�����ZD��յ�pǹ�a:���s�5Ϝ9.^�C�A���r^�4�׏��|Ch�l>���uO4�_��v'����\��ךuD~�����Q�R����|�\!ÐlKN�%�� ��N�DϲZ"2�.��������W>���@!�TT�$_��)�t������YD��X���b�������k��h�e
��G?��� @���_��>U�����h���r��pi�%�jgf������&ϕ��H�"���dhM�}t�j�ԝ��Y��T�Ch�{d�f��W��WBї�׸�c):[__��cq!�ǆ�H!	��� m�q��{x��`�����0(�j����#��h2Էm�v<���v����
���B>O-"���M���[���{.|��ߐ{ێ��ȱ䵮��w�uW���U%��$�ʈ?ln���l�<V��@x
H*X�Pd�Ϟ��8�X@/m`���&������I��0+a�$r���9��C��D�Q���`�8⡡��/8�G�{�̍�r�,����'�y?>��g��J�K|`���^4�M���+�.�tT6��~>�ǵ:�Om�y��+�U���Tm9T��_\���w4�յ~A�=ZE��5�K�J0
����a`��_������D;	b�!6H����[��:�����p�VV��%��$�5�DP�;�m%
^J�k��\�3�L����5���=�#ꛁ�s��S~O1$����q)F6�_�����\<��w���4YY[�|��w_yꩧ޼���)�81�������\��R��Gۦ��z+[p�%��gw_(�� @�sx4��Q�UU"��޴�|�P=p�C&�Ͳ�²��m)�!*T���X�$_A�����@B�5�%S�
a�
,Rz�D�2��Eޅr��k�Dj�:����{p�9��7���Z��΍�P�g�x�j}�˯�a2�i?�J��^�?�n�F�_YI�m,��(lJ�*�M� ��1ߑ����=�J�2�S�U��w����p�ׅa�Vq�h,l�6��~YX ��}������6�@��@�H������xr�	��4�xckS�� �| =	�E��iժ�I.)��rq�w��9O��X(D���CI�� ��#�f^��$�Q��Ƒ����:"	�N�{�B�7בk a�/zqݮr$�CKa�"{׫�9)�^F�7X+*���������L~���?x!��g�|�Z�?�a7�wD(M���|��P����3��e=��gx�A��F)�� ��{�{��x||ha����@���f�F x�/h�hNb�dCq��܉�q�!2R�GUi����K��S����PDU��g2 -��,d�^_]]��ù�-��itO���CiSq����:��=:��D	���C�9���l�I]��j�=>c7*�^�N/�}t�E�]:m�Bȼ�l�Na�m1��kEv��A0YG��(�s��n`�">���sK�!��(��lZ���g�\�����8�2�q��KG�3�}!��(�N�����d��M�*ĝ�b!�p<�0x��@	�	
D�	�m°$�ߗ��8����C����F��H\W
�UJ6��M�����}>���i2�B�P�}8Da΀Q�E�@����#L��9�U ���ņ��hE�y�4K��a_�Z�BAs)�U��6�4�׳P"ɁR�M����tA6Z�@%��	��i��kӯ�/��Y��ҕ+W$i��G�.\8's�|�f�����9*�/�
(t�ۈ?�v��eJ� ��!��a� ��`z >��.��\
��g�}@�b10?�26a��4��ha�{c8�a�c�zh��YB]��y(������#���P{ptΝ;=�51,`lG%ث�	�Z�6V%Է�w�>��d8��l�q�:��4b��J��X�z��E��;�*߱x�BS*��ؼܱ�'A���ɜ�%��!�T����z@�q�[�ssC��ϒ����$�!������PkQ")8�����h��M���x��m���;6��zis�e2��6��>a�]�������o�E`B�^_q�xX\���z:��w��x�'�7��������4^��ݺwb�,^=��J����D0�?H�c����nkA��
����.�����M����rb/�U�V��"�!�K�d"�r�"������)t��Q�m���R�ZZ�jW-�Ȉ5�[�
�y*������vil��3�`�,�	�J�/�X�EFh������X�$)�}�x���-�A��$�v�|�g���8
����΍���k�f��BX�;悾^8�4�>+f�s=:�V���S��1�F���� ��Yq^"��by zv֨����#�±*�$
��%��	�� Zѣ�|��*ސ��26(��|"��2���"B��!�Ϝ�;Q��F#�����3a��U��^O�мa5�����}־3�X���sU�� �=zb��E(�Ѻ/:��ĺ�p�t .ȹ���QV �D3�L����rn�֩%$�k�_U�)�*�sh4 l������Y�=������#��aC� -��h	dK���J�q�|��pk����yᚦu���^U��{F����{�=�0��&�Ҍ�:�J��w�q珞x����o~��
���|�~�7n�>������r@�f+�Ks<7���ztt �0��f`�D�?#ۊ"/�G��8:F���Z�gI�yk�[j��YB3i|�¼�2�r�J�[h(�� P`���6r=\Xis��a����nd�F�x�����ׄ��lԐ{���Y�IyR�Iun�ÅZu=(;˩��D�� *8�&�y�q��ŨFpI��R��a�7?��ڪ:�9�6
(M��;U*�����A�/l(�O
T*%|&sK(��8Ęg�m�1YK�BH�GI&OO�'o׆ eh�#�z�V+��G�1GE���d�9�3|�*��{@Z,yB#�%cƏ~����������%���^��gC�3��U�C�=$���z��G����cEB^P+����,���b����O(|FZrOآ�̞��{���hR�C6╫W�y���%����K����3^�4,��(�XT�i.
W�aY�1;����/�-���a�^N�oސ��Nf��Pv잺�F�/��J�{Euu��{�g'���-U@����w��ݯM?'���)��Sj��ԅ��3������-MA���Hh�7��G�(}z+�T��q� Fϐ�"\�Ŗ�RMO�:6��XbA7!�%^���p{��@�����\����b��ڟU礣Y��;Y7��O�-��Q�i�I���O�׮�}J��_B�\Kx� ��|
����S�q!�doI|�V�y%���QB4�o�ܕ0����Օu�����w\��.�\ؘ��x��$�bV{p�>**Z�	уe����{I�u��X��a��2�u�X,0��x�sNTT�>�l'��|݇G���C2n����C5|N������p�P ���WQ�����8_+���/������5��2��/��6O��jT>���Q��:=Q<�^�2ix'FLo(�	�g�J�8{e�2���>�r�DO7�b~dB�JJ^?�I�-��;�%�?c �Ytq�"����%�=9�<�
p�_�����6��(`�V�W�J�-U�k�N�)�L*�`_ʦ 8#�'�`�̣�0~�.J�F�X��4�d<�z���o�u�]o���-W@�����[��/~so�Ţӽa%��b%�.w$�0�$1�P����TϋƟ��;���_D�\�4JU@���VF7�no	I������ƖBT �z�d�"�M�$<!
(�ֈ���bӹ��|ldX��{JH�A�.$N/�EW���"Sq��ō>����*��̻Т���q��� ������mBm����t��n����4���	q�A��璮����fQ�6�L�#�yI��9hA�0a���	C��������po��9��L�Xfc�2����&�p�p���5,��y,�V����C��Pt\C��)�B	�!���OK��E.ݕkW%߸}�� ��8��z>��w���°�M�q�b�*5
z�yG� �G�׋���Qc�0�(�b{6���&��RA�ɰދ��#l�Ƥ*kx����Po�9�9��&A'C�܋����r�qz^ C�+�/	}��NX�*�5� ��{�I�H%[VJIc�l�f���B�[�#C�� U���ht���3/~�#y�+ ���Ϳ��׮\��|����{�z��0lnm�2���P�����H{�w{�j���M\Vnch��݇r�y�G�--�Ƙ��FRz�a���	:�� ,V�/��y�&'*�n�,�2��b�<,R�����;pڠ��B��h~��sO#®�{��5�pm��!+��n1�����"��G�{x a*)n��/�#lH������]�X���s�gP�_�!��u��W�cd�|��J>��:sY���&�u��^�G� ����?�d�����=��>kM<\��D���fc"�BQ92�D��sR\W泐ρu|��u�
 ��_(DA��C�7���=s^����yK�j-�ʲ\�)!oO3mL�{L;ׯ�BD8
f;*3Q"++���<�,��j�f���S4W׊Y��� :T) ��{B�����t���1��Lϗy�o~�\r��&���8Y��5z!)�h��|�h�ϕqJ��x=,(6�%(r�i��F`� jHH�r[�!;�@xq��^|��Go��a��
���:��w��k���y�V��F��FRf8L��&8jgD�}�� ||\7���$Ρ�6^�*������<���+��%��a��tKT�V�D�P�;�]x��������IͲ�M��Z�0�{�.4q���$u>�)R`�C<W�y2F8-!�bm��@�x���p�s#%豎�<�%!��p E����ԏ�yV�Sq2�ؾo�@������<�R����M������(�1(0��g���o�����:����s���+�a���V��sg�!�J�}�7���%E#<~����ŋw�����<P�Ws�x��QP�(�����ÙM̠����h��� ���ѾX�N[̗�W���)��ì<_)�r�����?Tm�'��p=���Ԑ^8=�
����ģWkei�	��\��٫R�{���"�����Y�^����3"y�x���I<����x/I{��ۍK�\;w��W����{�mo�z��|��|����hq�'i�BE���q#$�Y�����4���ܙ3�9��
�,��y�j�77�X�E'YP@���f�Gh�a&�l$XŋYԉ�C:v�I؋g%y�&%�{�N���JhŬ?Ƴi�P(Vu�½�f���� L�(Բ�]<)�&ǹNF*�_](����P~Gaǜ�oU �,_��E���(5����n 8X���R�g���UH��y�N����ٮ��t�6{&���2Y���s�Q��в?���'�1Hc��3�@�Ϡ�`b�?#<G�G�a3F*(zYޣa�ʆ�=_��g�g��z�`�~BQ mN�:+����څu�٤J0簐;�'/g"Z�0v�����յTi����[#^�N��A�$�����^8 ؚ˙�����у�I�4x��A�p0�\�6�n$_jQ����.k!
P����d�,2�W24��^�X���|0L�nd�6Q>��Ea����n]Z�ï�7�\�`�L�(6����¦���}(����$�l	��A���x���V��8�'����>w�����l�xٶ�BSr��y8&���%b 5�q��Q���7��Ef-�ͺ���X�6͓k��Q
 	؆�"�ѬX���bQ�U ���Ӄ�e/���>Ơ� ��aX�����,d�0o�|�������4�Do�sƹ���T,_i���@��@��
�s�	Ŋ)~��
Uz <���SQ��)�Z���J�^a��l�pp�������'�k�ŽF�}�2f�
���c��N��-�f)O�g`�+s '=^D�C�<%���vx���"q=|>�>G��0̛���` !p�s}٨�T�x2�0����x�E�y�P�Yu���9R�5�8E���98\��g(���(���eQ'{�q+k��BVzb��CnJ�	�|i-���m2&��%����Y�v�p��{��Gk�k�<�v=�+�w�Y��������uKu��E���?����0��q�=����w���w��?X�����:���jP�T8@���RZl0'oE���ň��N��H�As�T�=j�쿲PA�JS�*Œ��������O��/��^T&3�y�$�V�$�>vے��V�Hي��VY?>S?�.�`�A����F)�+���z�0#��:/���i:U��b����@�}���߽ M5'��+���ݨ���콬��6�d�+���
E������ST�w*�����
a%���l
RU.Bh�FscX-�y@S�B.4���]����_�]H5{�\@��$A,��M3T�k��0�WF�p�����zT���p�� �g�U�+o80�I����CL��e��U@��A�����Z�)Tؕ����R@��S[����D�����#�C�JY�޳�8�9R��r,���(ŀϨR�cc.�5��)�H܄��/�J���(thEh��{	�3�ćT��Y��o�c��9]ʔ���������<(�mM��t�������u22�lK�#�n��y�tz�!��w���}�c��mo���������>'��qҷ$�[�S���uڤ�f~�'���X)�~�d���ns+�a��e�!�"~>y����f�]*p󖓆:���lO�"�R��W��XXs�A�#�	Tg<X}���I"8%��%!�C[��jMHy�F�5�T��</�^F̼S+�K�B���|�_�D�I���Q�qk�JA��	>ׁuJ����0s<�	�u�����q�p�B��k^�d��9�̛��|X�#�&�ψArT|n��(�V86�{l�O�JO���=4�>��=�"L���5�ߗ_{-�d-��P,*���j`���3�2.�%É뀿����zV�� ����T%���*���	O�2ol��?\/kҙ<��~s\�~�k��^��=/w�g�
�rA�B�N&��l+���!^�A�PE�F���w�롗4D{��ۦ�0.]�o����l=�?-�-��L#i���M�ʃ����h��ڜR�x4��<��6Z3D^%�}FLq��A(�� H�����ȣ�ru�R��l2
�RC�WU(�F��L��!�)�3~�&h��Q�E��"�b#�?8'���b��8��E��CU�$Ě�� >>Ε����,�C
B�h3J�}�b�)!_uaC�&4@�^�0���hW��UIr��<��n�>+a����E�M9�$ޤ���4KD����J�+���Pz^���Wd�B�y>�H��0?��LË`�Ǉ��,��^XѨ����8�ą���Fñ(.D�H���({chð��Xر�]j�o�h�łx8ÁB��ު}I����<uZ�9^l%�1@����;k>�������-w��g!�/���ؕ�@/���¹�?O�m1Q)�#��£�<Z�>ߣj#�L}Z �7�	��]�"�chDEe���%����u��&�j�>�(R���5A]�x1��%Jk�aQ�^=w��_>��#��mo�z����~�?st�����#�>s�������t��A1��u�����!P\.Gţ���[ush�<$������ �M1d�
�n��8�&R�'�`E�A���u�/r�Φ�H2�Ja��Q�l�Dd������Y�!���'���g�ߋ2�0@�H+Z�� �h x��oISȢ�Ic�Jyn��pfIN��d��~c��JT�LQ0�0M��ʥ��C!�Mt�ރ���"a���<��d8����|[g����Z\�2�=2H�E�ݨ�[�{�w�5UP�zB�Q(�Yy]*/���{p��Hü��9w6����'�aV���!��BgΜ�5�$D�d�|~$���-��^<�ԄA�S�յ��9��0CF�;�/Q��w��L�CQTB@FFw�P)zClM�ϴgX���l(�\sp�?e��]Ys�1�B1��7�1�/-�#�W�mzΠ@�|M/��@&�D�)��a����u�=���G>��_j�?����٧w���&u{�s�2��հ���c���V�g��m���'\~x%��ˊ�������r���r˄�6p_���6f�d��J n�n\~@CYEX�*am,B��&h�� h���@�3O.4>B���AJ��!�����!�JE��B���\<<���!��C��Q�2<@V 
T�����������\�kP�:^�)���I�[;*��εի�2���åT�|.��ǐy����Q�sB�jT��c��i��KJ�!����|P��M��h��}�$�x��_�Ř[��_�b�����x�ThTj�z�A������Hs#���W�� �F_�<�-��\�mG:@���J	6��7�֢�n�i�j���kR�=�D���|�-�Rms3>9�'j��;B��J<+�5�5a����X��W���;,�wn�J:Z"�J���~h�e�@�gY~T��3w�ߖ�y���,������2�H�����:)�\A��F((�+蒢��������jQ9��6��Ua��O>����˯_y�ɲnOG׻� Aha�����wE�	s��ёP;>�1�ۤ�D����° f�+�(z�T-��K��PM�k�P� i��o�zk�V2���4�H�:"���P ��ǡ�N�)�! ���`�k_�����2�mV�{�v�7��_�� ��;˭R͚�4�y%�>\I´��L�"�'��I8�a��&�D�����0������ҳ 3�U޵��F���/���X%�8�uh���V|#�����X��\o�
� ���e�᳈��$
BZﴰ�%E���N̾F��i<��i-	���uO�F%E(��d��0}��E�H�S�4j<~O0�xS`��F���0��'��=��h26�*���t=X?�"�5:VP�|6]ʓ���{!8���8�θ��1���֢i*Y�����ؙ�߱�v����(-@����L�:ԁ��r�5�
u�׫R�oQ�}����/R�.�D�9T`
�V)��:��f�X�C)1����������p��[�x��o�z�᧎���~���7o�p>_���nՓ�Rc��Y��|7�L���l�G�p<���M�ɔ+_����P��J����$�t�$�tG���)^�1�B�>�*���>8�B1�Xa�]�Z�a�hAc���g0�j���TeB7Y,��ڃ�Q|�(�*0}F�>����TP ��88>
���*��ġ�tѧ���fQX�AhTQ$��fǶdZ�9��v�Bѕ�ps<G��D��Y�2�
K��B�x_���y���C ��c,N(/�
���|RC�A��l�PI�qx
U\o0T����H j��m����k�l�xNz	j�
�M����Ⳡ��k��"r��3�?s	�ȼ�/x�,��� \04Gԑp'�L�zI?��� Cy�ݝ��~�:C����xb!9��iEdJ�@���X�G��A������ %�0�@ٗ����1�� ���{C)���?�h��̹���!����~�{�Ma�|u2Ik�"0���ܾA)sp�pۧ��.Ʉ8�8c���c��9�\	eM|?�C����c���N��V�O�)�RhDA�b!X$e.hM���\������H��F�3Esf��I�0R�|R��=uJ�Hv��ё�0^�_��Q0��`F��b��(c�N��;�����z�-m��f�mW@w�{������O��ᇎ��@�"�X�0�-C0G�����=�ð��
�VZy�%�AU_Rc��x?n��岕!�.�;4$<?d3X�_=+ݨ��$֬a;���S7��h"�4S
]{eT����⁑���������γLa!F�7���m����Z���� q��@��*˱�w�H	n�[������7�00�Thũ2�:X���=B�[��*%s�<ui¿JE��8��l(�.���\{Qe�R�l3��XT^�\��]Q��=P~&=z2���B+��2b�.�|��H�m�M!���H<�����Q�r]Y�%y��,�G�����k�	����F��ܶR����5j-��n,�G��Ϗ��Ӡ��PX5��2D')r?\���a��']�_�i�Em�D���Z:Ը+��+�Z�t:dD����C����L�>����3A�V��õ�ĦBY�C�����(����~�m�^�qK(���vO�9��Q��\�̋q���R�v��'��m�A�s�Ԋ�y�R�Im�b���/Xm�IpZx-F�Ԛ�Dt.,O�	S`��I(�rwL��>*UM࠯
KV�T?B�޷Xhnt=́��7i��w�,#ټ�b��2,�S�+߱��Ƭo|Qs��Y4�I/�9
Oߣ����X�7)�T���.}>`�|�i��R=�T*{,䕨�u��Kir�*Є<�e��&��4�a�"�VO�sD��5�)�OT�ͦvLr�}����`!,�=� �*�#�A��ZSɆ�e	3-t}F֢�j��kQq�W	��9A/� 8��	A+�nV0���!��'J*��T��0�1w|�z�Z�n*��~�\�p4Hv���{�R��R�F�t:J�*� r�lIP��.ݒ�Z�|8[��5{T�"*g7k��PA>�	�VYN���v
� ������\_��cၳt�
���Z8{�t��{j�,4_�c���ht�z�[��������%z�����o~�[��v;��&	�
���IK(��$� ����Eu��!�i.hJ�%B���p�V���Bq�q��P�͌\�t�yvH��A�됒�ZQZmc����i�×-<��yZ�rHgY=���=,��2�V<Z��L'���!���)�/�A�@r{]'0\$����w�J�J�[�^pQ�z���T>�F�	cuu�\�"�%}���z���T̃�sy@�E�т'�*z �\��6����'���!~qo�FZ��˟�F���yJ&T+��P����GR�c((*]ϐ�� K��?{��CT�~���2���e��Kw�6Om�W/_e�������<�g��V���e����+�?Q½�і�=Ū��! ,Nѳ��N	���}.���$"y��}��J)�ڕ�[n<��mz��E�Q��L�#�|/�?(2Zл䞁�rY�5Ab��#ĸ�wp����z����m��¸���w�/���ǳ�G��陸�{U��\Hi'=��y.L_�"�¹3��J��2?.�ظ��v��&����@�H ��«Ul���쫌�Q��~F�|�{hs����z6}GT,#��v$�>�&R��S�/$i}ѣo�������ކ�esS��Q��k	�Z�'q�F��4��:=�˳-�Ѳ�����k�s�$>��B���Poͭ,���C���ZȴH\cyR�!�<�J��-�*�|�sH�a-�D��Y�ֲ�ZT�I��4=v-���$��w5�G%%��oo7�!�x6�����P�o-��&!*,�CX��������s�hH��\+
T����A=^|�y��⳼���⍞9{N��e�C�12�j�E:ɋ!1���?2@�p�,��&D�����P�sRѐnG�BZ�s�Ffk��B"$��O/�S~e�/:�^|�瓅�������_Y��ap�y�A<��#����J�7~ј�g{���}����~��oy㹿o�2
��'�����/~w�;qg<8�΂-�!l�͵�0����Ia2x GG��¹B���,w
<��i�P�>��0�
֎hcU7iw�ܱ2��m�:�}!�D��2tR��rJ#��jou)�Hf��n�UV(�Bݼj�Y0����G�� Ef����I�Bm.������y>;F�»5�k4o�y��?���壗ފD<<�`����ϤR�����!��0|C?WT=��y/�����Y۴`�^�����P�%����1�C��j��~�R���$O^���s�w���� P=3�� ��Jy稄t.���{�����=�H��d�D�LK���6����7�O��W�=��{M�b޵�s��7E��a�{?�������h���x�x?�=hA�:V<�����N�|�x�1�������>����%�"�Q@?���=��~#��5gU �@o�E���ŀ�6`���R ��dٌmx\��b��&���L�U Vt
�4T���K	��kܵ6!��b*z@ ?H��Y-j����ت��8p���;
�G9\�������4��a��Z14THM����G�h�`(9<��R�0�vz
)H+R	ZM��Y��29�Ee��Ul��E��ˡ��N�K�v� �,^�:x�We3�%/ǜ��+����ŢQ����W������و��/J$�`mVdWe'�����Q���Gù��ϣ���Q!-�u+%��s^a�K�b���%��+i~>��=:�k5K��2l<��܅�aې{�����q'�s��s��u �P���k�>(:*E��)�N?
8[�wE���9���BM-�H��>H,R�F(B�(��yYBReÕU�J��P
�а:�9���r� �9��h��P����y�Y���ȹ��@D� EK��Ӳ*��{{?��������m#}�qK)������~�k�G�w⁺3n�����4�Q1�E�7�̓�>(��;"�:�>��"s��[�����&� 9Ɩ��y<Mqb�~�A�YUs��)�2��@�F��[����:���]�I�����Ov�J�!�s�>6)�6Q����1�A!@j�=r�ڵ��|�s7|N����1|΁ʻL	qS��(%C�D;][c��Y�d�f���e�*��c`c;�3�s�S�{��?�s�G��L����,p���fB�V7	!�'k�����3|����u%��aN�:�ד���^�y�QȆ�#�Աh�<�
�m�������rq��h�c����.�ί=*x-Н��.�N����s-��2��ZA�}���V�A�Tz�^�ӫ����m)���:޼I�%�.ᨁ$E�����#�D	���<�݇>��go%��R@~��_��/�ٗ�<^u�M��G�������pc�9�Vjl��\�G�` V���~�}:<B�
@�J�J�l�����HWN�U��w:Uk9Ą���� 	��G��yϥ�����ia�TXHE��a��6bB�b���.6(���s���x@��bHH���&�9�ᔜ��SH	٪S9��L��=Zc^H�(P�}���'
7�V$��D:j�5���t)_��&�����5I^Yi�j�$���ai�<d��&$��1��ډ	��z!�Fu_ez}�r�I�D��������ӡb�ep���0�$/"�o���|;ݾX�$�d�յk7©3���Ф\���*�%�B�1���і�Ƣ\��SUf�
���d�@��,�y�=C*�����̢@���
�g���l$9$5�Z9��^�D��'��A=(-���p-y��2�u�AEՒ{?�i�C�zs������Xk��P� � ���*h�t.]�$�^��ή<�e+1�f�x_�D���}�{o	���z���������է�����Ι�yO��X<��o����h���_<�0�$(�r�/.ꔨ"�<s���z8AZ���ݚ���ēuzU9�]-L��; Bgd�.��@��hY���(jAf���`-Z}��x���t2Ҍu,����~�3�y���h�#\JG�pkcM�/�A}3;"�(Xy���Ӱs/m��y��$UdhJ֧CA� T>G��f�ϳ�a��1��#آ�~�<�WN�������~zO�u.̹p~�V�5�]�{��쨠��K�BNl��߳�6��,�9�V!π�B�sd��\����=�\�EK��Κ6��Д-Zk��T~�թq���@Q��]Y	8�~�|q�=�X�0��gQ�A){�!C*T�N@ 3t������!��sŽ�a���������F'��ȃ�����a�������9OG��'�x�m�}{�q�) ��z���}����i���E9� ��+����0�r�,뮴-�灃rxx^�a@(�����B��ةX�fl�K�����)��z���AX��&�_��,+ ����b�P[��A�_����h����[@�3�4���0�Zi缢��g��(�L����Z�1��_'�g����6�mt�3#<�����ahD�'��(묞)�]o��	
�)
x�`N��9�]SfiJ���&�U��֒�_���5�o�d���hB���Ï�f�_�fh>|���P�����\��{@�޲
˙�@s3�ҟ%��~�����P�Y���7ok�Q����j<�����DDضĸ/��Jj�p�;%�&�q���Y��:0�9�$g&TB�C&�{T��-�,!eC�=3�ZcW����iٱ�@t��r`0�H4�F��_�*s&�eu�^����&*uT�>l15v�=_�|ea��|`"��cH�kG�is��&�֨|��~�hoj�YB�b<����9z-�׮_��!'�Z�E��t��x�E)@1����S�6��G�e�o~ܒ
�����o���_z���E�7�V�G6��BMS�034���ɱ�$�X��XAX��G�K��c��~�3"$JO�p�Ihj�}�$K]���yJ!_�G'��[�9��h=���]0�$���$\=<��`ݎ
bXi�G)-�N�żAe���qe�Z�r(���S�;m���VK��eѰЄD+�9Z��1y[���P_$E���Ck>�"��f/�{�MD���;g�R1��#��6�;^�!/_����Iφ��-^���UϬ�d�x4������ubS�����|3'������'@��N>��bgoW�-B���a��@y���̧``/�㪬�)˅c���恞��<�I��V�����v��Q䍘��|��J^]�A"U��fq��{���ꇏ<xo�_�׃�����3����lx��o}�[)r@4$�����/��#���~���;��;������-8nI��ē_��'�|i��͟ZYnN'�#t�������-�L��/��*
��;ׄ���ŷ���XPX�v&��u'G�e���VWa:-�7n�Ҩ�^��֪�ѼK ��郈uwU�^3nS�6ƃB��K�QCnz��Io�#t�{�	%��M�R����s��-�zU�����<�(���ê6�b�jPX�?3gABW4����RB���5�G	>���c���օ�A�ԙ���ٲd��)�*u*b��g)�Oa�+<$&����@d�� `<�D�!��ʌaZ�T8�cU.�&�A�ʥW텽�7��ueR�l��F�����G,{�V��e��<�\��c��T��9��"$��<C</�F#�Kr9�>aU�0�g�����W�j�E�+)p&8��=��AEsż�@V�C ��R	�(�A8�a�T��4��H	�C�\(Ճ���y'�����~Q�?�������ʆ����3ѻk����xJ�aW��V w  �	IDAT'l�^ox����{���k�����G?��?�w����o�x&n��qA���h�ٵp**�˯]�FC5\����?g��k�f�C�),���Oƀ���ʉ�Z
�,�-�2E��d*T�2�Y��bd����iy_b�Ae(����3�Цpf�ڊ�E#���Oצp�1�BMB��y�G��f�����΀uRd�E���ٳKh��y����;y��3����h�fF�l]%����0&���9�.�gR�b��UϡIހ��{�\T�a�*�F%D���tN*(QX��Fpއ9���7G��ܮO HJ�׹}���X���h�_�W�k�Yܣ�>��m �Y�s}���nR�rʝY��s5E� .@ѿ,%Tdy;�.yo(��{��W����\��|�և"k`T�̖P��WFT�k0{E�<��^����H�jhf\�]w_k��i�1�����b>���w�;�3��o�vx啗�<��A�kA��*���c����<��O�3���->�e����������;�}4.�6�R�Ұ��7�$G��x2]:�8HW�\��-\Z�j5��N���&*��XN�R�`�1O�A���T��(�f6S�K�[hO"�Hj���5+�����r�1��n�)RM�v�)z��08����m���#�`̠�CYa@c>�VCw��k=D#���M�&`���-�h1pYj�0Zך�@/�ԕ)��zh;�;
<Z�A/!� |��Ԛ�#�I�3��C�/�

P��b�%�6}�z�|����}e|�$�*���W��;�}1��zX8�6�B����S�^a�j��)�D��P!Ä�ò&T�F CN[���!�W��4�;:���m�����e���|��!�c�^���>���3ʼNUq]H�O�sH�C�r�D�ጩ���o��zl�`�@sm��B����c��Dɵލm]��Y,�
��!z-��ҹ�/�0��=��#a75H�^Ir��7�7��o0���i�Yy�m�/?��O�n�qK+������_��W���|tcu�����AGQoH�AH ���@l6�D>a�4-dEA��
���5�u��Q(�a�7�r�󒂲��F*�k�%���yꄪ�B�L�����U`�=�S-GH�-Tȴ�j�v�x�������<m����)���v�W�*��"{T��&.�v�0�����x�C$��uoD������$z`��0iM���)��M-�<��N�{�#�/d���-F��(G(B�n=���T��g97��(@���1�����(;z^�N���Rl�L�ù���\�QY�5l=MSPv=������ϝOvjP|:�����x[��1�>�Q�,��rn���v#��GG�awO�-��Ϋ�x�` Ll@�0C�{;�B�jŭܓ��YFÕn��bXfNiCn^�p �~I�s�R�ua 
E����4��*��3(�,��)�c��8CO���sωR�\A�#�2 �~T���E?_4�v�}�x�˟��'nY��V@�����/��җ����hAm��������a	��[ Xj�#a!x���{��a<�~�Nj���4��k JF�R�-�pk����B��f�u:�%�O�夡0�ۥ�H�B�!�J�t/��Vki�Z���*b��q��'��,K�|lD��Z7{0a�!	�xʨ��c� Nmn�⚎GB��bBPuP����c�5,�v��UB�Bj�2"����p?�aO��@m�� @��*��	Q�����On��{2$F�ܷ�f��e���WIQ��`�DxQ �'�9SXG�6��}��Mi~H�W�ͪ�����jG�����)���U	�*� �I^?E`�� �k�@`�
�͵;�@�mon�^�?<Ly
J(z�x*(����B�S���OG"0;��|��i�����vndJ��� Ƴ��
����<�!��Į�E��͍�ua�&
��J}Z�އ>7��aj�=�|��L� �ځ)�(�|T���,a�����ko�T�v.F,�d�E&��v�N�0*��.�(x@!�=A!b*<?/�t��C����rʩ�FTe�G�ֱϰ'�}�YQ���c=��ٳ���k�J��f�I���8{_�ԧ~��O#���W@��/���������x�?��u3;��U�\��\��:`�[�ŚJh��m�-�L8��Z�P���
�\唰-E!�vٕ>�����un��EB7eʏ�B9l��c��2ѵ�us�,�v!X �4��Bg�*���
h����@s.�����)�{� %�E���I�)\�-2
�i|dL��N�7]H�y�B>�x(W����Bk��IX�.����N}mNNT/��$���{1��E�wp��d� bѩ�f3����B	Z���6P�a�X��<zQ>'Ƅ8���sW�1C��'���}y6�����W>?�e����IA�um/ � ��h��^��ء|��)t���H�7���x�������i��,��suP ��9�L��N]��{��I`��(���<�@t���aTYP��f�fUYθ�*eh)KF@itW�
�ϲ�uG��zѠb�=R�p�G��n�79ߎG�2g�-�s|<���������O����-��0~�ǯ�����?ͦ�G�bn��.������G�0�AΠ�,�W^}I6����S���H�6�5B�M�Je�յM�$$Mꏓ���)t5�#6�n5�4��x�8�xTe!1'���l��$	 ���ʌׅǅ�/ĚXM�ToB&ftt�U�김1A��rV���jg�`J�<��^�4	&{5�r��/:�ȻQ�J8�мg_8H��CU�	Yfs���BǠr�)T6�L� ,�'="���8Y;��<l�kQ��BV�غF��%�l
^B�.D*�fQ'�2LT�S�0C��b����5U�/-��6����{�i������(9	O�irҝJ6��f*�Mo�-�ޗ�Q�`D'�9G��>�"<��jDQ��kjQ1��Σ�+����|	 �[�`"�Ta�r�*{�<���	s�,�Z��8=�r�t���l�4@�m#�W�C��L�"�<N��A_#0���|}��ҹs���#�\���-�SO=�����旞��ӏE�pqQ�.&�]Z􄑆u&�i�i%p)�xkS{� ��(5,�ALq�����H��w���u)t��=��D�4l3�B�kֻ/���T��M�^d_�`KPہ��qC��qQ���?d����Z������ң�Jz�{]u(:�ʌDԐ	H���\"l�y�̍��^F���D�9+:	1�\7�Yo7�?76������%c��Okפ���G�qͼw�!�VTI����9f�$�#�c�C���1a��rN8Qq`0�2lc���
�4��s?�zZ�TҰ�i�`o1�rx��C0�S��f*~��(�����J����SD�	g��Q���z�o1���J��Cy�ht� #�z�s����ϵ�Ư�%���rKy� ���0��A�/�Y��,G�Th�Q��#"�0*J̏�w�ǺAѸd�,2`���\�s��������Z�sr�
���w_����?�r�����ߚ���Z,�@�5�!wv��ju#mfӰsGb�;�D���V���� ��Z�)�M�2��fR$[muBr
��ѹ#����*����ˮr�*�\�w�b.y%A#T��� rS'�$w��J��FkHd�Y2v(d�KLd.����h$�S������\)�$�1����ף0�g����H>���&:o�B{!ϭ��@�Z� ���>��憢+�%q��V�Vau�BxÄu;��j� �ԕU�	:t��r �5_���NAGe$�h���G�y�º|�GO&����R3����*yT�NǊ,�Cm�"�bC����FVe]F����TH�G���z|~�3jQ���gh�,e�S�g!Fx
I͑Ң�w�/�!TLミ'�6z=h��y��ʽ�P�
g]C�_xJK���ߊ"S�Da3�bD4�t�d��r
���b��'�~B��5�zp_c`4:�N?��{�i�E2b�
��YOH�J6�{\�㵵�����x�������mЃ~r�����<{���/�m}�d<���6l0����U#	�^N2���
 ��@���,s��m�	I�w���ʄ(x|��9������������i�{X2��l;��mT<���
�:��b}v�6`MѦs�)o�����x��*���M �ކ�Rb�����}Q�܈x7�̨M/F�F�[`�!\��K>��*�HWG���@`��qN.�53\C�'!���+��ܺ2.��)�6&z�+�>�5#T��	Ǚ�Ѓ�2!h���qz0�F��R*�9?��-ާ$�sQkoh���,ʢbΡG��"����t?�|���g��d�|�L�c��y� ����A�MƋڣ�C�����O��y����\�>�
�]�Q�"h��B`�ٰ�9BS�.���,�z�EZkii��c,Ǡ1�s�Q�|���T�����r-��˿���_��_<�ɸm���ڵk���K/�򾪪O�5��֜@hNǲI���p3������`/����J?��>7z��ź�|E��UB�S)���u*��z!n ���V
�0�f,�aY�	�E�3(�B,[��*e��&$�oRV)הu|���J�M��c�����c#7��A������,g덓�M0H�'�]����-VM�]>{��%�����q�5F>
�չ���BG�As��)�09�7��^�\j���,��(p�y�����5�_��嘻�q�tiu	2M4�3��V9���4&�\�J���7�9cA%�-�}\�`���t4��I/�#�o	��R�M`��+�{Y!�����k�0����]g���w�b&���R�8�CV�a�z-
Q/d}�KzN5�(���4d���W������H�&9���3��V�/�t�9J�g|g��;����eѓ�$C�a���8�	/����=�O��w4��?1�RY�"N��!��Ѧ���DR����k-_��am �N�2%P��ψ���'4�U�F��(����'��eY�l�V
�'�����ዯ�r�qa�s<����wpЊ�7B�Ƶ��=l"J��O�n�)��,"����R�Si%��B�ER@TH��nz��ҙ\��Gx���3�z�em�	���[�R[���tH���kҼ���;�XvѦ����1x�L��3�xo�
�z(�*�9�/����fX>���>�|2�ĺ*����c��s�wx ���)�iUbP�����L8�N_y`�x[o�^I��=&Z�T�^��#��b��"����!!ڬg� y�x���A*��`ǽ�-��p^�\���l��{+�ވaC�G��%tZ��0������<|6>�hUzb�{�~��Z{�ׅ�E�%�ݗ���sR�{O�w�m�����*D�bT��&��y�����^zP9���H�F���53v`�0�|�sc��]�x��߽��������gΜ����G�}��g�6�����_������W�����V��E��f��@pB�a�: w�ѵ}M����,+T��!j���K����V�GZ_�Z?#�,�t�N��Jh��ȕ����k2�������}|.\�&��	�.�mW�ĕ9��#9�A߀�K!ExuRN�~=�0C�k+�D����0-�s�p�lƐP�����	�����ZH����F�N�#��M
����Gv �w�����]�G��m!��#P�Q1R�KȦ�]њ"��y������Qm��� �@GQ �4B�*�0ѐa�P-l)�}_p�&���=E2���=��_\0<z݁2��]�u�#��E����!&*O
b��ne���/��̈́:πp�W����q
tx��_�G������m��<#Z|7¹�88j�P��@#��[�ׇ�[��7�4w�\�Z��ϙϠsR�'���p��z�b�YH2D 6��/H�,�g�
U�{EFX�^Ӱ=�4bI�
�D�{k	y���^ö���Q���������V��m��⤷��p���^��������`��`�\3<�֚�5� �^��ƪaZ��*#en�IsY��愥��ls��z���x��	�@k�¿(2����t#ro�\@�6&Z5�57o��ϯ�@Z�g��-�[���� 04%2D{�a�ߦ&��r�F
)>�Y~�
-��������/z>\*��x��X|A&�פeK���LAM�����o
Q�,$ܻX$!�+����� ye�:!�(t��B����ϫ�Pυ-4.\�C�^�9���5|�����4e�,Hj�)�GV���D[<=5�*iH�lO��;J��J�e�2�� ]��P �J.����<x<Ӽ�G��9`(�0��Q΀h�z�ـռP���\(��xþ����\���Ϝ'�5�C����B!������>���q���K�����k�6����ԧ~e��~����O�o�U�|\�s�(q�� ��3�6�n��Y������N��,�!h�r���ún�2)�`f���Z[@��ْ��6ߠ(;�[э�\����^��h��R<x)��z�Օ0�lA2�BPU*�_�^�������Yq�T�DuOC(�"����+(7K�B�y�J�O�HK�a;�b������(p0��S�B��
��<��,W0F+H;X���8�E��ŝ4��XIÂ�*yv���cl�0 |R{� ��)A�Y�
���a�|n
y�7�6�~8ʡ7���c`�^�tQ>c��PЂ��Bׂ�i��F��t��^�(z�q~���b��}c�l+���*��>A � OG�P�֞��@aUt�жo�Y��m,̆gBϔ�bc3<�Q����2iQ�r��>���%d�����puG
J[�g)�Hk�o=C�	�Q�l)jTί��G{x?�끞��W&�ܖA+Bˋ��Rz=zW�t�'��ը@�[F����&	/�������R+nC^�uV����=};��-ƃ>x���������n���GC9���>XY��I���B���ђ�^qq�:�q=������a9������z4���ϩR�w4.�M�c�T�T%k�W��B Y4��tS����#i��O�����G�)y���`G�{�vR��&��C���T��u��yBQz����x�P�^!{ʇ�0<��VϠ��P^�q}M���{xbO�z���ä��(ރ4A���N
B��q��E$�_�zG���u��Ӌ_�5Y!���1��\�3��k˜��/�[$\�SZ���D������#��@ϒ�u�-����A�2���Z?ʞ���մ�uܫbX��yM�����Ò|V�ֆ��B�W�X�S�S�Xz_Utҵ���3��|��r0��<�Y 3z�������1��~�����8�g�����tܶ
���������~�K��;;U�^���.,����xx�i�Sasidw��N�8u�*�;RX�)Q"p����M�:��G�u���d���)��(��@�Z��.
��E}3G*I�l!ú�"�!՚��p�i�L�t\���*�.�s&(��S���&�!Yk���U���6���g�^���Z
�\��*-b�kWPi��>	��-HZ�/y����S��E��pᶢLVcNWI P){���h<�Cl�vh�ҩ���%���wx⥴�O���q>06��ě�`���>���C�+Z4�sa��{g����~\�rPysP�D�q?�>/3rR	gs�A EYBAQJ^+*G2ͣ@@*#�u�֓������z0���g�O��b *�bkl���`��ʭ�����.��cɔ�
8E(��<������pj��L~������N�9�v� �4/"9�G��<"^��+�=��?��SO=5	��mƥK���u����s?|8.����h^6&�(,H,$O� �����=ؗ�9Xe=�0I�x�S!d���ŝT@�x��P���FQBu
7��bi�2V]9o��YU��ӷkKe�x���'��H�a�p17���"V^�y�¬cI�co��v�Q�T�2���������xV��ߕN�K�9�K�@4�/�rn)C����|��m"�3�N����� ���!(f�u�k�=��{`+�I�_z��P����~���D�\?�S����H؏-ʛ�/<��!#Q�2�Є�,�BP���^�B�g)9���[�t4Mk�{��3��?[�#�QBѹ�f���lT@��.�cx>%\� ;e�iz�ד��7˱�<��kg{楗^J�-�3x>��k1�D�q���܈��_?��_�{�F���m����_|����h��kW��7�Z<(�� �H��ʄ�>@��@j��\�}�Z[�Xx=�7X>B�ð�m.ЭV�����b�G�l%z!�$2��;p�C/'����Q���W�������g�q��҉V\�k�w#U'=�z�Z�ȢR%g�v�n�vij�*�����YfUa�'���@.;�I��Iz<��p�e���9�K���gD�� \�lYf�!5PV�$V�)L~&Û,Lźfn1]gz�#���Cc���BY���y��;�c��*>�,��;��qA�<[R9�<wz�Ya�pk�[��s9��Q�`�m�6E������r���`�CR�4�&"��C��T�4dCnB	���{j�v�� !jG�@
��¸��62B�[7v�rޑ�%��U���0�x�����(�ߋ��1ǰ���U6����y�ڸ��wx= �����r��2��{.��?��?���?�c��ḭ���v~��>�_~�GϜ;w���Ν����XZ�:uF������A�J;���k���ڦ�`�K���G�Lࣃ�	+��Lrٚ��~�� �܊�;��=s�3�gQw��N-�2h��:�ש�����Qst4��]��aA"/�s���Ē�򵡑���X��lU���	�/�D(�G+K�5�u/U�&̎��;B�xV�~H" x��$_i0�Do�3\IB��|�̨�8�,���3���!6$%P��0^��T�"h�z��b.�A��z�$׏�� I�[��mzV3˿2��mx�W����|Ǉ�(�=#�o$������� 	'�}�?�m\wh|��0�0���'�N�k�g�uOX/D�g��,�_c���d�;�t�i0`�r�e�J�j����B"|}Y�|@Z\��;P,��0\[�g�
�&y�Q������6,�).��ul�}�O�U٤��xwe&7�����稵ZM��^.���%��C��Q������w�v�{�����Ї���/�������y n�Ͷ�Õ�GW�3����0>�H�F���W����W�:�O�I�(#�2��o��V�-�VZK�X���԰@����u��ڣ�XP	M�j[�ʐ$�=���D�C%=�V>B��Vׄ9���P\k�5�4�R?"$�(�C#Z��b��
��A�t/����� ���2'}�pu%l����@�9�xt��(��9.��� ����P@��b��8'�,�G u*ݎ(�i������ X�0��$l��'�5$A�p�=#(�;�6%�1k��<��<<�(8��c8V*�K�,l�s�F�}C@�=Tn���7�JO�>�W*Q-��њ�+«���M�52�~ �0/N��+]��v��گFzWY��$�3�T����R�,m��_���o*C���p����@�����\������
�<��8�h@�@/���癀�Q��+bn���<��g�`��W	5���W�aE��NOQ~��F��hb:�U��(��=�����u^_�\lW�G!<Z_��5�}Xh~����U�TI݈�l���U7�0�ڣ��^�� ��}{{KZp�}�;(��w���9�_�q��Wy�?��_��+���n��P@���������o��gm;�;���Q������j���W�� m�Qet�C8<K�,��M�ND9��g�G��s�5)������n7]mb�mw��(��ģ�4L�V������2;�S�,S;��c���gDIZm�\FA��%��ka�2T�!�|.�4X_�C_�H �Ջ�B�3��$4Cf����I)r��CQ�B(C�ϥ"�D�M:�����D��|�g"�k�1�C����oU��d8�W�p�����+�H�ܙ��J����7��8�'�@�z�YS�{��Z�Gft?��R}I�-�=��*!��ĸ?Y&��R��--L6���vh� 3�.���x^��A��z٣���d!�=Qu�5P
�p�d{�@!��4'e
A$��E����y&�,at���s���=¸�� ��#&F�teu���:��5�ߩ:AKs=>����ʭ��u\����o)��n�+0����iPVb�mn���{��!�5?��[�0~���w��G�?��˅�ￍ�;Ba|򓟹������?��Oo��[�N���泥[{>
l��5��Ͳ��	�!˅uB�wyr��'2����[�<$�o
Xh�?�E��&����'����Э,+X�U����}.���4'��*�m�@����x��� ��E�r������9:�|&�M&�QGQY�G��BL*�-��j6�o%Z�ړF�y�-~�T]c.Ta G"D�X������,��BzL��(�e�&��9�� w�v�#�1�p��u��4g t:�ۅη�{z����1��Ut���j�,�(�>7����!֮�Z��\Nb���x;�* QJMf-���%T��a�pC�Rl;ˌ��yDx�&s�p�*P�hT�Ei9�F *S)ҍ^��@��W^�j9�Q��H3�6S�07�L�M���%�\X^1��|��}k��'ܑ�+�O�?٘�z�sH�#�3�ou]nU׆�y���#K��ׯ�����0	&A�+Qo�7<$��R���h ���{웿�+���!���0~��?����������{g��z�@�8Ԉ]c3��pA�62P<�yw��@"H_~��@#�s������|��P�^�rS���nފ�5H0c��Ԏ���������=b���Ent'qx����vo������o>?�x:�"� W���dX�A�E%���,�}Tx3���r'*42��_���h�
1.Ei���j8�g!9��6����΍ظ6|v���B� z�L�#�m�:�����*Y��<�7zl�1"`H�j�"+Y�ZZ��2q��l��^ &f���4��m�����E޳aY���ZP@�,cXG����K��"9�to"�*��F�I	ug.P��C�M������ BR��e�z�{x�G���H�Q��k��Ik7��y��ׂ�s����4���u�\P�@�]��Z�(F��k�q��+W^�y�҂�������p���|��ۦ�����R@��������3��O��;,z��$.~A��7o�������)=䏏G��um3)S�����X����~�|B؎c��~�3G�p�Rb�k�"����B2.<���*ta���IBS��X��lk������jr��heQ����c���_$Je<SR��/r���V!ZEdP�I+'�&�6���A_5rO�e���cm���0�H�De�S��t����4?�Ҿ$��d�r�~�=W�����w�Y
�z^��%�����8y�PԍQ�PQc��JyvP0���_1x�(��8�N@�9���0��}J��$4���������!�`mR�(�2X���0E�	�F��Q� ���h� 5)m����1���	��|��:� D� ��B���i�@V`��������\ìE�Z������z���Oax���*�"'*���c_ͨ�NOX��KŅ�Kaj��}䬹�̱D)
�z��Lm�e�s�={:�}�����@�x���i�76���J����� d��R@���'��������7��'n������BIA��@ gЇ���pՂ:y�h��!�EaeC8h�P,�7r���3U l�@+�r.���!����p��I�f�|�&�UX�kTh�R�G��*��.�J��a
� �Į��1�8���r��Iz�Q3o��0	��A�h���l�,��T���l!����H%@|�-�9�a.U$�e�tQ&ŇgX_[K�b,l���Ɵ��(���q�Xc$���^O�j��˅��ҳ�۴�z�>O"��@1�Z������$Xk( xz�dm
�[T��3���[E8	��-��75�'( \gogW�sj|N�_"I�?ڭ�g�Y�1��i����;�B��K��\Μ9%
��ũ��*O�mV��?�%�O���ZdeN�����"�\��yC���װ�){��u�G���G/��?�'�͗>�O���S@��G/�����^�'.�Z\��H�c`���gOkW��x�6%hE�]�@��B��BTR��u`� Ȃ�[U*ZA����%ֺ~"-�B�=�Q��#%.-_��D�SG�$��C�y��P�61�AY���� ��k7M�C	�C[�)g���$�-l��K�2ѳ@һc�;Y ZxH[i�Q�p��ޚ	t�fenH���^"�`ɖ����8A)[r+-2�h�֪DK	�N�\nDB�����fQv]��jvS�Z�T�,�jll� ��MhB��8q$d�$tq�K2� ㌑�<��xx��9��s�H'
8@`�c�iDlcL,����TU�nW�~����~s͵�DB�`[{zl���k�vο���s��O����y T�Bɫ��S5JN�^l�Os�[���#�pQd�	���z�.��g�9S$2�C�a��.�y�,	#����ZJjK��\g�_�a���ii�u9���
x�������	������QC�=� ������DNۊ��ή�*~��@<[S&
4QcLzL�{B%=r.B�0��3����61�@RA�*�������6
�3���Pk�w���� 3�)jӽ�0  $<uI�
���y�HAM>���r&����W}��o��;���6^�
n�ѣG��^��q�`���֢�<I�1W�ظzuQ�[�F� D������e��߿�şe;��,W�Y�W��!���0AK
���7�uF���/2�cX�P�&�X��>�Y��H���{�ڽ�(�؅ߐ\Ǡ��kT>/Wr�2KShP�ʾ��g��l��PD�ن{D0 Vp��0�����1u+54'�k(����-T"���#!(�G��~��6��o�{�_��'y���ưֆ�C�
���>$a���Cf�"�^�ܛB��^���N��Q���۶�����I-�|�7�
Y�Ǥ���ųn�g�XO�C�H�A/gȜ��)�Q��r��X�#s6��z�%Q,�ű����TJ�5cA�Р����=K]ʼ�J����-Z�9#Կ�d2 �����(j�(����:�B�K��ק����w�w�z�6��x�$�<P?r�?���}�3c��3�v�#�˘2��+���biӅ=P�g�	{��E��@qX�d�%+U����;��0�h7�Z���R�G�PQ�9A�����n�����>h�g��ִ��J��׷������H�I���x�9fM�P��Ү�橄�M��7,ڧ"�Y"L 6P��*
"�vԊS�J/�1}*,�&&���6�ſ�@ٯ���t��ܖ�Ŗ*�4�:��m?�BVQ�b�X��e�9�$u�BCy�,�!?DH�je*V)��Q�1�^X�	:�g�}�}\�v�,�'��S���U�g�HF��
�j)�������r���_�h���s�h��cȔ�*�)�ƚ'��߯����6��!-�|���~�?(r0�M8�A*cv��s2w�|M�D�ǂ�$A�
�Ԇ�-Y� eF�.

uz�6�k�jϞl�����%6��=��wJ-v��`"�X#���ڊT��u��&b$H]6�]SA�����ں�/%RM�敛n�I���+��s�m��K�B���SF�|�����Ơn/��U@��{�������S���5�3� +�/_����$XY]s��hh%�hf�bB�;wN&�B���h�i	r�B�+b	�~���Ru��@�MC	�d^�	��P|��Ta>��$�R*��K9��,�E�8�)E�F ֍��d =%Z�r� K�cP����sJǷ"��!
O~��� �Z�c��N���d�Iz z��e�@#��#� 
 l82���'%Tg?�w��hY�}�	_拨�0�ܙ�ΐ[�Sa�ug����RXʨq��K7��1�O�)Ǳ����!"Q��@2�N�vz���OMC�A��.�<�M�T2~6�5�g�n|�v(7U<k�|��ϔ�X?�P��@}�APdJ��� ��cM<w(v&E���H�n�gx�` �@k�l�{�`�왳
�c�L���w	͠/--�T�Ԙר-$?���v0�ۮ��<�_�xBs/��g^����|�»����:^�
㝿���������;W�Wj��;E�+�@{��w���[Lr^�pI:Q��Sz���^��؅����5�
aZ|� %�&�5��� 9"���zYT�ql�'C�lW�5p�X��~%����]M��kڐf)q���'M�rP���Sz�3d��DP����N0V*l���b��8�|��.6y�\�]���4)=Z�z拺�C�~,j�+H���ײ-����H<#\��`7��ǿ����<�`�P8%���X�d�*ǌ��!�8HE! ��x�%��0�)fɫ����a@Y���&�{�������"�;Y��0(�����q$wh��n���P�I�����uO��0�B�A��iF�)�Gj���p2di�A����[P{Y�t�,�Y����y�yJ����_t�
1)YL�8ԮOܜ���@!�ȶQ���9�X�I��mqi%�$�Ms�Cy	����Qi��s��.̺��ь�9ڱ�����;��R�q��о׾���#G�������n���x�fNt;� 6����F!��0辆p�J�	t
��ZM�$ik�#��*�S�C�	���#W�1k���QH��w�q\��e�$=/`A� Ѿ5Z���!?$.|�ŧ ��&�U��[o�%A#{����ׂ��Y��F#)'C(�m֞�e�Z�RԺ�������"�J<>=�w�AX�E�(:+6�
p`��)��ĵ�%(  +l�bc5>�*
R�;�@�Jf�K�[�yT���r�ږ 8���|ZdϏ^`	��Rv^��:�ON9�#��t�����.&����\�7߫�����j_��s�gOǇ�Q��Uw�J��ٳ9M*$zQ<�+ъ���~蔍�bzb����0w��)J�l��Qf ц���$��cת5w\>3�Ն���#���R��#�� J!jߘŜ=p���߄�t��xIl�n��K�7�o߾㓯|�+O��L�/y��ˇ/������j���$�1���z}�:a�	�z��(q|�ТXl�Q�� 
��.X �D�S��FeZ����~��F��
(pJȇ�bP�p�CH9F�s�o��_X�?-����`Y��X��xF��E�C=���aݎ�B�B�W�Kб���:�}��ޤ�r��)��$�@I5��#&u}����B�pҀ���z��	a�8r!I��Ԫ�\���&F��%�(�_7h�����܋>�	��U��rD�쪺\������q��@���������ds�5s_���fѱ"���@42�"�Sl��9���R1�Ꭵ1"20(̽8��0�y��u��Bעβ�I�4b h�����3xE�;�I�K�uQ��܅�j����-��ܛ�^��x@ݞ=^ʈ�0���ø����'�3�HE��<Z{0����,uf����B�ݕ�[�$z O��v+�Y
����,���K�+�~�������}{��7�����������x�ޟ)�{�yI�|�q]( ��>x���o��s'N��gfиy��0yĪMꮳ%��ϟH������k!;E�ud����u�hb=���hy؂ï� �0��`�V8��Jm��A,C	_$ٹ�5D�K�'6�λ����N��D�>u�\Q�pjղ�g�	��HP�9�Q�᚞O�� ��p.����{��aj�D/�y��28|l��h:�'� wO�*��U������,p;V�ӊ�+�Y�#���>�g�����m-y�y"	�~�\g<W�с%�����JE��F�y�K��7����wzd>E��0�ό�ͦk��$���܀s>h��,��s��<Ȧ�v7�zR t@���y�~HP�6\X�d(���a-� �C�\pe����&H�����g���Ȕx�������^������I/h����<YX���a�]�|7k���7���/=hdUp���Fa��[�rq����#�+��̺���n. �0񐟀�|ٸ�ra�$D�@�a�@Y)�X�I�I��]ۘ;U��Zk�C�)	����Y�h��L���6<łRW\6�����J�z��;�~>�+��娬|a6��z��QV�X|	�Z�#F��I%!�^b�G)���jZ�J��^��B�RLz|e��3X��,ߕ�U�-,5P`�(~m�:�aP��:
R����K���i[�R��/���&v��~	�-�N�[̼��c���~F�`�s��(kh'ޓ,��0$X����<Ĝ���t�H)6��$�J���
��E�q�h7Ђ ��a�`���m��іa}�)�z൪¶m�5-�sR��w�� jp�dD�0J��S�Hd����o�7NOL�S�F�k��W�����
���,}��*�2���Z6��G>ߍ^d݆�cb���^�WV�}C�<���l��ݷ/3o�ϝY��5a��a�ٽ{�~�~�-����˸�X��;v���#�k��;���WFFfXw�h����rAr���s.wQ�-�/_���^8�ƃP#;.ڷpQ4Q��JS*Zp�,_�͉]�Q�g&��iN}�c�5,��u7��^�	�R�n[ w!���$[KI��!BkQv���u��$I؈.q�:�;�)�4�yr`[���m+C1�Q�އ:@��?�� ��w�S���/\m��b�x�8�ꤥ�� <pU4ȳ��0Rۅ+���X�(��e9�U��<>(T�v
 ��m�N�Ӗ�!ɣYT�	� _1�E�ٯU�~R^�J��VR$��<K����,��}x�@hb.!4�S���Fp(Z�s�A���������u��"��ж�{�W�\����ֈd�\~E���2�{�l�n�Zz�|�|'`�J0�eR���6v�G���J�!^2B�%]#e���[Z	�T*�[�E%���4(�Gʄr����ҥ+�^Kc6����Դ\# M
:8��l;g�?b������-� ���h\W
���[衇�K_�;��o�t�w���+��}^�m��$6�m�V�i�tEx�"ce-Ⱦ��Q�k���RT�0�db$�?��iJ�_;�VD��N�a�����,}UFp��S��U��lZ�gjh���qq!�"Cf����!���n�̊Q��Jw3�Ff*��E�j�S@.	y'8i|�����c�L�wh���lA�m��c���[Rk�+�F�L�`vc	KE���B�t;Ay�,��J���"τ>k�ubB���٩T��Dr�~|<�@�c��Ґ�����Ё�$P�k��7ײ�WyD��@ �T26��|�d=���\s
=tZm>���]'bN��a륄��?����#���JM[%�HR�Z���ꎌ��<�Q�k���%�ꧮ�_�枤ht�L��Z�xF���G�'I�KG�bL ��B�q%����u��K B��pŘ�����v|�$!���4��ym}-غeZ�h#�^�̊ ��.��J]�{W��0����c�����ʖ�tQ���W$���K-j���~A����g��	�MXq��(�Nc���m����o|�SozӛV��l\w
�mo{��_��_?��c�Z�ޤ�r/_]]�*sqW�� ,�'��i�Y`�K�JY녚F�Ï߈�E���jpZ�xOA%byi�K�F>K!ϰ���x���b��آ��Qڻ�$�:g.�J��<�#e���m�X<��O,�Aٞ��w�����pZ�������m�j]iG�,]f�]k)j�Ըl�!,rM�~��j��Z��zꍺ<��I��yLMM�n���JO��w
�=7���=ך(��4K[�N�y�ˢ������M6��
�>�uX�����K�xQꎃm�[�o@Y
�@���lN���k|tJ-�lS(�J��K�'�6xe�w}�5��[o�\ȭ���H�vD��U�1h�B��Ey�c�y�]_�����2%_Ƕ��6d��cE�YxUљ�l�l�0��-��(i�8pP��3g\��z����Rj����_�&�m��1��T>h�"��,]]v�+���|2�r ��R��[�k�@yj|t�����|��߽\��T@�|�;/��_��g����4M���Wo2-B�H!�e��� !&K�@��n�'�.�bQ��&$��\�"��|�b���ڽO�L	�ʅ��d1�Q�N�<h�+Q���w2DO��ғG@D8�y09�\��B�^F�n�%Ud��V�GqŅ�$�aB![��:11f��zbj�l`IJm�a$E�:
F�xy��%t�� ���Q�s��A[uX��eA�ި�%����{n��c�q�#$Di�j6�0]���Ep�CPD]+��@�	�� �����}a[m	�5X^Yt���0��!��^�`��b.%�F,,����)��w�C�aO���K�2WT+Ƌ	�k)9�g�u���q����&�׋�2O�6�)�Uq~3L鳆H�X�&}�z(����<���t��,�x�$M����	g4�5x�VX��J�yS=N��f�M�*P(8 f���%�{<�}����Pk�P ;���R�l�s��H��׿�g��O����u��0��h&�Ǟ�������I2���&0�3���$a ;��J�������Ӑ��X�]�y�M34�?����Di�;.���f)^s-8�a=Z�l,�9
zH�kk�^���wk�>+�ŚX���zs��Qމz=<B$(���H�j�[��A��뢈&b� �> ��Q_��@�����(��D��c��I�6�+����fR��盅ಞ0|��Lj����Jw*(��~3��l-�<�t|�98�v�]Ki�B{�]^C��5��)+|��h��g����R2�:7c��P�:�;���|�\X����ݦ�[�h(^-=P��)�s�G}振P�d���F����K�{��2{��P�J�ޱ!�\�0O�JT[1��+%���=��w�l�C���d�n8�g�}V�n�c�u���g��ȝw������/}���q]+���ر��.=4X�Mi������lx8n�gvJx��:����B�P=p��&؍�A?(���U3yW�B��@�B����I�>����>����������)0�D� Y���gE#�e@i���wdփfu!P@�+�j:τ�&�B,�^�4���R�i��=�V���������0Rv��F�/@	���V7�fu?���=�?e��"g��mk?g�WXˢ��D,b7����͠c�ja+��
f�nqD�[ :���=f��(6kY@�!�ͭuWZ�5&����`(Z�P�����WV�J�r]K�䷝�S*�-���G�)0q������͹��k�.8o�/U�f
��
�m63:�y����)6�sH�4��f:p�+�׶�oF\[s�јsx��+��Gc
H�ä��^?3��[��<?�0�(�r����@I�9s*����y�Q#����+ O|����Y�]�����J�r�&��0?�n?z�=�̆/q��k\�
��/|��~�K_
N�;=j&�Ϛ�4�	�� L>X��b1�����m�A��|�����B2�ĒUu��E9��Z�9�Z��=O
Z����\�daάN����AV�b�W�+ �S�������>�2���mk���C�J3��K��BxeEQk"��qp�d�f�!K���z(����\���[�Y�2S��9}����}�O�
�����{KA��}ޑ�˸{�j�-O��sD���>��3��v�Q�Py)�M���^Fg�7B�U�vr,~b-��8��Z]�:m������ID�ѓa������s��Vir��܇��ʊ�q�E|%���A�w��J��W�j�\Ysw��!�טu������d��?{��0�u)���5rw8O!^%�k枧�</��ݷo�'����;��t��|\�
�O�ӏ7���}u�긱X��Y0�|�D��1 ������c�XP4l�lzz�ĝ�|�		* y��M�����.|iO��^B+����sSx��B�AT �ŧ�
��3`�H`�q�Q�����U�ʶ�^6i���	�����T��Zf�Bݒ�&5�vG��̵u�LI�_NCG[�~��W�� � ��/��cj;f��)���Vag�[2GS��ޑI��@�U@�;s^x��c�͂K� X�|6ꙍ8����朆w�Й�(����0�ֻ���a?��D�eyi�%=��5HYX8���V+9���Q	���l ���4�� _Ѥ���G�%|��91��Q!XT��K����SPm�H�
�XF��:������<�G�7{�.\</���5��?��f��t��s���!e����=�g����}��'��ַ��1T@��k����C}��_������j��y�Yh��2����X0�/z�|t��$����=�:�W�"Ɨ_�l�ˑ_���+%�[)���"dX�/2�5;l�&c7�_*BlGTR�\v�8-Z�p��k��Z}8>�\��>��S/�6��X�xA!����Rg�*�Mp�M�����$і�xn8	�T�Ȯ�]
�j%������s�~a���t+�q~8'&�Z;q�̕��	�\�wu�Vwΰ��Q$X?�j�{���sb��]N�ц��nv�V�-�C�ќ)�T���k�v|�>z=�D�o�C�~}%�=f�{��j�z�c���ewOyny�6v�A�����x���;����#U�k��>|�pA.��O֜�{��1�a�ka{�wB�ͽ\0�����u�+������!c���񶷽m��~�����A-�o7�y�ߏ��Y�9�X\�X6�k�����.�"$!266a��j��q�m����ĕ��-� C��l�0��l��A�1X��6����=!e!�U-��P���0K�����D{�����l�ji9���o�0��~	�d�x�~����[Y\��k+Z*�+u���=
D��1��!Srm	��X"a�ۨph�n�*$ˢ�����mq�p>*@?�୺V�,~Ź 1�k�9Q�%�E��޽7:/�Z���EC�����-�&"����?��!)�Ta����s�G�\oY�u����P�� )UJ���χ�&�W^�����,�
:�8�Xf sS'�x��5D����i�����}���5D́���ն�Z0����oF��[Yˍ�'P�!�׮�U�x�x�l!k�z6ط�J�=�#�Qsv}���ed���ʯ��c��x]­�5�
�0 �����?|�Kc���ﮯ�o5h��t`�c�A��t�A�z�:��̽�MV��P�P�X�[��4��1���h���:��f�%�ϥ�]X3��C� ��l3;*/�V/-�4 l<p7��<?G�Sd�(��۝�@��Y�7����,�D��`�,�$$��==�a�|��I!�gH�����w��`��
��`��,��-�h'���õ����C�'��$��aO4,K58��xު��.�Fe ��U=��*d��jS�J#.d�=P)jqL�r�Cg~�>G�T�O�)-���T����-*;x��'�<Ҳ��O��?�ܢ|sF.K�Yj[z'�7II	��9�v��0Q�̩�!#kQ��+�Q#��
zY
��_�>��(�G���#7�
h��w��ſ����ģ_��R�Ј�6��j�|Xd��ÍGr}v��X�B�cCW��V�gd��������:�r�"�l�:���'g%�#���І�"Wã%}`�K� -��F�x�N��c� P��<�N�
� 	roX�<?����2�㨹T�H�.�F��s�Z�HC
�V���m �I�ұ�A�M���j�~��������s�"8x�;_$��|(�`��>!�.���ڠ`H�#ű"�D����-,�$�Յ%���M�&KLcUK����	5�/P6l�^`�q@P�W*��t](L�t�U%'
��'�:M����b�[�H�kR������2��G�a=~�K������w�Z�Wa�B\�������<�%�G��A��Z�����C2jd6e��~J��x�$E��<o�GK����2'q_`0���b��'�6{��~y�|6Ct�����QB{�_IZ���I}���5����w� *+vY�]0lk�Y�9�c�bQ�2f��\�
�\�����ZlY�PfI^i��(���	_����֘L�]/�x��Wy�	���`�e/?D�cR�B�3?���w��ќPb�uKsao��r����y�P>�~i�m�%:��E��*֯�zR�v�$��%-�m��z\#,g)ҵh;*]�;YXT~��iz�&��֠^_�yE��-=�ȴ�sGİ�3T�*~���۾����g��/����h��H�
���K|��<(�~����K�μ|1��P��T��ǌ�r'v��{�y������+:����ks��g���n�|�1Oh�`����A�� ����˲��3�������5��}������������t��PB����䗿�h��n��Y�7�zݚP���� ���2	M�ᅠ�DG�HH-��ݻl}�h����
�Lc�������rN�7t3P?O�oll`�]q��:��u��������h�z.�.!+�j١ʄH��H�tR��@��R��<4���R?���uK���� ǃ�>GX*�2��(��{\pc.�e��J]�:�n����<�huTz�B�FI ��`���5�S/�/
MyU�GW�ߕ+s�CP G*�Z�&@�1$'h�xP�JoM�U��pd��O��'V�K���� d��O�s��@.<��{ijȁG|�
/�W���C<nQ����0qs���������4��x�_�WP>x�\_�/x�7ܰ[�gx�  <7��(�Jx�bX�������[�~�ox��������7�����[�#O=�xj��w����laeaaU��~�U�\\s�� PP�J�.-��z������\�m�Y��(�j���o����K�������K���.�y9�S@
�,8��纾9��~¬�CY�ɣ�͗�b�H�0�O�sH[�n�㒱����@�JB��n�¢�Ք� ud��Wabr<Ђ��Oa��������5~ u�,�
��Ĺ.��L����ـR[sT<��4s����R��$�cmNٲ��aG��$Ȁ,����KY��!���S�28G�7os�ls��Nd �K�`���Ð�۞s���|t?�<Z�1/��(Z��J�Z�ya����(�G�@Fk�ڪ�d����j��S���W�Ї>t)��;�
��f�u�������������������B����,e,L�����$���`!�*P`����� ݜ��-q�	� ����/XQ�?�>̺��beD�"�/"�(�54���	Y�����ڸ���t��� �^�v%�W�d�Q��އg��ƫ��%� ��b�$�՚V��A�B���(�R�0�
(*�H����*�3�M/��A�>�C��1w�#uD�8�� � .P%��?B��j
`�lkQ�|��Bl��1����[	�Y�O<#B�{
�(E��}:2Oy%��:S*�1���9�Oi3��`��ь��a7z�<�:P�ơ�����{��@A�|�5~�i�Ў�= \��=T>4�p� � ���R�B�(�f�4YI���ɉ鏼�w}�/�b�|�=c����L�J�����5¹�_j#c�̢��7:���P�xC���b�~�8&0�dF"	vZ�EњWDT����,A/)�0	�1D?a��
_��y��7�D7������[kܳV�pM���:sZ~nʯ�Ea�:Ėj��DD�!l�9	J���0�Ia~�!��~`/����L�n��������U�}��иƿ���=���r���6�=���eG(<���J���� ���oE��H�⬌lח�Qh�}��~:9��,s:쳄�"ч|.N��<�Qe2�P�����䧑�1G�@]:��E.@�oZ�����q5C���Ќ)"��'��!CSQ&0
&g'U*4�P@4pb�к����#+�n��-S[>�����~���F��o���w(�cǎ�3��o�|��A��y�Y�7�F��V�m��0Q�w�a������H�:C��.]	V�V��o��N�9�
��Q�ږ�꣢�8p<Q6�v����3�B����Z|�{]�٣W��Zk������rP@
Ho�?!z��ɺj�6f[��m�f�k,}Z0�~م�JVy��6I��Ͼ�
�.����Ϊ���V�4���T���vi�秂�:��}��L�C8��9��(Ȉ_c�=��8:�R������MB�x�]MK�(�&�Q,�^�A���m���ą^;R�9aJ��vӾ���#S2�(I��p�}�w`n�,@Cm`x@T ���<�,�Bz�$ڌ.�@����YGy
����O�]TCaG���J�k��2R�Vh.y��9�M73���(�X6@�Ǆ��tyN`�P��{���������|���Y������C����Eq�������7��E�[�V��~/� ���a�wn5���X�	4`�id[>{�9���ܹ�UNk���
;�X�y,
Y�=�F6�����$z~u�_U���n[@ 2DJ�!$��|�4����o�XM��p_<W���OٲRd9�|S�"�����j��fs��z���Z�^��9Io�>�P���(z��L
��J�?PT̛0�oK]�=Zv���һ�Ⱥ媲!-%������u�=m�^�._���wou��'		Ԝ���
�S+�m�@�A��Jȉ�����b�-ϓ���fX�!Xc>�����ْ���0�z�)��TY@�1�l��;w��ȫ_��G��3T>?�*�p`�O�93�?���|����j����z��r�=��		��ݻO&,�|�ʅ�Z,��1�^F�:n���"��ڒW�PU�恂�Ӟ�~��|���Џ<a�b�l�5(~�j���Ǩ��sʭ� ����s�Qx�Ip?$�˞���/A�Yt׵�"�2e�B�b�.�����U�T�Ҏ��!���*�lg[a �˂�� 1+������H6��^������̧0l˜��}�@�B(<s4"�S�NBa%챐׋ʑ��Fm���C؍��v�͊U�p"+��y����!;6̇�ѡ��6èl��7�dN�<���X�ux�O�`!gx�-�� ۞8q�xJs��_�)/�c�6���]�����C���?��`8~�1T@��O��������>�裏���U�2�՘"ɴ~��ɓBю82jU�O���v,��9c[2'X]�X�y����'
&�G�*<�2����V��bb�$��&����$`��eRO'���}�\a�P�M%�{T���Ǣ��(qP��8E���(�RG8
=V��X�]ж�
-p8��(��]�$-xd`��y���c�`��Js[a����8����n������xmE%���{�Sȳd�eް��xLB�G*#�jI;��I?z�󌾷Q��3�a"��J�������;�+iu��}W��RXo0 �p�����χaq�a�cd~�l��7��5_~�{�{�(�`8~�1T@��q��w��9r����#�<�H�R)�#�[[��$&0��^�WŲO��jU�
�
�� �Hl�`u��i��WoC-6-^�f��,F�/�C�H��x�<����szl1�EM�i|fsD�2�Sv�!
F��|�������~�4Hr���4�u�#�6ԭy���!����#
�
h�F�+᳤�e�H�HA%���aV����;�׋Z��.�j���{��A��k�=��(އ���Q�YVO#Y�WI�C(5j��;{^Q�P��b�윳0 Ώ����͟7a�W��p(��D-b��UY3V���X(!��3��Gk|�EA�C¶�����h�uٜ�cf�������?������ٟ��C�C�Çc����G?�бc_j�����y�Q0��v�%B��D���"�v��%�փ�CiAx�(�ݲ(��$�
��U�o��Bχ�Ԯ��2��/.j~�C>����L837De�|&
"���1������#$���`����M�����z�	G�`�Y�8G�Z���ǐn���	����1B��,ґ��������ϲg�lx~T4����[y ��
CX$�Ss}��R�ۈ��|	ك(u�=_!�i���~���;��) Ė���Նu�c�ύ^�Cʝ]�vH�@ �J
�
lO@�E��ܞ5���[n�����sϷ��:?�*���������ԧ>��O�]���szz��f�o��A������S�6:��ܱ;(���V�˹X7<ec������ED���H���|�^dk=ٔ��ȅ��/?��ׂ`Ppc��;�ܲ���u3
\h;�@a��p_�Y������_�_�t1��}!�R�{��h`CTV��B�������{��%��u:sƖ
&�p^���es48r'Ű���<b�FG�_oC��W�����V�}�Ph��1���:�YZT�(F�T\����>J	����ۅ��b�*�#�6��䯝��T���m�N�rT94��y!ܶ���|p~P<P@)����&�q�Ƙ:o����o������{��;�s5�zЏh���o����?���}����/��,�ט�w��¤G�Pk '��������	aL~x��b�(�|f�b��@�-d('�L o���sBu�H�b�LQYa��b� B����c�S�`�SB��&���X�s�z�/��b���I{��oC|�X�
��$���s-��D!>�����F,[(�����4+�?;*Pv����'�s�?_��-&Y-ϋa6
s?$�yi%7'�H= =oz2Y�D��� od�=�O�1͘/��%_��<F��ΠHM@��J���a[�ܶn�"�Ƕ\wҮB�]Ӝ�Y3o>���S��{�Ç���#C�#����y��ѣ�~�k_[?{��Z����A��5B$DPm( ����&}M���ރ���� �ZM����a"
\�����$� +Z���B�ɲ_naL�	[@��#��~�������ͣ��Ä�M�f���4����aG{�T���!*��DZ��e�n����aLQA&8U9�=����������<�����:o�?��s�GG�}�&	42����z<cNY�����!��}�k�#�}���Z�  ;�r������~4Ș�<_{΃v�2*��A����^;���F�7r�0�0?�t�!��Z	`��-�n�}��cw�q�~��p�������5�
�G<x����Ǐ�ӟ�����kf��Y�7�:�R�b�,-��g33�V���y�;�c��z� ���u��%�C[w��D�:�R������x��ڃ����(
!��*���ДZ�Y��]Kٷ����1�Rw�E!7�s��%1��J�(�ʅ^�	z��Xr<����c~��Wꪐ�N�&�XE!L�c3@�xd`�Z���h�c�d���$se�,��d�f�M�ߌ�ܿ�ah1�3o���
����O�����'h��r=lF�5�0B�4��őX�/�eqN0�����$�Z4s�E�'����;�㋷�~�%�||������z��w߽j��'��4N�<�\��=*Ň�4�A����.���"�q�Y,W��ϔ2mg�!<�][��I����V�\���,	��;��@�6(�b膃�����-s���c�f���%� ��9���iP����>v�MΑ�Q<g_!���c"wy���9"*�(��	>�F��i��}C^�7�9���x�����b��|�&�����b��ߡ�Ǒg`����A��b�E�1��"Wy�}��h�9�)g=Ǎ�"���|�}�[&�;Hs�0SX�����!��m����aT a��= @x��Ũx�9E	����c~�xI{��^��!���7�
�y�}�k[�zfff�=��c�fa��Y,w����~>0m(	 q��Qb�/���	����Xd���7[��XA�v�G�D,( �Q�c� C��F��\���])�b��Gk�ے��P�T@�r����K~�JQ���?ύ^�UQ)��C�ض~���i��,��MQ�/rr�)lwߢ|r��i�Y�������x�GMv�á��y�J5|V̭�}�Hœ?����T:>���ý�����mv�Y�S��7+�V� ����6\�$����91����?M��K�w����o|�S�z׻��x��P=��Bf����|�;�Ϟ=�N�	�n�:�� X�P*XDTBc��5�h%I\r����0/T�`Z@�+�
�P6
|H�8a�"�4��7[��7F�>������|G��Uh	3T����R�V�M���v>������c.Z�܆�"�\�9���'����q�uF֓
-$�*��c'�e'a�e���Y�1��A����V�@l��+iM��b��o[����q���5XaHظ-�`�L�n�(Ijl��ɪ��dJ&.��IR�#_�ɹ{�F��w���~�0�����bD�`s8�{�|0�0�j� @�P�E��&rϚ�}�xJ�1k��Q>+�p<�c����jEޥ/~���կ~��Sg�b�� ��u;�R�Xv���l P��L,��Sϟ/�>�6=����,�}��In�A�+IA���{E��M�a&ҍ�z���0���Y�����8�g��JE%G+�1)�ب�>aΈ�W٨3���{~.d�� �[�K���X���0V���*�ܽ�(�C�d�ٽ�{�"�.�y8���d�T,�s#���}���Wŗ�K,{y���k�k��o����r
wC(/���\U���@����D�~+y�7v���=X'��WM(��Λד333��;>뭷^9|�p+��}Џi��/����?i&��~ꩧ��V�j��^�=�X�(��,��۷I����l�B�0Í����������7���c�|Wߐ&��nD��_P`��0�x^kP�s8>	����g�^_����;����.�f
�S��@�>�Tτ��Pb��a@��O���Y��#|��%�̽�Vpn�ߟ�L�_�y5���)��'���懲������K��`C�?�A��=�c1F��U$�Y��(t�d��"���]-�?z��lll��^��z]�4(x0��5����,@�[(D�z=PVXWDSZPJ߼.��?o���ޯ|�����6�
��8�����Ǐ?k������b�Q�M���f�m7
(�pT)�h��0d�3 ���Zʾ%�������R�ܒ�Ȣ���T0i8c`;���3�f֭_;�**�=h�c�,&��`���0�d��O��"�����/��'��
��@�EBBI�wm���/"L���R�m&@i�H����[:���G���w�ŧ�PMC��(@����e�j��h(*�z��c�5@E�a3��^���s��W�@��mf�D��#�ꕽ}�&����TJ���U��%i�(ǈ,���X�}�Z�&`���@�����x�p�馛bc!:�����뎻n���-}v�����3?�3�������`8~�c��~�y!���'?��O|��>w���b�����,���ʚB͂/`�XX�����:o�Y�'���ymm�+�ر+`�\�;&A(T��"�A�ErQ�q�Vh���<��%�3/��"��J���\b\�Ԡg������� C"�m�ױM��9��uT|�!��	�*�b�J���E0��
�������*y�1�gԪ�V��]gU��B�9���>�DT��I�Ц9O��^�� ��~�g?��ē�e�uڵ]F��ӂde�F%�@rX�S�)�d�@J61Q�	cp�EB�n�,,,�n�j�D��3/p'⼱>�� ��E��
0�h�x�sܧ��Ͼ�e/��]w���;��z0?�1T@?��ַ�u��ѣ�MOO�K�L}���V�f��&����@�^ �����NMN�eW_��"{�G����'�v��1T�B�b�1��y����8|Hrޒ�S�p���b.$�j=��ַ֓�،	B�(j�zT�+@�o|�����ޘ����~/��K��g�.2L�H�{� ~�o�﬎��5S"a016�%�o�����e1�V��Ԡ�(���P!��q�&BT�@���6�qN+��me�/U�{%^\I�J��*�b6��2�pEBg��P$��4��JTV�c#�����K�[l(6#|v���1�g�����<x���۷_1ʧ�Od�Op<����Ǐ�x�'���y��w��{�����%̇`!��ņE����܀`SP���E���V"X��&k�O��C'�}�Nz->P�C�`)?�\��͇
�53��~�|8G��A��)�)1[}c��/��)���p7+�eؐ�����=�yn���"��/��H� O�������J���C��|��bP`��i�m?�qf!Q�զd2���#���u�Y#�E�,�FWV0h�����NIÇiI�6����3� �޹>��Sb��۷G�$xI�ck���\����c������YG�������Ot�Oxؐ�s?�p������Ϝ�����7�E���%�4�ٰ���=7�����$�����!��7�����z�-`����Z���eST��.g���}aD�S@rh9nN��sE���Y_@Ϗ
��b+��E���2*��$T����r�����^.H6����ϡx���>��A������a�
�/߆.��D18�GJH����[N��3t{m��(���j0�ȒQ_]VV���+sn�aD����9=�MBnxa,..���<��c��tμ�B9�+^�/��҃>���'>�
�2���y���ܹ��7{���j��OE�`����,@�U�����e�K��ːxUv�9E��l����	�uC�;B�Ƈ9g����^��3A�� S<�u��9��B�
�4��W��(���q�:ʢt;r��<���/��B?��\O1!O��P�8D�'�}�V����rהZAiH,�`�QT�rnER�����u|�V�"RO2���� g!���b�(��ey@�^>?�ȼ 峼R�d����=�S��iju��Ѳ-<x�Ղ"���P���'e>��eFy�r�|��1�>w��~�����`8^0c��^@�xCM��O����Ǟx컧�=}xl|�g��7�0Jk�R���^[_����*��Ok�N�X�x�$-
� T�����p�%Q(�x��B�)�䀂(�)(s�����A���C0I�`�����H���sE�R�80|�����p��$�(!�����^~hοF����v~X����>�[�C���}h�<"�\G(��Hs^�y9r���ъ��@T���f%l����xG��� s0�׃��d�C�!̆5@��>�Pj�uż�2
	E�_2�υ!���7�
�6�P��>�ɯ�/�·�������¨s{2Hv�6���:�K��딫�A�7:��b-b�@���(�;%V'�~�o�!�Y������Z��:f��ҷ���$s��^��؄Q�C	
�*�.���j�\�r�.�o�(T��s���>�i��eM
�����7��A�~@y��H�jȪ~z
%���+�:-�t���Z������C�}���{�t��Q�瑆R/��D�K���I�oTj�"B�)�u7��>:D���E��Xдu92G�o��򽍍M�����q))XX�$���rݵ�@k��s/��k�-�[eW�ץ�A����nI�i��ni���ARd��r ���Q����s׺k����}�>�ޛQ5TZ�$�*	�=�_C�����y
�����|�ՠ��?������衖����^S�>�d͆w,p5�L|��H�ψ�r���,'Q��znD�~��UWS+`5J^����5��r}x%�;lNN��&�H�٪_>�,u����AUD!�e�0v�UK��,S>;���@�BY4,���p4�E�㵿"����w��Uٯ�Q��1����z������q��n�_H�̧kTҍ^��\۞�O�S]�<2 .�&gPB�6�s�r����.U�0�[��أ31���^�M�Y�N�Ǳ��t;��f��_���Y�re���4M�r;��_�k_^�C�ן���6�t�}M��}�s�C��`+�塡`1��ܪk��j�d)V��{v���uuu̔�~j�b2 �>�����t<�����ԥ،n�ɒ��!/�e	{���;x�H��tA'���� *�R"gI
$J�L7X vu)�`^��)2�"=o�גB��er��<�(�Cm�9$�����P]� ӻ/]]VB�o+tmu��͍��li�"�njF%�Q��?D!;��԰isOo^'	 i}y&̓���P����<�d�~J���S|xO�.�i��ɸ����5UN%��4�
�yw�����W����6ߍ!W��1%�2[�υ�g�Q��S�P�����HZ�����@��n���I� v"0�<�Xn�&&��w'�����B>��L�Zy����L)�l�&L�0���3t�op~� f����9<=s�׊�)g}�
-�&>���
��(;�~�nȏ�Py��e6��NO�n�Y���;��Ӂ�V�7̣o$H�@O �}�Q�k��֠'�l�6ֶ8����i�N��=�#��cm���!�s�5����k��9���O�xL��(�?���,Z42*��[5�(�w�I�����|��)�$%�����M��u��ߵ^�������K��
y�+&*�QZI��^N�so�y���� ��&&m=�$�V���N�`X=jQY�hR�ֺ�����N�����}����ƹs�ē�k?\�|5+C��j��v����+؀`��e�bs�54���f%6u��D\6>yp+M�7�b�Π��:w���M�=V�GӃg�j�����5��z�gYϖ�,�[�XV�)�b)f�$�h@��f���)���a�»#|oa�wJ�?p�m�MpD�ݦp��N���{���1Xpb�uMs7���9G�U�8G� IM����FE_�u+l!ކ��tm�E��H_c���pP��x����x�=dB=�}������	$'p�~M����u��c]���V�����Fb�����zOi�A����g|�mr�B�\���)c)=��{/zt"}0�Hf����)��ҏx�(bT�=�j�=����$縲�6�R��G�t��@6���|s�3��(��[�`�Z�,����zdy����7fl��� f�W2i��T����[@k��9W ]���y_��L�����U�3� z��"x���hC0c�(��r�ܑW�vn��Os����'ՠ�E��OM�<X�Y��LhPb�C��\�]��ֳ(IeP+���g�o���'j[�ߐBQ��	^b3�0Op��vْ�.�;W���:_v<6�c�#9�
Uv�B�3n�ĸ�j(NA\P��[H�8/Ur��/,����m��N����''�����14�xS�\�!hY@̭�r�e��ٯ��XÁ+��E|-�*_�8�*����eaU�������x5�T�@���థ�}�'� �KZ�u.V��Yc9��s]�p_O�Z�T
�?�-sp�B�C�T�R	����F�.���>ֻ2�}.Zb9X]�^�K�����?�C�?�[ܡ��j���jh/
�IZT�=��� X��/�_����k�E��Lt�L�v���|��;_�}��`������K���|���M*L��у�UV �\,�1�|r�ː��AԈȁLm�~���i��M���z�)͈��eya9��k�Є�۬������\��IRYr|�2?.g�FO���E߹՜.w���D#���Z?�Ì�Ϙ�
�ì|'�~~pr8�s�*E�b���������sp�v�9�<cVQ��'�]�߈I(����~i:d>s�VV����j�=����R�l!t�kA3��H���H7@u�tb!�?^Qt�?�^������}^��RH����œ�����2�"<lA�*&uR���E��?Æu>�(؀6�%��0���wZT_i�䊖��K�Nu��GуfG���1 �{L�x�:��E��)\%�U���g�͜hM;�瘎��R�q ��z�r�Z:m@�\�`�7,��<�B�JQ�F|�e����鏖h�_�z F�5��6��m|��n��@��o��#��μo�FB�eS�D�L���OG_�AD�}*K͚:���I����W���O������7�s�u�
d���+3Ɨ�xF�����C��/�.y�i�
y�qk��B� }9C���/~�R�@�o�O�q�Z`��A�iX)fz�g��BEE�	_��s�%��M��`�·�L&����}��҄��O�r�P� )�����^qr���$ ����=�Ҵ�9���uP*��8��-�xmv�&��Z�N4 r�+��X���!O��!m�~q��m֎�F�g���`�UT�
�g鬽����A�r 株�sq�����q1 5_��/i����^&S�c��V�1�A��P[H��K�?]WT�$Ү��}�$-����"�R�W���.7-���f�Z^���%���sO��:a����`��O�#�?����kj+!�Z9c�C1ٙkt��0�7���Uu'+ݔ{�����/�R�vU:doa��w��IU�*�3O�:8��1��h��͍�IE����\��#^0Y�&\å3������*>P���0����� �����H�����w$����it�Uf�2>�'�'�)M�䉅$|eƹ�k��E2svR�{���iF!q4�}5y�es��&@�E��)�W�o�oL���z%��%����ƽ�"�th"�q�!Aȼ��Fdg�d��9�n/D���C�Y�q.x{�{�=d0�#�y��k!tzd�c�����������zթy� �1z��E�J)�v(���+D�8�d�B����^Yض�Dɂ)������Ǥ���	��;�&��o�A�-Јc߁v��t�6����*�e�/5�B$q�����+�44�-X_ޱr��P��]�;e:l�.�Uv}M"����I9U��#i����Ɉ8�]5t���|]�h�����^�r�ŢE�,�"�������uw�������=�n�x��ܡ)ؠ6�Oë73��<1}�j_�_�4[m�9����Y�B yỹ\!�-�:�Y���NV*��ߖ�KIܙ�㴈	>Z�U�������F�%������iH����mٔ /��y/�[����%G�*�F����X}�B�0���#�I.,G�x�wwx��)��]��{n��_���F|���d�^�6+��N]Dm�X\f편�K6=%4�7�};^��< ������=c�����r�%�I�S>�������J�HH�ߞAt쏜�By�5��;>��i��I���l��$�j1@��~W[|�	��--��s;s��/���Í�ӎfz�f3Ϡ�[�nE�����Rl���u�������	qWm%�0���l�t"^���@uz�Uƈ���#A	`?���Q|��M�3�owu����{M�K��|��2u�D�($�7��mA���Qb~���g�<V��%���-�aL�W|���X�a)?��. ��ײw����et�����"G�hR�,��P#�8_8�Cd@G�%<�0|�%Iu���JgMM:1jO���i�N�b#��ԴS�͜�	���P.�[��q�X2-�s^_��g��"��wYZ܅��1��u2�:��_'pQj��ꎗ�k�듣��wBW��8a�V-����@(�$�V��٨{����|\���߻�������0����t��O[��:A�qy�☢�8�&ȵ��I[n�9J������-c���-�y-�;�7���Q%�$ο��;?g���b|2�s��ƥZ'8���
rhZЦh�$�K
�t4K������U?>����"I��|ô9�Cz�=}|{�z<�X�Mg�g�bt�D�&i@�����N��c�8°&�����FS]S38h��Ds��,a��!��;�7��s�ߖ0+�u��O�@s�C���X�����¼v}��I��6�����
�4a_1�V��Yu�zd}�s���qc��%v�V_����ilT�/�	#�2r�÷z@����t�/�<�)Y#���+�
k\���X��RZ�����µv��� ��n��8�ǥ��)���O�L���j����	#�T����Q��ޣ���<=�P0w��良�W<��jd���e����e���J>��k��Ӣ�u����(�}�`?Z6�Lz�M����4[S8Q'�ˤ��>i̔�4ƞ���|�����Hܗ�LL������.d���YGh ��)��ݸ��K�_v���������L���J��2�(� 9;����l��[���j3�����E����7"���L�~>� ���U��1�}��׫Eo�Q�q�0��F�RSV6a�~0bT��)��s�+��/9,��h->�N�F��#�p%�WcH�s�=#��%���ۅ�F#'Q+�������'�|�#����/t�y���g�����!��lH�k�m> ��ǿ=7�Ѿ��_��t���qn�ڟn��8���x	Ϳ��Xt�&Wa��c韄7ؖ��e��Y��>�� )�Z�?S�ƴr.n��?z"�Y"��ou3���r�
P��+����z��E(޾>? �\|�/�U�Q�մ�#��c�29�X�^0��/EһӍ�s_	�<�5g��̰�|մSΨ�$��J7��h�R��m��\e��S��u˼�W�ц�C�~9�sIX���+A�+��O�/݂���vE��g���(��l�xW���[Y��D����UD�d��S�>~��-���n�6�_�{��i��pz��Z�x�阹��	� �v�P@�#��V$�ՂB$�Y\��|.s�>��MB�w'3��KG˽Šd��Hč�++	�
?Ë���@�ך�1O;��K�)���,
0�n���G�U�0�}I"�¡IH��S���'� ��$�f�+�y�� 
m�RԒ�32���ܣ���RN|H��x��d�ρ�7u�0v����
�&�ϧO×e�rȓ�%�|Վyd9�<;�m�������H6��5����Y���A3I�"5BQ@�Q��?h��/����Ǣ-���^^~�w%U�f����c#��6$E���^���*���|?�R��kfY�Y7�" ]V_�G[�����[Dwj�i��c?Y���m^t�:�Ӏ��.'[!����IM��C&XJ0�x��Z�}uub��ufQ�"�&T����v���L|ߊ������cP������S���$�\��ވ�N�;������յx�,��;�U^�_����T�4ϻu�)U��v����f�cm�Uc��6�������`�e�B>�;�@��&*��[���rċ�lI8���	��b3����=l���~]��I�������9�d�?�
埱��~
I׽c��Hn�Dq���N��%6������	�6�Ɲ.I�����8�NK��Q<e4�è�[m���D	�FZ)��s���w�s��������ȯʝ)�V*�2�\p�x/�w%S��\<���VL�X@&]�o��`�ː����o'[�4}g��Bz�˜�<#��7�Lx2$(�i�g�j�q�����O�);X̷��հrmҢ1
�a�"t?����܌L2`��b �:#H6 V���9�[�u�1�$'�8��U#7"(���wbl
I����Ȗm�%f��ר�'dC�L�x�c&�P?˦2&�\y��k��e��v��Ō���2�mQ��Y�M#'�c�ݢ:A����d�����=���xڼ�����q{P�ۃ�
�z`���� &�5���ψ�%\a.^������]\�e�6��F~��\>�G�㴭�'���R/�S�Ɓ����K(��wvnG����z����Oٽ@�ʩ�+�C}r��21w^��j3�n  ���rz.c�\����q�1��L��T>�&��ǯ<l���a?W����^���l!-���[�ǎ! )�o���zS
��ɅA�����;�5�/o����!v�'xC����o%��7�P7_����m��=����"v�-%�E���N��6�����@'�}n��n��P��;Ğ"�얽�;��k߾�y]�s�L�W$�^OOO�G���E�^��_v�\Pp_;�}�E*��B�q�䗽�@2
z=�rdl�6��A}�b���V�S�7R��Q�7��m:�a�Çl�95�ҩ䄏z|cݛ��0��|����e�d�,7x�-7�:���6o��
Ѩ�|��q�i33�J�矐��qS�p�� B߫��C%E���.���Y���)���י������<����1/谞~�pW^�F0؆��
����5�f�7߭�Sf2@S7^ӄY���H�һtj`�.�o��9~�sb_�����W�?�쵑H ��$��;T�J�R���ԥ���T֔8�
%���_�﫜�O_�Uz��fdiG�����$i����w-*�������]ddd�=�;�4_2�8���G=�R�d,=�$�#*N�f91��o j$2�߯W�|�Ř@�"ɜD�db�Z��2:�5��\�s���9��@���A�u�;9!W}�M��?ӕq �_��²3���et�Z�7��}���Ի�8��<
�V��_�K��þ@}d�ݘ���;~��3�x��~��@J͇�45��j���������@m��$';omM���`��~��H���L߅e�ص�۔fx�e�|O����U}�=c�;����	���O��|*M�#�】�K5�D�i��8�/R㭉7�t���(��b���$c����޷2������c9f��U�)�@o_.�����-�L>]T��j�O$M��c��]˸��!a�RP�ξ�M$.-��{��h��oŶ�Ϝi��f��O^�����$Pi�B��|9�8,j�򲳲��vvƏk�L2ƅj�ż���4�D�����W�o�R�-16�����Z�?�z�zU��8��o�����Χu��Ca�u����4�V���v#��`��d3T�mk�a�bޖb|s����uƶ̓4���g�ӧ(&��~*jg�p�/�χoe"�OĨ�R�ج�r��Rtx��9����]T7�O�u�	�3�_Y��_ޏ��~n���UTLç��wooo���C#}����SV/��J��627�Z3:���Y�N�h������X�]��gx�G�he{�nD�Ʋr՘��ց�h^��虨�+u+��)朊�`	�æ�O��������B����C��\V�H���w�a�n�`��W'ݳ ��!��~����sAX
z�9�J���#̄f��Jg��f�)�A5�X_:�����(+�ޜ,S������������-�W�:�����ܟ�V��{���|�'��7G�i�ڤ���z���J�-�V�n W�i�̃U�mߴ�2��_�D�|��#ա�Ԟ��bf�f�c>�G���;�sv4�R�!mR���
��:G��&Y3�z-���?r���ֆ��O�6o>������MBgj�|���rW�3��>5����)������iob�&�����=�W��ioK�?��n�?��6$�����p{qy||�R4]�Â�����NSWC�m�_�=� !�o�h��n'EjP��x��y{��(Q���߬�N������6��r��;��K���3�)5@�?.�*h��q]�*G̞�,�٥����J\�U�G�b�:da���i���AJ�^�k�Ǚ�0�)z��?���u�4QG��{7	k�@K8��f1z��{˖zH���:��=b x8�}�oyXC�ش��v� oZ��?e:��4�~�M$�a�ץ`�O����6$}ֻ~�����n,�`�@\���r<C�G�b��J�ڥ�7$�-�������a���������]���h��;o:������;Mt8_*�qt�S��ﺾ[�E�@^i`���ٱ�ů������B^��]=!@�����8��EU?�l^tç���d�jd�ڹ��O$:�\��6惻��h��6:�����e?��pO���L��;�߹���=�U��.<��OY-:��u,��,f�A���[3�`�r?���+ Y-ɇ~""m2<B"�=��c
�u�$U��(���{�9���PK   ���WX���� 8� /   images/2f18dc81-c63e-4164-9e24-83fe71d4cc63.png��s%\�-ڝN:�ݱm{Ƕ���ckǶm��Awvl������s���tV��1W�5�k���� �����7Di)q�o߾���la~��������}wQ��V;Kp��ۯo��"j��=^�^D����5�U-U��Y��0�$���H��r�?�E"�~���;E��l�k��&0�k��D졲��f\�^��՜��9|m~\ry�v���QD�xW�	8�,�m<�>徽���x�D�~��I�'
� b!��!����c!�`�Ѭ���7<�5���'��a�(�p֠����XZg��7�Dl�_?���������:���%
�!WROiijZT�%{$Kۮ�2L)\$o�����Nѻ����6�grh?�UZoI �%)��Yiɖ%ii�I桪��|u�SA��Dܵ6|ΛӍvcuJa�Sp�5�����HTt�u�ѿ�T�ho��T����_��H�l������1��3�uw��>�-�ː}gmՆ���/U�����[�m���i��^��qP+_=�<}B%my%��]=+�b2�,9��@C�X!5��,�H�U#4�Z���+��+��:�Z�����	��r�[
Wά�Tewe�a���!6-����{�H��Z�銹����F���?ȥ��P���0�@�vm^g��[���Fz=��>����#���+W7�J[����O\k�	�]��6w\�Q	Ԛ۷�*����V�ڳ"j�}��F��4�[��<�[��Bj��VC	����ﴟ0�O~/>ʇ���)�/0�ډ��Y7��uM[gSlT���������(��lc&�A\���6�;��f�ԏ�h�g^Csu'�������a���io�H�>£���R/?OX��ǡ�K�u>\�!�a�������V�㥕�� ����ʔ���C�l,c��hu�gkq'��;�x�1��ʨF����J�Z�e�{ة��ZH�\@�>&\ ��'|%m��m�� �g�ZUu����������B��z�0�ڽ�ռ8*��JauL�s�@͔^ݒ8�2x�>��H;]��J���F1�?g<)g��b��Rw	��Ѱ�C��ԒW�� w}�޻���޽J�)�C�jZxi`D���Sv�;��BȠ_!W>T?țh��0$ny�3�^��P�H��a�&�U��o|� �o��E$#RX��>����xSG7�����}��
U�[�{f�ytO:��xz�A���#��c�����9�ܲ[�O�s�u���dʿX��l�s�����!�,��I��I3/`<�"$]�D�7A6~�e�����B�/��J��S�d���.+�oQ���;]������;n�4�gn�
�|�V���e-jS*�d�rc%�#%fԏ5g4��~�;F�����Wݩ�+�]W��]��_O�8kȤ%צ�*��''��7����q\ѕZ��]y�ZQV�@z�Fv�(Ң�z;b$D[uu�Xce�DM��b���T���󌔣]j]�L�=�_�Q�vGԕ�h�N�bz��� �O$x�U�!w��5Ԡ9�K��w��ЌC�S��g*�2��_+J�?�I�G�(���Xy��jw糆iXAa�����	������K�d�=�u�'�  R��X���W3y��U53Z#�q״N�5�����+�ʪe�4o�6ʽ
�L���G���	'�8R9�~qB*����	O��`��J1]����?�O^E��G��r(�W4cܙ:g��Dء���>���%�hp�h Gf�!ՈpB/��lM8��?a��蝃�='��-��)iʀZe���4��a��Iy	���ccS���B�y�n�w��K�5~`XWi��vr�����S��<�ً͑_��>7-��	ۢ�̟S�WpM���>U���]^�Q1���W.�ji�m+�e�R\�\DJ�5��e�F�8i�U���'�~�}6:�a�!����΅p�U Nԣo�.~�f�bf���p�0�qX�{��>@\v�ز)kjۧ���0�h6g���������'lh ��X�І{DyF��ǮU�be�"��-,�l�c}UQ�DЖ0���궅�J	>L�R�ҏ�R����ԉp 8�2՗����tx���>��}�8�H'+�ݶc�
z��	iV�5�9#���X�:��C��X�V�Lx/U3>��Ph�.��I	�g�P��>�FUH���t͈(f��k�Dl2��W/��0J9-�b
N>E����s&#�Y����Y��)�޲��YHc���@�54��$���X��=j թQ�8p��9g�w�~Զ����k�uh숍H~>�pp�}yE��q��B:(�r�lY/��G,��u�O��R(v�EXe1��'��KE��Cʢ�	#�#3p� m%�L�x5��]�
]�8���<X؜�yާ}�;�m�\s�di�����6��?�l�N�O�E���v��g,�	�v��ǽo��>�?�`"�I�%����y�3��hE�#:S?$?/WN1 "����4:�15ڲQA�򧼩&�V�S��܌��̳E�h�i��l���_�hl���j��>/Wo-��-z��b_	����c.�����&^�|����q������鎳��hܯ��px �XU��ޕK�b�T��(��wҐ�W�Өc��Ɗ�����s��m���و�ʣ�z�I���[�&ē���MA4�@�B����
��|�L<k�͙�-�?�!ת��E@;��V�I���`,t��A��B�_( ra��ѧˠ�O� ��Y[U������'�AM5l��5�ә[ߦS�%tS	��J8E6�X��!��!�ￒtnԮ�����P �%M WŖc��vl�z��@,��%P�=���{.Qʩ�����1Ű_P�~����&)
Ğ���>���c5�!���P3S�G^Jd�T�}l�CVH�O`{��Clp��fw)錑�+=�g�p�����O����8�_:��ߨ�o��vM>>�ƪ���?�\�խw�\���bF�$B���r�S�$B�U2���B^;���6�����9|A랓[w���?�F�&?��pX9P����ƣ�'|W�^f�:���9�y�������q��^��&�x;���|�:j���c��q%r$Wdv��%�G0M�m�gٰ���z:*ķi�u����R.������Q|��uh�� ��.}>���:^aQ�>zP�W'�W�q�ۤ5F���C��An����/�Qlڣ<y�����U�3�{P�����q�֊�w�)�IM'e
iƨ�+P�o\ш%B��#(�eJ�:B��=��YɌ � ��1l�X�?)�yUj:\���	a��F�B����NK��R��b¿@v�|�L��D:5o�&n=cE~��3.����ga��9���M�z�D,9���ݕ^N�8g�����
>���0�����*����v���9���U�(��ɓt�v#rLN��3V�z�=��I�ý���$�O4���x�W�1��D��ԗdQ$7VH|FpIc�����������;Ho�/�O�@[� ��J4!'�;A������55U���Yތ���K���k�4��/��n�����&Z���*���cc#��Ĕi��������4U��y�[=�<6���x�MFc��.������
�~�t�t]���+�'U!�<���d�IP����mJ�4g~@�zA��)X��.��ɻ�P ��K,� ."lq%N�8
?n�u$��9Z%1�<=����I�TqS9��[obM������M�2���^�]�+9��'T�����`�ϋ6ƞ�pxF����+ӳQ�}�Wdm��]������5g��5g�	v�Pvа���j�;^���JOL(ȼ#Up�r�p'�iL��h���6w!@/`�5Vǋ�D;k��� VYI��HT� �.�Ɵ�8��!������;f�Y��U� �|�Ѯ��}��ova�U_�iB�0�T��ݐ��A�@���h�z��hQ8]!Y)����_z�$E��m��ȸ������u6����"a
E��K��$��^b��1�J���:c�E�f��зr.�ja̃����H,Y��~�1V^���ݩ�OP�GG��
%t�Y�p��2]�^�f��N�}}LG�ӣ��2�ꨬ�&����L}�n�$/$\���IV�,d�.y�K��lY�4o|���K\�}�oo[�g��}=��ǳQE��D@߰�g������9G�e�L4��$�,����^48J )|�HY�0o��+?���N�'��o)��/�x�#a��
�K
��;�E�2�_�|_8	����ʂ�+��9׸��v�"��H^��W���\@_m<�y��> �� ��A#qo�tr`�}�������Ѵ
�?�vޙ=��O��w������e����h��sym�r<#����h�5�-nК�F���EΩ��藪��g���%*��ɴ��F�l�09m֑���!�C�!-}9��1Xž�R-ioB�H�n�;�:R/7�Fʣ��kZH:2�����ڇ���ƫ&�hύE��CM�������3���D�\!S`o=E��/J�u��M��<ʪ��,�Aͷ
kK\i	�k�ڔ+��^J��و�?��yY��r�>s&�ɠc��?�#感��1k�h$E���.5d���)L.�8'�v2�r�a ~�QN���ɽ���pR^�M�T��脞��*�6r�o���6�l�BW������Go��ۣ�����7�p��vPn�Bbҥ<��i��3��1Ie����ͫ��5D���ey/L�{k�OĂ1�/�%��i�'T��wi��O|���i��
�ۤ�Z
�ܸ{����d��q
�4u"KPm��1�#?��Y6v�Uh͝K(�im�����f+n-U�$ʤbj�lݜ0�8��(:�b:Ϟ4[��x+�ArC8c�Νn�b	u�覲�ڳڇ�t3�3�t�f�:��yG�K\��z�f/�m:��&\����z����G��⿊ˎ��G�z��Vp��HF�}�*+;���:�춺��^�i^ώp�������l����
[�bA�!_�o&K�M��I��r4:�K%[�
w�b����v�?d��Ȍq���c���;::��;E��ڵ@�(O��;7���{��X&�ư,��<�F��@(����Y��#n����{=!�7�j ]F�ttyu���B�����%04����ۋn��PR�uJ7*ѐ������G�G¾��!�5�`���q�
��A�����Ն�$&��d�/�	��	3n�?�
�ͶE,pVY��0a�����kf]��Q4(�p<�$�h����m6��)�
P���<lb�O"����������w���[E�醰c�O�Z�<��3¦Y���h��Մ���8�g�5nW�?�N��7�*'�wg�}b�>��4����E������Ʃ1�BxĿ��^$&���`�O	V��`l�.!�M�6��cU��_�1t��0���X߫�-6��f�՞,MЎ�ԃ���˿=Bi�a��p0�|���I���1#���S�s<����.��b�d�P�(��]�|)��MuJ9�`o|}�"��������Ju��a���@�g�c8���x�����k��w�#��8z��v�W�����m�>~�2\���Y]�Y�	�"�����l�ߦ�����O�ַW�=��cO��/]��v� 7k��ӈ�I�f��,����8t�Ytnh��x�%�#"}4�������JqU��0\���wRJ+�W����ll���OB	8�T��KA�yC]i�V�X�h����_��(;�Qn:\��K��QY�����5�����7�K"���	�k����ڞ�.�2kЯ���)K)�|�ԫ�Щ/�2ԡ�
���_��j��8Cx�J�h�e&\�X��Af�U7�M&�?I0�d�1��X��W�7��l����>$��4dAE��bα�~��Э �q�NX�W�ܘ��>��4 ��7���v�P��q�lMK�,�}��H������^���7�,i�c7x��A���������l���&q6�	��:�)+2a�]��qKN,y�LZ1��Î�u�7TV�4�&42ISʖ���|f��Bސ�L�4c:��0�/�<�t���ֿ�a���
\S[ĉ��X���l#ť�5���t�h�����,!:Q=�O�7t]RO{tg����kz:9���]Xf:=3�K�)55�'=//�9�X�1U3U�i8�I��r�8�ED����rtyS�Z0ĥ���������1��y�j��d�t���%��O2w��gMKG(�&��G^E�$Xc.���V�3��?\��]8�f^Kj���"�`j��2*f9����+!=���Jf�5��77������]H8�2#��QUU:����t?�h-�lO<�O�U��,��M*j�>,)L@a�3�ΓV2��:��=���n�$�2X���C�N�`�2��\)8�W;8n�ew���Ʊ��b��Yˍ�n�2�k��4�B����S��s��o뢊�$uJ-4�,��h�^���x��h�J��B��K*8lmk���66?k�uU��bF��?!8:�j�3�����o+p�7m��2n�*�%�ό�g����E�9�SZT��[>@>}���]�<Un�T1}G��>�A'�8W�%������h(N�����Ƶ���mEU
�i⅝�U�4.3J�j�[�#�(�"�_�7bXA�(��d
�Ƥ���D�	E���v��I�3���4�F! ������橣̅���o�z��w!�|w����籴R��Ѷ���3�4y?/�N�jp]���Pz��h{D��kii%��"���/�Z�z����z�]�{~>�e�6��-����c�='uu�}������j5��@�B
%���D\���/��T���(\CAe�f��t�L)^ʿV��×��i�֍b�]]�
	`�2���5��le���ז���U+T�����)����9�g�3`��N����h��ba�"���F�˂�H�P���1�:̽���# �Ȩ'&��8�I�	1V11%��E4�p�S�"ggX/Y�X뉣��0�+�2�͈U�=�{N#鸋�"���R4u����3W��	��B�D�P�V��S�iB�L�;ޙ�B�|O\-��.ߚ3��i����0C��$�RP�u�r~�<��� �԰��D��!�*��Yt(մ]�����ٜ�
�jS��dj}Mz0{\C��Ȩ7��ew��Q��{hӟ��ڻ=��G�G��Gu �����X����"��az��Q'N|�	�?)���F�����6ɲT��ja�!f�n���d���Q���T�ݣ ����+�zm�󲷎�����?�����K-�ᘛZ�`�K!vr+A���ywU,�xVy!(vE[}?X;�E�k&/k��"8��?�*~�.$d���Q�Įī#um=.O
�DT��p�U@?@vܨ�:�}JD/SB(;��wP����Npy>8��_��U�?��q�����not��{��v�������zP\�d�>w�n'/t�m7|��Sʣ�����=+�9���`�KNE��'f���ˢ�b��b��z6��X�S�n`.���i0��$�#~��S�$�^^Sa����QE�����)yy�����'����#�;�Eq)����2����Y��c{�����j���a|jF����H̅r��\�f��(!r��f�)�U�&��8(����f��Ķ;��)��KkT����O<�!��;�S<�Y@�lCJp�'�j�I�	�13%^l��t,�]�߄�(��CZ��ʾ��, �@�yKj9�l�H��,��$D{��*�6,P�]B}��8X�I��ñ>�%��i��>񍺳�RJkցR��	~�y��{������o����t�g�{�����rvZ���X� ���|0 �u�qf�BޖQЄ�J��YGo��5c̵���M�� �E�TE���`)uR��[��|�.1�S���rLKz��=3�U`�Q���+/����3�uao13t���$P�̇���}%���xYZ]���|ݛ��<��� -|�Ua9N��X~���vr�qZ^���b�x��Z�_�ᓖE�㇝5�Μ�x}�/p��{h���Q���ߠ�	w��:������������ɜ-�"����cD�+�a�ȣ�i��j���1�Q�~T���%>[&�\?H�N7&��K�P7S"]���x���b4ݰz&�ʎ^"�7өIdYh`O-
��2�����㋩�.�(�`��"t;~*�zi������CJ0���f��q��9]^�CRX%����ňP�E�ttt&���z5V��I��Z����n-ҡ�ܢ[B�4�=8�DK®Sq���;�G�LĹȍ�XuJ�,5��1�*���a��r.����ޚ�51�Lp�R��J*bB�'K*� X8Ú,2M��X�A�t��
G���Q=�h>S�'>�Dt�G��+	�"S�)`�R3aϕa�C�H� �=�w��i�4�L�V��Z�]�>B�n+���/�2�|n�|NR��a^5����#�H����4s|�ܸ��?�i~��m,z .��]8��S��	�����e�BQ*M)k%ĲO;��%��R^����*2���3�ͯ�:�[�Jt�H��z�p�jpg�1.2��DO��iO�Q\v��Kg�gA��d)V�)���t{�B����!G�#{ب����� �:� T-�Nuq31�����ԔU���hݪ���������.��S�c���|.�3�����f�U���l�iyӋxqxp���j�a�_�歹M�17�(Ph�n����A�M�۰��G�����l���9��2�N�8L:��4隻h�d���Q�1ʇ,�8��YS�^����h����Iz��JX�8kIYT����ov/z ��@U���8�Ӧ������U����B�S�+E�j%d]]��;�x~Ҽo���"�4rHjp6G��@� o2(��wo�LERx"0-�yd5�F����H�F�Lϭ���WO�����W��ǘwy18e`��y!�yԨ���֫6T�R 1_kmK�)!�d#[1��v�G$-l�(�A�-t�1�cH��
83e�/��?�v=����~�GK�3\�Jt�%�E5��J���v�˃��*��h��'OO[7u�ڽ.�b���nkԊ8�3�y��D#�u"��ƶ�_�IX^M�Y�[�t\�ܛD�Sq���%�
B3x���ޕQe8ǣ,.�kaM�o�d�b���8� �Y+���	E�����;�0��S�H��F�up�;�Y{��n�X�+���y��׸�L?�cf ���L��XMj)�F���?%Y����k�fP��V%kfv���zgnWf!�d�أs�H#'xiK[W��*�?���/��Ihk�������c�����ᝒ�������,����+�gy���;�tiǇ���=�o�L��jy&?2W�x��8�=��:a �3c���PF�U�đcRk��8ǘ��
K�lvZ 9%e˛�����*�L0�d���"třixK�9�#E�4�D�m_���<�в���2�kMQ}N)f��D�P�㗔9�E#��U#�5���M����4gaW�q����J���,�H
SuyEl�̝�;�3�!�H�o�����Ņ���#$;s����u%jdf�E�������@✿�RWp��D���У�����:�q�:M͚.�uVڢ:h��*D^������g�ύ�������/�HHc�[����5�Y�r��v��,`ӮQ��@�,��3��ů��������+Þ��<�G���f���W4���q���ض��:M��eo`6���rIj��ל�.�����F�&G%��u~d;N�A�Ɯ�S�G4G������%�/,i�Z�~	��kޜG����?񂌻(�R"�j���H|�?O]��܎.��lc��F��JG~b2v���{�Z=h�
��
ۄgL��3_"�u5X�et��mn-��̲�Gy�
M���n�)��P�m��E�Q����ke�e	8�=3�����]��\|$�q�����Ojbc/C=>!|$�k´QMF�Bb���\�<��݋%T�ZB�������V�ӈx|г�����F��7�]b�ađ<r
�>L�ʍsS��e��s����bIb��U�JT4}�^��4��G�y{AyW��;z�nϦ����*K�4j���$@���q۔��_S-��
�j
�b�w�@S��C��� ��yIbLS��%ye�~5��j^�w�͵��(=x2K����cOۭ`D�r�~��3�������`�n�1R.�-��x߾B��B�L}�S���-�Ļ�\ xm�~Q\���@J�������}Q���~���
��;ϵ8��B��7��Q��{q��_�2N�8�V��bm�,��qy���xQ�̓XyQl
����0���ȳ��Y�н��C�����]�׭��[_s�����ɷh��b#��+�A|C��迍�i�p��n��j�lꔔ��	>�6��Њ���}^�>a��H����ͤ9�%����Z�&�%��e���rrN��a�:���l�5�-�|!�/��ȯH������!��x�[q�V��Hd�{r��4�e�\���* <h�ɸ�0�"��g���q�`Nh舎�a�|�|R��Ϧ��O����&yn�ӻ�؋/�)n[��T��,s|j�[�bu��X�.
�r{��^߫�y�_㛾�K|=S��:ۺ�NvR�W\����K��`V�#�)�P����B(ύ`�������#F��݅��=�OPV�v�Ę�K0+�t���(����Y+�����5�P#�$EC���v=�1�-�<��P��j�6��R�d��@ŎD�Ny������,��U����nGX����@��g���zJ!���4`E�J|��"���qJ��Ñ�9|�6&�+��1�T0P�c���<B���{t�#ON��� ��"�6�] Z��z�
� �e�Z�9��y���$�$��
�Y�� ���޳�y�q'��c�xǿ�{)�"ƞ�P7>��_���<L���wq�ؑ�M���=�Kˏ�N@��H�<��K��ь�ip���-t���q�H6-l3}��{k��}n��v�^b�}�nĩ�3jYA�޳�Y��G���bo�/�n`�0��ٓU�E�JOﰙf&&�r�J�|�Z�ʹ�����?;��o�r�5K���fu�c((j�)tg��j'~������Wz�opZ'�Al�d?�^���(�bo��F`�|���f���a��<���G0E��SZjc|	���K+�@��7)@˓Cr�VŲu��N���fD4��.8���Ua�*�ٶu&��0. ��g�y9D�h7�m�]�,ت�ߏY1�</�j����Od�?&��w��S�GG��u�LSp���M�@����W��Z���t��q�iD�>aӪb��}��i��R�*Pd�nⲡ�b�ˮ���4�i�ζM���X�c��%��Mq>d� ���7�#�N���~eT�'S �Ь���#�� ;���@��	�N��o��n�J�	�ke5�8=���k{�������Q���+.�E]n���v+1��k�g���p�-t����:L&)��0��#��
O0���I���b2����+6A����=�����nY�?���-�K���y�Fq�ޓD��`��^��ץ�,��T���ͽ�^y��WY���%�����v�C�^�˟����Y��;��wiI�ėq�~����V��?j�"��e�]K�-)\�� !��=&!�����g?����/��)8��+��#��kSK;��6�Epg��'EB��ɂ��l�Q�k� w��K���|h�z�ƒ�<X��ʭ@窆�ǡOU{\�C�R�F�겳p�x�Zy�2�Sɸ%+kk���MX{���Ur����d���� v!���I�G����:Y��iC޳�/�ZBtx��CW�)K.���5gAN���n�ZS�I��-6����5	�^�31�#�2��q�2a�A��g�pGnÿ��&��	��5X�a�������3W���A�ټ��I�����'_(�~0�_��i~ly�������;��Q��׹� ��w=�k�z_߄�`-=/���z�]�>�];�=�n�]�HPXX�L�i�<aי�MK��x87�2�$��Ę(��w��UѸ��=/{'S��Ժ!�Pdr�<�I0i���U�B�0 ���9{�������l0l���tx�0SĝC��ŗ�%1�q1�
����D.������{�B�A����zƶVw��"U�e[���c�~ʇ�e����q��*�$"��V!'��s��Q�R+��Q�G%r����I�4�B	0��{şɥ-��q>��r
ɨ�R?����Ѓi b���s��+��il2uBU)��C+�{S�:�d~!�]����ds9�hw��i� �������3��_�"�¬YUvQF��SQ��q�.6]yΪ|��sT�/� ��в;��*Z���?�}��ٯs)~Ձ>��R��M���<õ���kH�@ͮw����ޘ�R���</$X�Rz�|�i���v�����No6�1�U��ٳa ��{�`qe%ՏJ��J��]N�D����>�f�7 ����k����_���]�A�v�7��R����q�pNp/%G��b	&�)r{�#+%�$1�o�{<�/r���+�:�wɾ5���Ԡ�8s����qs�v�W��xs�'��=O�W��-w��_�*r�3�H	z�����й�x��2���w���|�%2���#�y�J�r.�p6gC���k��oU.�r�[Jl�}I�����1�S1�u�f��Q4�BI���Qf�ڈRlt9	������ꫣB���4�f�/�A�M�mѤ�_#���X	@�
L�nR.�����uB���������{�˧Y���
*�sG{/;b���-?��o˝`�F�GB��v�;�|����X���1��7�*�Y����4��'?��� �T���]��ʚ/�
�*�uнsW�],.^u9\�A��L//0�|�B����d=��_R.`}Â��w������C�ʾ#�5R=�ʪSԲ��!�Pfc(��"YQ�u��&���[ת���<r��J#�3��Z���/#)V6k����)��v;������%��pݿ��x8����[I{VӰ�B�
������1���)l'f�/�g�J�	Q@������+�d5������6�29��5@��GC�&^����L�!")
yčv���mt�ch���j��T��׮�����D�+eg�2�3��o�Ƅ�[��%D[|�L(rl#ݟS�
=-�V��5��=�j�cO���	��kůkh��������>'�#���&C����mo(z>t,v0��<r�����(7����.��ֆ8��D�E�t��%W��NʕFj���n6��.G*WCqX#�nb�frjx��Y���9�"�D�N �7�0�vs�k|B���f��X��5���T�������o6suA4�K�[��{�����9rS�	���P���k��݃hm�n
����0�v�q����4n]8^9N���W�L缾�Q��Gm�"G��\���\��L���%�t,����6/�V�Y��cn�pn6O��-ￆ���y����\�ES]�C��A�c�=�4o$�w�R��a�5κ�$I��jq����@�*��?8�,y�3]g
�U�"������s���<�~��D��K���ߔ3zD��{-'�iΈxA�%t�6�!���N	����ݜ7�6?$,{�hiʘyz�y���J�ϸ �m����ot($Uc����r�~���yb�q��u����cМ�^�eM ��q�ᢕ�g���2E�r�ĵ\��#¦�(%���Ln�C@V�f?�>��c�s^;�j�$qE� �/��A<U��ҤqY�-Y�+�"0��V2�u���N?�K�f�`0e������!y/�{����d�H�����7��ɩ#��t�Ұ:c�d�x�ʤ���w���V��\��P몓�u\N�C�4i�<Ib�*X��^J$��sa��8�#G=���{]������UI7���ck\w�hG&�X�vWl&vƯ��Vvٳ�(���`�!(�!9��a�����_����<�={#�n*�A��@2�������$�M�\H������KE&�� 
��d�=v�-�?J���׹���H]�5W�k��Z�92J�� �!�Ÿ�� a�OK�mYPOt�Ҋ�Ռ������������b�aQ���b��1�K�M���t�<c�Ly��NN�R:������aƒ��P|��:�uw?��N�m�&�p"��o�~U�,�'������ub���/>+>8%�Е�)ED4{rtp�Gc���_|��R�.������L���J�=x�T:ƩH9��H�C��Ti�<<���&��s'P���qKVg�}d��>�q	��u�����#��͡?�R�E��M��gW���OD�qXM�OD�@�Ɋ:DxC�
�xB��`���	��x>���WB#~�|�x��ᵞ��f|���W�L��&�u-�b��xbB믨��
�USfD�0F�+aգ?�\�΂�U-e0'Q"J���F-��mI����� w����cm�'=c����w{|�ET��x6EB$N�<��2Iy��I�,{aҿ^:{"I�{r!
���'��mSޚ�Ł�l8 V��~�ڌ�9�-�1���hjxq�IR���Q����j/��岹1�.�N���񵵓+����,��&3�U��tI=�3&ka�ȭ:'=�ђ#���cBS&��~�g���JY�|���U�e((?��{@+�<ގ �,.#٬a��WK �tL�~�&^�2��۲����n���Vx�h���
�u�_|+��D�B����P����Ԇ�p�%%�˳V�Y�0����58�-Ռi��X��'k��Fm���."ҮL5�ʧ?�q����&J1�浔~҈L$���$XOUp3��HYd�`r�����tl�64�,�m��\�~����]u7݃�F�<O�be�zu��P
�D�*��hY�T�=PL�#�07뚌;�u�E��ۀ*�X���Dx�qE��}<Ă8���f��7E�����n0O�o�%��~Cرdg>3��Lx�@~����_�=�"�&��x�J���u�a�����aFХ�O�������ۗ��-Ȟ3T��D���M�[�V9������V�Y�+��~�(e4d��C�ĝݏlX�*�I��D�p=In�|��vԂ����.;{;���pM߶���j)�:>[����ͥ������<<�l�={���
����kWҊ��W�'�Mۀ��o���g�J�?3	=��9���&��M�`�e�N��m� L���T�-9=�N�c[0�$��4�R��ˍ���	��ܣ̇R�x�>�}V�u�\�Da1����5�3j.��9?^��ܭ��a��y	#���o~�_[�P�Coh�����:�� n}3��<v��ZX�l�u#	�4o���(o�vd��T�%7�S�'*�g (0Jw���9x!��(=ȐX���B��&���>s �U� ��,GK�'�-{t���,]�'ʍV�8{��tx�[Z*n�5��
��q�[���j@�n֮6��Y�=k��3�-�7�����������5
˂'d^I�
���V�SI��  �J��1ޠŉYy�p�:�ж�N��d�GV��F<ٕ�c].`�x�N4��g`�9'�hJ��p(�K�*�e�[&�zo5ej7*a)��4�o�R�: @��h������+I%���ț����p���cIz-�U�*�'EP5v/!?�����}�χ3�1��B4/զ`mO8H� 4��\m�[�&�����a�������y�	
����؃W�WC��J{e�-m���H�mbg�P� j.��@n{-淩�.R*��1ȍ<�LFx���a��s�/y���%P�8�aoۈ�F����g��.�f��]��&�/��SBa�����9�7�e��5S��ܱ��pO�yE�)^1��>�k��.��-�_����|�w��0�M��G�n���u ��)��
�r9�B��G��?�c��!�\�^N�I6�!5�L3�tT�d��A@����F\��;@���fěk`c��$~	��9������f:�����X[\�}����Z_\�~����<4c���}������y����ڛ�`R`0��X���H�9��3��H_Q��H�<�1Q+ƓQ�0�X>��(�D��Kb�^ٗ��d�(��˺�7�)�|o^�%��U�����(Sp04Y�����@��=q�2?&��L�'N},���؉�n������6~����Γ�Sl�Wxd#��7�Ǜ����'>����{ۘ�bt�D]�2g3fMkml�H=���,5/j�'�x�r�5;R�[�ƓުA �SY2C��k	)2J>�׆��Y';���J��ɠ̿"�ѿEE�5��n���Q@���}���ξ.(��!jwE��'�4Q_X^±c�1��$��ir��투���Rơ�ox��
V�4�)8q:�9��"!˻T�B�T0i��S��Q��c�d*.͙kBWMr�B(q0��gJS�\�(�o2���mEC:e��}T:s��_�,h�/G�p�����(��TYq��@	m& HO��Ij��,�����r�E�ӹ�2�5�,�H߅�EqnLsCt�J���c��G�$�I��)%A���v�>>{����"w�����3z���t��9<e]��!�����v����Ջ��F�K��St���NN�Ŷ���G��a>��P��o%��/���ZF�,���V"S�ٚ�_�Y�W_^^�� ]�Ȥ5-8���;S\/�	M�D�-1�ĦƘ{�/IGTJ�b�ʔ15FGO4	&5a��ͅ�ˤse�{�_?�<�P�Z�ٰ����f��*���������	t�<;�&Q�#+:F���g����(�&Њ���;b�hT�ql�_�������{\��'��wQK#v�^h��D�^}ND�u�ԟ���ʧ�|��L��z��C3����'.����[#k������P�#���X� �Z6�gD�$*��JY�*�ef�0E�ʈ3zXlR/N��du�喝���b0���V6bLjd�b�;O=GF�l�.à����VF��;�(S�"�d*.8Q�u�&�X���F�2�ʟT*�`ur����c�ͅ���c��+x���յ���b��\9:��/�G�x�²���U�2h>�x�f#ؘ�L����Ӵi�=h4�u�T�'��O㭷��D尻��ф,fH=�#=e�w�r��]�Ӭa]@�"�a��ȅ��,�����&P���6pj��9�>;C)�����a^��&z0
��+�4� ^/�@���4 
K'�؜����<��,}��4#و�L���a)�*��Q�20["E��	\�X.������.sZr��'Ʀ$���$u,�"��o^|�:RU��A`a2؇m��1N�H��LzJ���uW�/�Hٳ�W=��FuZEJIsw����5���z�s&�c�h�"&ASX�u�0N�98���ގ�X-e�EԩSJi��'������>��R��U�אx+�8�� �ܱQfcD~�˗^���+�	��ZN�f���h	Z��~�{��Z֥�9N|�׾����̚�z�q:�$�ª���M�Fo���HD��SY�1e:�L����T_���ݏ���Q�\�Ζ�:�:�G�m]�e�Wꬫ�2<��/��n7ɠ@H��HFѻ.�(�k a�-����i�8ǔ�'��Z� IW	Zw�����9ƹϦ�WY��!�m�L+p_	+����|E��L�+��\E��.�����m�=�`�Ւ�`v�:u���>q���z�y�C3���w�����oM�����pc� [�c&9J'�=I�K�QL��Qg�����r�J�[��đU����V�E�����9m�f�s�n����ņ�T�:�y9����:�F
���)�D�9F{��=F-��O��Y��!����a��+xfԷ>:���=�H�ή�x�9�\y��ۿ���'Н���P��f
�V9�LQ�Ub��vD����/��DI>�↣�k�RxuJ�p4��³�(�?�]�)Ċ+W����B �b0�["�dk��BRZ��R��=�DUu�{}����]�Ѥj�[����1D�%��0����}γm��Z��P�Kȉ�9�@���N5�D�&�qM
���(� 02a�����~=���؆�u��U��y��AlH���[Z�,
�#�r5PQ�".�V�$��ܾ4 �]���Ӓ��n�d� t�!f:XEA�%�(bĳf�C̦Cx>��S�;���5VYF&�\j�!?K�q܃t
m������p��D�+*P�x%"�tDI5��K�B�YrL��Pc���B2�J�'/<���F�K��o>���v�+\ߛC�c\9������҄�Q�ȳ]ܼ����a��O"Z�*L����>6B+�Y����>���_���x��Iч�!.2�c�i�Z���.��¶0����4P �K���BO&Ҹ���f��@�D���J3�4��Lg��졂��F�FO��\~��%�n��QN7�no�F�aA�dߍ>�&Nw������@E���&0Db�P����)7m@Mo�p���(�IN��-�r���:�F���5�R9���|j��ܐ/Ab�;�1�#�H�봱��r�ԅӟ\j-�� F���P��̓��=���ϼ{}�w�Lq8�8�C�D*�v�H��b*]`E>C�̈́vϼ�ks�i�0p����ގJ,�	�92��Q��gI$!�&Đi��4��lin-��H�db$��$�1�z���twѡ��đPŊa��ʺ�A!ܘ�0q~�S^i���e"s�=׿���Ozx�t;������p����[��Y�I*��eÕ41
K	:!���Z�8�$(f��>���c�)_�g��9�fs�`!0f�݌�y�9ﭺ3҉S'����ap(����DE*^2�����B�BH�Jx2v�q|���8�ks�'`ۺ����R��zN""��� �@���!kB�F�\�a|��n���#�ZDM���q=*�A�<��vP'��˫�P�C�C��@Q���&�o�L����aIg���(H;=����h�����M=�y�|���5�����\8�nR�1�H�=�A���c��2BUY�yȃ�f֩x�|	�ñ���A j�d4�EE�x�E�c�)�3�j9G�]�4��s�֍}9GƖ�@c;�la<}�|�,�����v�k�}$�
��+)(^S���6�{�18��xpe���9�K�߁Ocfhw�2R�R�.��.�}�
^|��iv����(���8�w�JJ
��k�b���H��>�5���ht���v�!�Q6� ���Z"��)�2E��)�ؘ��</Y��?�?�Wd�jo����%m�+h��!k�<�������9	�K��C��)<N�N�q�ghr�j��9��嚟��z�9��͚?B�qr�@��Dƒ�s,1�Ry�.�C���=̵��u��<q�=}�?�!� �{��v0����7�>��{װ}0BZ���I���<s���PY����4���q�D�"'M>ƙD��B�4م�+��8ue<�!K9C�B�VH����Z.5���Ɉ��q'��g3�M�3������.|K�V�}�Lg�&VN�-9�l�m� k֟�be1եK4Ƅ^�\M�D�Ifw٦�;��ss�z��뿉c�Cw���4�ʘ�K��¡lI���$���/�DK�0"!S�M���d��c����S�'�h��G�p4J������0$,ݺu��v0�d��Mm6e(ʠ.�QcƑ�\gY����� lV�0Z������4�g�K%d���(���^�!e�I�Bh��=��μ���Ѩ�Q �7g;l7����2G���h���ji��'.3�[q��1!rF(YF��D(O�Y��M�ɂ��RD��<�ñ���|O�vavVZ� h�d��{�1큽B�t�~��l��x�bd)73�<4#d�3�� �7,��������`���х(S��2��K�{v\a���D��R{mOg%�(F'�}��/?���f�U<����8��>�K�}~��	��Y��)��6w�C6�F2څ������)W��UcK�����c'q��"���zo_~�2�G>
���)"Z$X�k�Ddb,�H�Ock�
��$�6���0O��v��G=?�9"�Xd��ɣ��hܸ6�Hd�\��zx;#��U�1B&+�����<�i�2��{�C�S]w�����S�$F�g̺ں���` �ޔ@I�r������[��2�ׇ� ��@T4�::R��H-�d�F���t8�Nc�r�,EX�_�9p������g}bnn����s�C5�;��oz�[_y��m���A�F�{�Bp�b��:��H��������2���o��XX����<ڝ��o���<c��y��i�ݽ����h�
�g�J�o$Z�e�I�8؅ȕ��9:�P-2s�lB�E���r���b�/�@��h�u�fԒ�9�G�@�5-��%���xŎ6�;�ɓrB�Opz�����w�ó�,ڝShͭ���fY������:�=�D�K&a@�cW;�RsĄ�/^�(��݉P.cl%��r��x��ǫ���XYY���L|1����-)Sa>�^��.�(�q����F�,�bT��'�]���No�	��Љ���h`�O �.3�W�n��z�E/_d[��3'�I���T�J.!�J�Fi|�Ύ5���8uꔠ�����Q2�f���"}:�X�,[��� q�G�#}rUY��Q�LF�Q��wºJ�ὄ�@`�ٔd�)�vnbwo햇N@"�\uJ���N0S7�D�K��,M�ܓu?eu�ԩ�r�Krq]mu��8/��*k;O�ܔ�k�U�ח���W�̚�[V�����	�4ǉ�'aWc�g����1qn�씸���ˀ�2�
H�p�	F�1<��x��tv��a��H7*:�_��*�l��e.*�p���e+�_��w�ΐ���k!&��<g��/r�l�g>u��Q'y��%���c�YM���T����Z��3��zz�V	~ aT�-�J{S6��t���ق@��8�&��}F4��ƼLޗ�!)6T�_�������ily���v�:5��t���)�3s�Mg2	�đ4���2k��)Htťj��F��)�E���k�9wѥ��ř��(C2�C�ȅ#�Z��X���4���3�>�a�y�C5���ѓo�w󵷯����!��ڤ����V�Bb��P���޺����=Y��īK��	��$=�[P1�P�L�(|Lxigk��Wnawg��r��$Q�5�(tvU&2��%���D��w!,Yw/�:bh�s4�u�XZ�A{�r�!R(�,Be�j�8٧t*Lnא��{���ǲ7��B�3��{���g���u~o�����B�#Q�-76�g�e[��t#�-��y�b�r��_�tI	��x�5���d�<7d�� !E1ʵ�}��1&N�=�]q��3ywg_����J[���e��Ls+^[�� ���G��. ���+R�Y��/*C5l��!�n�&$���a������)�X��~����fi
���4d-v�l��TrČ�5R[]]�.���@�.c �W��=�hiXh�Ln_f猠1��5���q�;�&�όZ���4���3�w�s����.����9Z%�dz���mv�<HY��3��\]�9��Ld����o!�5(_���������6�W��N>��ǐm�.--��c�F6.�$�ШӨ��T*q��(sF�t�N�<ךb8yO�<Z�.no���Gᮡ�}��#;��O��oc6�������l ��~���|K�r�M�+t�̳�R�B8�!�pd�i�+�^���"����.,�%3xMI�1bt,W�s�G���K�F<u��	�Y:�2@��&5p��Ncks�YTԀD@M]��(��D:;&���%���Ά�O#��s���=k����`�@�ƸXWs��� B8)�hEA��>&R���R�o���GJ�<W��}�э3 F�LݾO�Zq���f��/�9�l��B�L"	��sI�r\i3)����vK䳼��;�x���� ����P��`?��ի������.������$S�P0Y�������ʌ�߿"����,-�&a�)v���Y>�u^�!�,����{Wq��f)��CU�E2��C6��?ܽY��Y��5v��O{�&nt����Y}�˸%�w�����H�$,����iH���dTTٮ��&��"#n�����w��7�Z�^��ʩ*�T'��9{����Zs�1����Ѣ�N��v�]�4!pZ!�UX����"�p���N�s�{�����̋�̍QV^,Q�����d�`·�Z��Q8��Ղ��>�w���J�K�v/�`4�d.Պ�`4�!:����@5�����\���z�\���<�3�+�\�~��$����)�tE��n>g6��0�4��EIE6A��f������_R��2T����*|<Z�?@��v W\U��޴����&���5+3��`畂-Y2� �K��lA3*�x���>��L9�m	0��f��%h�;օ�J�zhyd6'����S?��	�Zx���"�����<s8H�]�F��� ��>1Cy�	�k���{�"�^� 8_T��k��c@���8��s���Рxd�ޠ�|fd�J���{��h�3R�%		�"�,�̆�+%�rq+�R�łl���"%��s ��M�Fn6OS���������U)u>�To����+k��d�G�]-k)���jh���X�O>�l���d_�y�h�l:rR���te��O���&�mEM���<Rت�T�5U���G�>�w�D�Y[�bW�Κ��,�1��<��̎g� ���s�Ĉ$b0J�Vir��h�v4q"q��ف��`�[1,	V8��9���Y��-�}T����"-�W��ǹ��������j7�+�\@pA*��s�tE��,��~�|�z"��l4t�?U�{���i>7�yhq8y�JY)����J#�u5�RBA���a�Q��S�� ��\[;���_Z[[{���?�g>�`�z��O>}��G��?TgcC�.L?�E�$�!H 㐁]lv�riE��~�'Ow=����S
;�wl���ʘw�����d���A_�����=�&&9�ﺪ�L-.-M]����զ����"��3!@���^��B4�����^����J�OCt����Lr�4�F!+3DM"����T�b_��D{�ӷ���%�j��:A3U%5o ^��f�A{��3"�=h"�Ύ?��ή�e	�>H��}��K��dd��������b���g�޶���������=߇6*�KɁ���Z�z�6���R�i<"J���x4��)2�1�3��s�}p�E����F&Xŵ&7�4L��, b*�Z�1ĺ�34�迻���8�ez]�[�~H 8Q� 2s2
C�Y>�{A�"B���Q�z��'��d Ͻ�k-�0�kX;��� u�6l��'�ݩ:�._�����h(OB����H���MF�*����q����b6�P�{�K�!c�)U��LФ"��W���6��pȒ.Y�t�ge��Y�5��j�ۡ+�[7nK�S���կ}Q�^O��`��iq˕-W]���j��]-gZ.N5_�b84y�۪�@U����,�h����]z�բ�{��N����x__�Χ:��4Z4�^�������    IDATEU�}�,)dH��4�R�X�%W�9�2}��r�	�I#�
���" ����s�%8��5�a�2�D�g^�$�|L8;s��Eg���U�(dl�8D�-Κ|n�<�.>CNl�����'�t��<���[o���fh��5�g>�y]�sw&*ӘZ�f�]����ؒ/�K�����q�S����e��_�l����=oY�̺s���\�t����������l�ξ�����{�ɶ�<�ޚ=X�NN�:�?��'����nG+�����>�G�7���E���J�����K�7Ԇ$U��?���@O��ѣ}��?La��Gv`�-t��^z�VW����J�D�Ұ�&P�PY�9�F_湑��T��������C8�}��E��a�����ȼ�*�O����_����P�����H�eQ�P���((�Ž����MYy�%���"�~�T?��O|���oR�8v���E@��@��g	��̞`�x�h8U�
��ۼ�Z��R�G�m��U�\���%uz=WhTk��Ȳv$�4�Wt��<�*���q&%�L�΋� �>	)O0��Eϋj�`��|�����v!�W(�"/�`EC$��	�G�l�l��m�g�g�y�%6���_�ו}k��iTD�o'��z`,#UO�9�w��	�a�\���������K5����DC�eg:>ڷ(�t6T�ϕ
����+C����X�7��i�uDnh���aR�l+%��V�Q���z���hͦQ)rJ�]m޺yS��������W_Q���Ӄ���64���o�j�t�S?�X�J�3-�c���ը�]�߸To����w��V;muZU����zE���O���vO�-���.��ZQ{}��c5�/9�8`�B�����,��x�[F�������&�8/b=gr_��I�6i�;��3��<a��u��<&����O����7�E�J��1���o��$3��_�hw�Y-�S
�	b�P��p�a��� �彙�5���F�n4Y^��(&Np��c� 8�a��N2��I(�v�C�d
�H69W���%+J!�����JO׮\�O^�����E���3�k��?;{��w?~�����vVT�7�������)4#�ʥ]����j׋��?�'�>��ma���1%g�뽖�7��|eݎ/����N��w���ܣ�sO� Z��%�]���M���-����#���&g��I-�0Fb�@}�v�p��`D�v��Q8'�+3V���l��:/J{�2W�<Q�p���P�'ߔ
[*4ֵ}z��|�FuŔ���C�p-��׭�KU;������&����?�0��U���ֆx��l���X���چ��b��&X�M#��b�g��ve��m�t��CB�u�kBBs,�`��w�`�(U����=��|_sФ�K5���9�Q9��bl!����0E`~7�A��&�%H�ʓ�6�a�ǙHr�L���1b8?�Gs��b&��%��BRU-�qd�^�|�� �q�����V)[�	F&�}fV!Op��V	IC�J
ؖ�?���`���_H���N�#�WKe��#-ȉ��^p�M�����A#�3������f�������+f�'�~�^��j��^�x����'��oڄ��_�����U�� ؎t��C���X�©��h<	�4�R��*�ڥ�7a�Sf��R�m222�Po�j�T��?�@��H3p��P��|~���k��J���ό��ԪʉB3\/��h��,{t��G%���*�+Z$���^0��Y�X�y�&$,$?��Y��?�܉	�>'L8�8���1ߞ����z�z�Lwق%�'`�#�l-!=�b$�.�D����Cߞ/*c'#��ˋ��B!��4*��B$>z��ޣm�+[��IY{��+��{�\�{�$l;����{�����O��ȿ��������w���=�� ��U-J5C�'�=}���y�a�Pҍ뗵ui]+=���������c3�	�k���������ZK�:Y��b���G��=��ޙN�&�M���h*[�Lp��`����#��y���5�,4M-'W(�q�`��š��X,�J�k�W�V�
��gߓ��r��$o,��H7��L��P��L����o}���7�����<���>=H�C�#���pH��$,��������w����8z%il��;f%�J���/�N�����
����C������Lm|p,��[�
o���T�~.�����j�m�PW�_����e!�H�/�b�J�@��3���]-.�a��� )4��/�� ����H� }���l�@ܗ*��ȿ�*��<�������	�=�¸��ڨ\ �E���f�����X�ӛk�5� �P�5�.s��M"�r�3Ѹ/A���>�0���C�E��`oǁw:�_Hx��d�,�u���j
򼎭���~���A�A�]=��}x	������VǑLp�cr~r�u���/_�ȯ�|Y�bѢ�Û6u2.�P�b�k��{:��T�ٱ
�s��&YZ��c}%UjS�����|�.k��V�^R�Y0��Tmi4o��������P����m�m����s&���X�L(;h�Q$L�R�I:�.ݫ}� =�,r�
̞�E>y~�?���<��8|��:�$Q@�)�1�8��	�&Aг�H��C��ݞ�J��f��jΊgDP�0��E/8��\�33�ԲL~��]��Q��l��i�xu�7=q���e 8ۀ�c�����4e�bn�S@�+H�b��D��(�_��W����?�g>�`K���O����#W�mf)�̖:=X{x�w�D�q��U˩Q�l�{�=ܶ6-?	vO��֬q�lU5�m����v�����1*;E�q83�k��5�Ƶu�t���X�ؒ���t~6v�M al(/.��L�	�$p� t�T�V��8��J�����A��u��ly�r�X�W����������V���������*s����3l`�jŌI��y�-[�=z�H?�}[�e�(�lT��b7s���R?><���-���t�F}�,���b����e��]�&T���! 9"B�#1(EE�G�ר�u��e��I$8 �9�����n���s�ъ�E���9ԚBR���u	����D!��0������k��*�k�|(���N k�Є>�I-��FV"8��C�j��>Z����\%�v�s�-���L��ST�B��Xr�q027	,�%c/Z�j��b���{N��볓�*e��ЕA�^P�=���{���|��J[�.m�����ϭ���Vj�4íe���f�M�_�c��(a��#!�s�E<Nw�W����ك��k^��q�nhr1>�Ï���}��'*�U*��E_<ty+��.mu�,��hO�YR��0�kľ��j�!I�U�m���}��ɱf�KZ����ݐ�$ha,�	;2��r-�9�l[N���U����b�x%�DA�<�`Ԃg#Y@�N�1j���&k,�R�L�cS�x2�p���j%���\
Ҝ�8�$�
��0�Y�C����k̜G�62������aW,��1{#�Bf~�~=��D"���s )q� �ks`䀯��h2sɣF&=7�\@�-�D϶��Uk ���7��T(\���?ǯ�5�����{�~��ɞ��C�0�i�\��?h<����荇��ϓ�[v>�R@���ˊ���벑��'g���C�<_˯�Z�3���>������T]���uݾyI���Y�(,=|�X��:;�Ĝ'ݑ>�Q��q2k��9ż$���4�D/�E���S H$���<7����yĀz*����s�|����胻�|�Qc�����FjW�Aϟ� Pq"K`�#'g�(�Z�����w�g�F��s;�D�b���p����PÂ�X%����YS���tV���mm��tʆ����!Z�u���G&Hۑ�b���tO=1?��a0��ZN�Y�G�$������E�����*�ϙ�����cw��_m�ŵ��#*ѓ�+�TQmi�	�m�G�9��&�*�+F`�J!8���>؜`���מ�:�HDz��,�9m�DvIs�������r�v��Ns�Ǆ�nQ���J-1	Xh�3W��
�ۅ�7:j7kf@O�#=|��P2Z�^���$���40%GQXAFϖ�V5q͜E&�E]�tE���^zq������`��e�fE��R���~�����m�P<�!�G��%�tc���a�To��1���ޚ���|k�U�jK��^џ��~�ӧ�4oj0����hu}�m�>�*%T<C���Z��^`V�#��ӳs�jUW�$)T��&�q.�ll�G�e�ӭ�E3d̓�o
�v�0���?�SW�����Bk��J����c؞�j����x��dd�� �FŞ��R�NVz�3M�X�FA|TJ:�|N.Ir�~o�w�e�ӓ$��� ���لǀ�Mt4b����	(σ���|w����fK���W�����J�3�9~}��v�����{𣧻�:�����<f4{� �1	
��:��
���דǏ5<����F�m_M\^X��sΟ�X�n8�k</h0��dyZt?��t��\��BW�����k����>'���<���{O��s�q�S�:��-�A����G2"8�(	�F<df��b��W�I��
�3M��c���f�JeR=�с�m.��/_������k��Rs��T�g*�cp�*��n�ᓧ��g"nv�HVzY�>����E��*;�F�G��\$̀+��o��5&�,���ݻ�ɔD��[�^Օ˷5.uڟ6��uχ�F��"�����Z�b�&�5=>�5�@٬&�d'f�K�%�8�0!�ѷu�^L=��ly''�~��L��B5�A"�2Y��/{���y����T����D#�0��h��+9�ġ2�n_���c��jk��>gט��c�5�<����څ�u��Ey�D��y�L����^�}�^T�h����;�T-/�������с��Sk�$~�0�������'U&�{�Ͻ�j��ƈ5[е���V,u�ֆ�6����#���4*�ڑ���сv���=��T8Q��9��|'m�Z��ha؀��\���׻j5�l�\jQ��M�����R���a$nm}�m�=b���։���� /���m8�x�?�Ē���g�^��ͨXN8y����%��U������'��,���N�h�䗝~���X�qfe"�]�R;�3��`��D\J�[�<[�u�J�ɳm��ud*�Xp1`�\�0�]�Z�UG,��G����n)�vr+������rz�K���}��tz��FS+�6���/��r����s��q��_�_��vw�����O�;�-���hLO ���z�,Z�w��A������"	����Ug�d��<��C��޵�9}.z[�����>"dFf�a:\Z��VO/ݹ����g/y������~���5A���aRYa1DO%���������)��Uт�fZ��tѓa�r(�o�f]B���ED&؎G��\�o���qx���,_Sm�GC������y�
��ս��Z�D5kW�b���d`>��ѩ�y��q�y,�yHֽ�D��ل�a��:^jjw7�l�i����\՝_����Nφ:=�j<e&5�w�a$Ţ��l����_�HD��QS��٨<sW����s�B_�z�Ez�)�&������d@Oa���x��.HF���J�Z+2�A���I��"�)_a)�d8>��FEQ8W�E+W�������l
�9���hR����q<�ٸ>��Q@ٞN�������L�l>�l���֦XCXt� 19�xt�f����͍��\]�t��ӧu|�jbc�B�/\�����rH�q����FI���c��C۰ݸ|]��P�ځ�^�j}���xW'�K:��4+TTo4t�����j|���鶤3Uk1S�#s`$_��T�3�d#b�:��uu�u�q�5��6���ww���~�j���������kk���ؚ����"A���R���5S`��N�Jvz9H�����n$ey�D���>s�)��ٛ�fB�A�Y]�S�Y�6������ܽr��3]v���	|��Iv*K
i܋��!�)	�O����yA�֛e
�)����ovb���nʜb9Ɩ���hAb�]U���9�@����}P�gH��BI�Rɕm���K�o��v��*����k���;�������ۇ0gj���L���27tq�^�<Va���+.4|�ڷ�li}c����q>!;>>:"I�c�b#�X��Y~y��6$$�Dnݼ��UFL���{�����]=y��L�������I��'_��5��F���`����͟+��wu�o�	�X�&	!�q���;����w�����B����u�-f�;<U���|<��J[kk���7�����Z2�p�t�u>��`�P��ַh���p|���Ԁ���.nK0hޱ	9\WT��2^W��VouS��^7�9���U��z�/6o��L.:Yn1����`��c�Q�020ߣ�P�/���l��h2�7+�uaiƲ��Q�ED���ڪ�I��5h�5�=���0Énq
�����T��4O�p?m�@�!	9W)3��|�沈�V�=��?[`J��v��{R�u�q���W�6^���u�m��<O-��n��e�k:G2�F�|����67V,�_.M���t��F�s'*lhf��}v����i���?c�H"�{����my��-t�����m����O�u2��P!����LO�}��ў�����6'9N4"�Wt�RG�&F���րg�be�jk�Z��R���>:�7���J�+-�v(kt:L�����M!�n	�Er�J�~l�D�`��Q�]�ZXu�	d���(�y��T	�'P��3#�����IƌL��!)��\k��=����'=�|�9OB/�I�����7�ϕ�mN�9k�x�{>��d��/T/�]�dc*eFي�l���;����k��@1�^/�����E߻��Ҫ�L�BI
tq��=x�K��,
ь�s��\�����[?z�mi2/��~���d8���{��y[[Qasz��p]���u�7��[]�:�4�%�����mvY*�/<m��`m2�Ǹ��҅ɷ6״��o)mo�꓏��`�X�1~�!������Բ؀+�Rn;�K�ٮ���ᨒht;�ؘ�L�Ҩ���z�Ԓ�gj7����_����ӟ�\��5��R_�&j�ZZi7�����3L��:><
�i��	a���>><�~�;�<l�&�`�P�R��>�ՍMǘ�
�)�T.m�պ�jeM�:P���/��Vbd3,�TU��	��L�"C�`����C�3�Pr
X3��м��JR5g��?E��d�K.s�u�O6�V�U5Ϗ���υ�H�.�O"^���#�ST��9P�g�+Aw1Oͧ��MCw62��l&���r��WH���!��z֢�T��w .�pD`ϐ��`�×����G#�J�_�H6�-��B?�N��v�h�e�  ��b���P�GO�t��f��ץ� ���	��IJ�A����d�`;��
L��jθ�w�s��M��u�&&E�Jg�u��]l���~���i��=�TP�Lc��<aߎ����U��j�^�+�a��v���JI��Ted#K}�ɱ���O�,nj��jQm�h��N�٧���J�qIḺ2��H�i� E�v���s�l��X�<�ǹʼP�J�s�9<��%�����	3��L�+���s��`e��k6qZ�m] G�fe6﮴o��R�ͣ8�����,xJb>��pȌz�2��P݂��V�|�IV����*/K���������^�/ɴ��	���h%W� ��F�*��ѽv�ї��E�m�������l���������ޑp�[ݸ�r��Ó��������ƺ�V;�s����ybG���am�[���ىHV����p���G ��&���'}���
��    IDATd��x*�
��<}�v�i���S�c'�6�@�� %XgH%W����}�Yd��ć*'m/��w0|�!� rx���|�_,�U������_Q��~򓟫P�������D��\�暯�۬��ұ��4�f�>>w�����#O��g{�>�!a��@��l��C�-��"2w��h�n�Q��z풦��*զ^|�ݸ}E��P�(��a^HP�ҳ��a'��L�ǝ%�Ph����EUi�W~��Ȭs�6x�� 	4mVwѰ�E�M:�9�xB��Î+��`h��x���:���g-o71D$��I�\]$�����I�U�:sb�̱�/'�v1�~�ǁ��(�D+�9C�U*a�`H�ڤ0�{Z��Z�8����`�S�(���ԂlV?IYY�FYW�����4;~1g<�DG�Ou�lWW{j��=� >@���s���73��PN�o�f�cL�Zt�B��X-�ҭ4��V?�+/]1\Xm^ҬI�&E��^��o���g���F�#�zс6��2n���ZK��[jT�����n���+��]"�/6��G'�ỏ4_�4+64�5�1��j0�����}E2/n֤l"ibW+!CIki<]���cy/��\Y���ps�h^BRN�U�aפ�����Is�oK��=��S��d<�!`sO��t��fd	fz�Ȱ*��D��@��޿���C����\h��y=4����8��}��(��$Qc��'�}�F)�{o@�5G�t�?�"dD���XW�� �Nr����~�W^��?���}����O���ޓ}�G5{�*W[:8�kg������X+����cD�����;:>�`��,�`֝�^&���2[�a��uvr� ��hxG�m]V�hպ���.����,����
tba�̒��������7B�Þ�� ���B?���l^��p(�BJ1h	�z���׾��َ~����P��Ხ�!����$)8\з������q��ݷ�!w��P<����H���7=�}�8@���"����;aE�F�G�q!?��Z��Z��p�̊�x�K�zc]�ѱNώL��"�*����d���� ��D�;Q��x������%,�Ҩ �6T�<_�WK�l��h�{xv0��{�)�0$���`>��3�{u��o���ȣ41���:Y��S���e��ah`x�9,�*�"+������N��i�	�p����oJ���T�:s�E��$&�H~�-](���T ��I?�h�����ǩ_ 1��Pם��ToP�=*3��i-0r��xL[ׯ^��3�{��bv�67�{��s��з�%�n���m���'z����P��^S{�.�������?����X�>����|EUAj��p����z=ie�ι�L�o�K�7�V��4��.�z���6Ng]�0��N݁�d>�E�����$+��V�v����Ҏ�'��\��,��d^b�4ɍ�f�lr�Jթ�sZ[�2�b?a�f2���L�_F�SK��#)����EAr�+<�A�	�|�P��q�_�Z�!i	��v3��!�h�T��_�� ���vm@��DOַ%`�5a��X8<�d�#!�x�� �l+!�wS����߻s����.�no����>{��G��యj{E*�ut6��щ7��J(B�W�e�%�Xĺ�O�qQ�2O�!��(�v��2E<U��}`KL�B���9���a!�BT�b�#�<#�`�N���N�*P�c�j��:E�����;�9�<-n�K;~��_!x~��(�,�����ٮ��+�z�x����7���;��H���k�9>���4���@Z�����A�Rh�����	��p�-)T�rO&��l��*�$��k��0v_,�a��Z�T��kp0��^z���4��?��ҋM'9Q��tv��h�c\"�L�
1�j��p�u�4�ϩ��0n��,�(Ȝ��x���� ء�$�*�,��l�
H-sx>FG
i�'Xd�A4��ωT�q-
�d;9t�[.Ԭ2�u�`k��FqPf7��d�h�}a��aȿ�$n�H(聣%��^6��>��jN�Nfo�+��'����u���-#D4�
�nl�O�lTu��5�jGd�^��������~��4��h����%�~\�+vNe&f�ް��wT�!!0�u��3����l�O����Z��]]��+�U�,a�2?���?}W�������5_T,�A������U)B�*��k�K;`��n+��
v��m��R�j<��?~��h�P���e��!�P�nf5d?>똙l;%�,��pש����'�������m�N���,�m�>�.����5�Is����!c\������x����3yŴ�f�f̓`v�cj���V��FCB`R닿�}�xV�à!�-�'���h],�C�O���V+�|���T�	� �S�: 9���|'1�y�E�։
6��aʄ@M�y��Q���woܸ������~��O��}�3�;{*ԚR����3���&q���-�)c���o��uB��Y�Z��b�ˇs�`���f�s�Ⱦ�&NO�U*׵���j���Au2)6�e쐻ö���j���Ւ���K3�`;Z�y8 [��E�Ep"�V`N��8�=8�M�/������f�aQQ3��8>R�6�o��kZ����7��j�����x�i����pb_^���J�(�Z2o�.��:�������-l�L���6HR�IU�	@?��t�;��6U.�i�l�\�B^��Н�����p��gY
�;��'TWx�f�� �P��C&,��;�)�.#0�zGٍ�{�Y��X��gL�Yo�`Wp�d�Q��kZP�d!��A�
�RF�¨jb����p�Y���=F#�N�TŁAK��u��Ledy����C���?��e?wNK���pO�G��$���'�l$%=�^�`r�O��­h���M�`A�(Iǂ�i���--u�ʦ��l��Ug�h��=�'���Ό�������6*�����=�*�0W��F�R�VO��Wze���:خ�zj�.��������tU)ڳ�ho_������}�y�MC��yz|�Y,�}i���#7k͔-�H�m6���^ok4m��?���H�U�]���Wg�-L�
@H"P��y�
��.�IaZL�3#s9r JU0ךIL9�fd$vs�ڡ���ל�9�4�>?��s%i�;`�K>{�5�ϑD<��fw��ɉ�ǅ�$���/��`S�x8�-"y�,�^븀�����Y���:R�U��k�͝��D�wplH3�z�m.���P(�[��U�W=��v�B�lL .�͐���	EF�њ]��zk}}�������_~��'�!����)UJc������/&�3�4��?8��ٱe�2y�,;�[~�i��=9>teB5������~uK���`�rp�Z��ɥ��?�p�����7�x��vux��>�+�x�!�ѨX���&3;��
�4c�@�ٶ�~�-y-����)�镊nݺ�9E�w�`P��?P���_��_Qqz�?���R���j+W�ɓ�BK��XUg�R��PB���T���J�#6p,��Oe������tɒ0�Q�2�PM�j�(��P�Tn{̊M�uyS7o^���pt�6G����]o^����c����8�3��Ts��6g��|�$�o�g��|���!�i&q��/q@��J���$��P���s�Θ/��\�һb�(�n{x���XKC�A�\��`�+�ܻvp�(T��8��Ę"زv�~�3�`��V�3�����r=f��� ���Y@��@�V}T$�:RaNL��xu���@�9B4�:9�C�6ħs�Ҽ��&_Q�f)���9����	Yn<I"�ǌ�-��/���l	�o�~Ǫ?��Z_Ҭ�����I6uN���������\��:p�j5���:3�K�n���Z��Y��J��ҍ��I��bC��C�Ov�*�V�n&#C���*��%���"c��Σ?$�La[�("#B�Bv�s����=62a���j�!,	�D4��.ƽb�܉U��٫;%�[dlML2��Ř�}��n2�u��2��ѻgLdO�m��m�m���Oςmm�񑸛Ę�ˉꕅV;5m������vu�c����ٯ{4/�PF�gc�r�^����X�`k-�FӺ��D/��MT����k/��;����_��Y^����o����?��ގ��E���Um�=��~�Ȕ�4����?qi<�Go'���є��B�cX���z����~��fz��u��U�n�`�¢��^��{'�����v�\�n���S�������&CD5j�Wc��F;U�����{0 ~Gg}�y��@�&�� �"�0A����3o�˗/;�f����ݘ��˚������:+���~S�>���`�f��6~����g$���#�L�-������9U�w��]��N|�㪏({�{̘UlA�R��b������������+�|y�..�� 9�P��z���� ;Q)�=��F&��o�H�`��c�4�Xy���ΑXA����r�5Q�d�!	a�ڪ����A�[��4#��b����^�ٿ��,��d��g�"6���r��6[)f�X�٪�	J��<l���9�Yau����9���䮠��,�����t~����^�Qz����To�u��Zu�����qo<8���JŅU���W��o^��#QN�3��ؓ'g��*6��I#FLi������2�>����N�Ӛz[oi\hk��8:�$fӉ���?�g�~�b��s��N��J���f[kkܓ���.b-��\�n]���������~r���ʭ�(�L��}�Ao5�E�xF=�g�;��s(j[��9N'H��X7&-�p�Y��-J�r&.��X�6�-�R��3K~���(5`����wb�o"F�r��F�8y��y����~�\�:HO-��y��}�g���bb�r��VY��rK׶V��b@z��j����?;��|��yAG}�[C�jW*�\��l/	���0/�*�� �S��QG���-�v���n߼�_�Yb�/�=�k�}�d��~��ӯ�hW�ǧ�3#�+F��
lׁ���P�~�}M<�7vkb�4���e"��Z�'�p�"����ƕ����W,�#��JO�s��Kz�w����D��5����)嬛��d�.Dٽ��J]����r׺[�!=Y��.�&HjD9seQ�w�i]���+k�\�Z:�X+����o���َ����Z����=F(d�Ta��F��4�Xx�,6nf�N㐆�������w�����)5~>غ��P:>m�i�*VVT,3�ְ���k�zu�c\�J��3�?�ې�3|i�ڥ+W��ی�Z�����[��͌ݘ$1M�@~�1���`��`�j4��zV/UI;�Ƭ9���|��9�/VyQ�P�"���҆�[�����l�� U��T��F5�����q6�X�5���R:>�6���a� D�|y�u3� �]���( c`C��h0���ٱ��,�hiL���xaEY,.t�rO�N�������%�mOu����2�~T�T��gH�����c�4�sX�e@���&�b���k�O��d��z��U��tr&m]�UMK=� fcfCS���Cݽ�c͗��yň��rU���Ҕk�-���7W�47�&r��t�E�\]���X�r��{��]-Q9sЌѯ��~Q��!�@:��,�rJR�=�|Dp�T�ه
Y�O��Q��h�+<�|&��� H`^ǉ/`T�;$�9Pɴ�b0��;�/;�������S�ct2?3"�+ڋѽT�g4$����T�$|$��g;�q.�w���_yK��nh6>�Γ�n݄��23�e�����#���T��i�Nu[(h��rlQ�c����Y�G�m7�n�<��������{�H �����l?�����m�������R<�u:8�����)6��c�ր��	�C ;�p0ځ�hx�_��z�擾6Vz��/�ת�g[).]A�����^��p�w��=zzz�,��
Yp��0/�t{F��P	���/,�n��k�/i3���T����!�0B<�a�G�,���x*CX��@i }o�_�+o�8;�O~��f�--kk�>>բP��J'����zjDnշ��(fU�:=>�����la#{󑸧�(G����Z�N�#��Rq]�2��b�nH�_�k׮�Ǵ�EU�W�<F��N.?|>l?%fv1��w�ѓ�07cW��8��m��b̢�`�A����T�ANlߗ�%\-�'g֘ǳ̆�ʰʸ�{<Ahمk �8�.��%�,�'):����Vz����r����X�J �`�w�{S�s����	��#V]4Qd��UQT�Yc���gچ���a� �p� �S����f�g�X���"L���V�]6�rv��F�1v�Œ�����[��l�W*[~%��>�&��G@�=��� +��K#Bۯ�����O�{�~�W���h�K�S�_҃'6j �l��#��'����C���JTTT�ބ��By�zc�v��f?ՅZuf;Q��YEˎU�u�|�O��{2V���y 2�\�+9���$�Ct�S	su�(�I�)�,�Ņa�s��rd]"��`��W��0��E�Б��I�����L��8�4�@ӄ16�'a2��e������M*�A��X�!q��Xo�}90r 6a5��hK��3����@H22n�R�Z5��/���W7T\N�����vT,T����k�oke}Ò�}vO{�g*׺���T�45�0����&�rH���f\*�:���z�6����ҭ��?K��E����{{o�p���\�9{t~��;�z���ó���Q�z�é�7�QcbB?�H@���q��3i��>�]��z��֗���d�l�Q��#g���X[W��P���?zO�=��d��V�=$T�X(g�����}M��Ƞ�U�RV�m��[�ɏ 3�pZ�9&db&G�`�3��Dt8��~���]�R�/����'O���O5_^r�}�wh��j{�=�R7�MlPf��O���{��d�lh����s�칂L+%�p�9H�a�(\,�ZH(6U�D�-����*Ǳ��KRx.��>J�o��%6c� �%���`h��P����ru��9{b>�3z~C��Њ=�-CН
'�9���
����U���t��C�]���y�綷w.�u�&��tJE�>�<��[��\���|0e8=�������ID�gr9'�I� ��S�y��� ->z��֤�&��>�S!����$1V��o��S�S��iՐ8횉ܪ/U+�u~~������W�\2�L�1�QO0e�?��e$������F��l�$���嗾�5W����P_y�:�������%k��٣}�H:� �������'{j:9U���R�J3z����u�Qu;X�a ���v��h+������'�;.i��iY��?V��u~�$~�� ��L�}-�SA�(�2�	u�z��`Eu��>/��sf&���%=���ae8%����@&)ԙ��@s��Z/�{陂�n����pw�y�P��$3�1��5�S�)�{q.g^M&|���s���t�S�D��B/�pC[k-u�������6�]m]�jE�k76����Olk4.����i;A9Z_]Q6~��[�j�z�=]n�Zoe�iw��+[[������\�����+?z�O�O^|�dG��>u�v��@���3B)�����G��E��a��ɢ����4��(�0e��&gz����=�Z���՞�[�����ֶ������O��G4���lYf~:X�ӑ�zx�ӳ�4��<7�(�����0�_�����`6���3�ċ�1���N*Q����EݻwO~���S�x��/�zM������?Ѳt]��5=����`���%U�U-�1������o�*�e3����N��e�}�����W�d�g�`E�X �!��S���ru��(	�����7�jkk�ڳبq=�	>v��2k�~��j��ȖN�
6�����Q�$s;�CT�����D�m�/�_    IDAT)NK�_�`y�S�g��D�c��-�	_�~X��fӃ�TI��z��Bp���=��	�bD���d��#a2��i1���M�dF�~i��H���D�YoW2��r��Q�0���8=�X��쾓M�1�szt����,ˍ�ބP�"��ɝ#���w�Jy�Q�н�juf7��b��E�e]�믿n� ���<g:]�ּ_��Y1X��4�+z���o��Vc��O~�/�rI����w�jv��R��>�����V�]����ѓ���ϬjU+�T]Ԫ�M>ϰv,jm���u��j��-�9��M��u}�G��?�hQjjV����(]͆��L�?G�+�Z��U��Z���R&@�g��*_B1-�;��1;=�L	��G��^��s���f�s��T��f�<!)N R�6��ٴ�חU��(d8؞�	�r�O�g��?{�i���D���������+pdK�j��f���n=�KT����P���N���^�T�Z��G�=8W�
g�n��J�:�j0�G�A��8�2�UW�QR�����n�o������_���l���ƽ���ѽ'��~���t��ϴv���^ߦ�3w��]���LJA�/.�O��FZ��6Wѳ#���"���T��mݼ��Ŭ�ʈ 6r6zF��5�R-�spa�D��SF-(���4����P��WԮ8���&����d�ui�����o�r��XP���A���Z�pнu�'���'�v���߸���꽟}��|K��[���51Y�e8o>sU�����^z�:Ҩp� E������Z.k�9�>x���➒ 9S�T�����b��r��[�b��&���D�z���5��WR���E��Y��\!`����e������r��-����U"?g���=���oz�O{�d��*?�a��:x Ӧ@约f=A�������V�|f	��^H� g��U"� ��>}�R��c2��瑐he��W&6�γ���8����d(=JǞJ�$�;�	,Ge�����SL�#�E�6�C�cW2�
�����f�cMGG*��j� baW���FK/���ʵ��$>���ۦ���v:;g��R�\j,��ٹ�ܺ��^Y�G���ׯ�=<���������'�$�� ~��Y�����~�}}��FT���g;�	��^]�^Y�f\3c��f�5;m���U}�ǟj0nh`lM�FS��T��]�F����v�� ,xJ���3gbg�Hu�	G�g^�9J��E��ύ�2�v���b=%���re�4���g)W<W�#=��D�o$�Y&ДǯԪ��>c�W��v&b+�V���0'���e�d􆳓�!(�So o+�
���@>��ֶ��k��JQ��tS��CsmŶ��"��s���%�j��Am9��6�4j�������{�k����'��>�������?��ɹ�+����c�
wd�����������6�u�����LY���^�/)��Z�mH���d��p����g�6L���%���uX�ѧ��X&"N/�g�@�yoN�b��'�^�ge�c��k�4>��� f���®�h���F���\ԛ5w����zI_y�g����~�j��J�MF�Mjŀ;rq��E��o�=H~tr�
(�C��HC�W}���ٺ�M�X6X�B����f����e3���s�b�*|`��;
Ÿ99%oǠ~hU;0Y� �p?2���$`9s��C� �!��]	"��3)R��	j��0	XF������ox�1�
^�g ���`$A9;>��2�v�dtb���`���	#A������O"�T��4��J�I;��y���.k:�.��NV3����fT'��4�he�F=�=��̽���3s�<�c�|8�`�h1=W�)u�%���tr�n^2Ɉ1;��Vt�6�`���n811`>�	�@sH��a���s]����^E��w��_z�,��:�o�T��ݏ?��u�^{��豷����������Ç>�V��R�奺+L�\-ը�-ratաƊ��>���OO5�b(RW��ִXհT�����yI������j�P�Z��#�-����������cm�B�HUb�Hi��ƺ6g!�Ӌ��w���<��q�ԯM����m6�P���3�BN�B}�����BJo摌Є�<����LF�N�h��6F"�eNB��Y���s<Z<8j屸���p����h�,�vc[mVum���l������?��MkM+m���ԫV�R(���H%.T��j�7�q������_�`���w�[?����w���ǟj���=�%�I5L���l9��� r����dFV5"��q�,ؾ��ؠ��ek(��z��<Rc�-�Z�=A2.�l���o���꭮
��A]�����l�a�u�yz���,PK�R1A9�����Bzo*2|�����pg���kβ�9 v�o�?��jA���W5��o_��*7ֵ}x���Т��U9D��,�Y��ny�~8�j��@�څ0��%l� ���{�ϋ���\vM��ֶܳ��E2 
��jO��aR�R��\S&��3J�f�GJ\-�i:�2b�}����r
k"�fmV6g�L 's�<p2l"'^����B�B
B��)�s���Yq��\�lG1Ve�fmGs���O~��F@�Y"؁��dy�\��E�6&��H<L~1���|�<�D��z��jUQ�J���a.�Q�J�$�$��;0�kJ�0�p ,�!�a�ld\�>���~}u��u3?0t{�JO+�������^�����sp�N��_>W��`���3���C�>�ǭ���i.������[wti��'O�Ui��RmK�=|h.�k/�ѯ���t��5W�������7OG{Mдog���Іh�j6�KBΘjkU瓢>�lO;�@��g���|�F�V67u���߿���Jg��<�}��W0y�1�:A�1��_�o&��\�:��i�P�OeW��,^H��M(�	a������I^Hj�5�%��5-����3̜�Y;�%��&g��5qb���kO�:+Xe7�����&
&�4JDی}�|��0Y��8K�0���b2�a�f���zS�7���kw�� ��۟jT��k��˕JE됣�e5�UUͱ�t�]��ֵk��l>�Kl��e���������?�T{��8�U��9؃8��҂j#t���F�H�qH�[CH�E������;��,�S`��GσyZ6=g��ں�nm�ǐʊJ�pxx�jr��HG��L5�x~�P��Poc���6KF�t���E��bR�s�ų�Ţ+�F��K�[���l��p�>.�Vx�{ݶ3^FF�˅\s�z�L����H���;j��ѽ�����Ț+��M�����-t\�aTe�J�/�J'Ñ��9���I���K�i�=�R6rO*��c��rlTw4p��|�%�M(�#=sH����P���d�y�$�(6w�D����qh�^��[����b�U~}Ɗ��B󱀒����3G�@��+`d����ZU�Q��9x<T����@�|]���̑��<UFfC�5��ه0��{��C4 �<S@,�q��:ۜ�e-l��s��b�t��mg,���g��;݁t�؜�9�<S�{��V�����Hv�5C�;;O-�ꫯz�D��&��~#�-���9�]'��M�R�j�U��+�ըNl�~뎃���@���j����z��W�9��������;����O�C� Z�V��L�U1��E0S���O���������ǻ:��U���?��WR���~��v�����`���n��ӎ�*�J'=�>.�@C+�� �5/!��ݟM�vџ!�"��N^�zp-x3�ٸ� g��3�8�b����6�#�:`-g「bY2D/��� l�$!!��@n3����Yk��#M78�sO�/]v���s�� �r�����\@m* �͕]Z�h�Y�W�|G/�xK����'Rsê_L���jZ�p���y�EԼs�k�����/����@��.0������������w���`�3��J�L�s�@h̭!3��9S�"�ȼƪթ�g�׮;c��ӏ��艡�+�/��iyޕ,�﮴]]z<��憾����O�l�0t�����q��#=|�H��{���;:8>q�1!D!J5��� �{��<=>�X��5݆	'O�QX�\�E��J����g����l���f�����q豠W[,�Uց���������}[��j�����c������n����q٠GX�<�Z�"f�y�	O����Gi{{;���Atb�s�C�ֺV�*W�UA�Xb���k7���K!�?��6���B��g m#��#��o*[*��Fr�B�X�ͦ`'���{�
=fGC��I��dT�>{�;�8EbOb�� ����	��/�D������x�1k��d�ʨ��Y߬Z\u�S-��촨�3ٶd�	X������G��k[������z�&�ʶ��z���`Kekq.��,R����x�8 �� d�{'Gjf#���G&*K-ɃN���[)��g�:ؾ��[4������D�7G�E2]n��׃������	�_{�
R���\_{���]^���B����VupxlR�+/�v�mTj&Yq����w�{���*,Fբ�����q?�jR�B��W�ù��'���юΆ����k��"��$���݋��m6Z~n�=����l ��K$M��A�K�o3Iv��>	�ϋG���a���D�2�T'Y����5���_ӮY	���:�O&4��Ԛ �®ϣq&h��������V��8=�j�F����s��qKː
;��9�\Y�~��U)͵������m������Zi�h��R�8�k/l�o�n���?֬�S���5��hh�^S�f]��UMSp����ݾv���Kl?��������~����}������\�J�C�E��y�@�����;��`G���)'á{f�k��-Uk�y�n^�n�/����+q ����?;�Q��Ʀ0���ik�X�d:�x޺��Gz�t[�~���:<8ָ�N��vwAx|D��z�D��l��e���	D�2�ѿjhmu52��B��3�G�;x �c���a��i@�����~���P�4�7����/��vK��wt|6���rٛ!�ׁ�!@r�ФZΛ� �f�����jgg�BJ�:�Ϥ�zq��Z*�*��Z �wUĘ�V����=�D�s�`T�vxˆ�]"����3�4�3�Q�3P�Y�A��Rٮ� ���$A�
?��^e�/�H^�5��VR�+[�E�D��pr�5�Um�3��ƨ��f잳�1"��)[�nX+6�y\#��et�\�᭟�ѬP �nH6�'�Ϗ"�/�3�!��l0�U����lT;|?A��J���9F�U�ɲ��1t���f�s�[$ACU+��C��s#2~x�����v�roo�{��h��!h�f�	�����6[�MGч�w4�����+o��WzM�Z_�`���ٹ�ĩl��o��I����b������?��@��T��-�-4����+�N�c]P��0G�X�����>�τDA�Ɔad�����*ԁ%A���ϜZ���,.l)�n6��Q�I/��g��('������%�o��v�7�ap6�b�,�;�?����a��g�nY�-� @�$Z)A�4�-�8z;�b��� ,�g�N'i^<��^�F��F����e@�f4���NQw�l��*�?���NH�q����Ӯ�Z��fY���7�������_q���k���nj���*-@8;i�x���_޼v�?�Kl���{��~�~����U��a��)d�bE�VK�"Vp���4�l[�=aJ ��dp���o��7�_ѝ�/hsk�� =>�G��yX�?�&.�%��^χ��0���B�Nc��-�]�p:���u����G(L���޶G �@�@�;��17@��?Oʇi��X�#fUɾVV����L��r23úU�F.�င�!
0��)�+G���|]ݖ��o~GK�ȫ7���T�C�*5�`˜*=[f9$�{L0����wo#Yzf���qc�#������v�d�#q�y,2d`��'�oҋ˰�7�!z�G�˚��1lk �c�Zg��M��ޫ�k�̬�3#3�}1���?+���9l`�$ͮ%3"���}�;�X�Sܹs�=�L��]�$iO��J!�ɶDH�Ϫ�Fc��_�x�B�IN���E$�qY�Z"���B�,��_�tk�iq`�9�h2�p�Y���qV�xjx})ӕX<yX���M�F�4ǃ����/gL|�%	���$��b�co@S�a��S�������0����?�>���Vb���E�|e��;���>3ٲ؊��x,�2����[58"�Y�=��sŖ��'���8��R	a����v�D5
���v��x�|Ld#"/b����ݯ~�~��r�hȏ{���SuO����<�Kg�8bnq��W/������]|�sX],`<1	���'��v�E��|��_GLF@w��w��G���oc�k"��9�8�k&�PV2�>��%��sgq<�:��N�~� �`�TA*[Ĕ� �-��P�b�L�S�'By��P6C��l���|�%s���^܎i.������S^-�G#�W7f2�?>�҆�����{�\2�eb���C�}�����Lg���
�Ki�3͚��<c�����l�\�ȫS���[��"zt��51W���0W�λo���=I�"�9������ �^�u��+��8���H�6���<�J>�j>�
�*�����"(&�ouy���R���N�n��ﯯ?���;�����sT�aw��8�n1L0�B�H0C�XQ�K��4�{���*���2i,���ƍx��,-.�桉X&|�f��ԝ7''W~ѷջ�xƭy�
h�)�~k�5�����?:��~w>����H)�KK�
���F��B�?,˃˞;y3��2�7.a�j��݊�f�3�'��h�h�රpn1�R�>����bh~ﵷP?������y���f��L?�/��/�M[���z#���C��{����O?=ỗo��m 8YF�Fh_Gmm� �X���w�
����w���ǘؑL�?&��z�g� �B���AF�u�.���@QN�f�A$��l�%֩���D�1W��b�����Xt��7(U��r�&���{hJ�/�GjmccdsI5�I�!���%�Tl�$BYԟ��l_,�:�a���z^;Q�Ѯ=����V!�
�0�"B���y�\.�w��!L�N���o[OֳI�>;�r�}�;�d�f�
u�2�0��&a=Y�R�nGH$��@Cyr�76�輾u�>k6��jY߃�%5zZ	�v����=��$O�����s�b�i�Q��[��B�a�^B�F�ݑ5��kW��[�����iZ�>�z�������`�)R16Q���6�L*Pr|�M0�g��O���E��,F��$F��<܉�Qm�>�a��y?X��k(=��_����h��,��y�P���^�����S�l`���
��	���a��4K2f&�{�<�Yt���Ş��3�-k����՗� ��ĂkB�=��pr5��)���>�G�_9ƽ']�V�&�(��؈V-%͚t��恗_8/?��u�{���?~��@��\��� 7/f���\�Bi��m�X�*�m&�@�+J�Jγ^{�t�o-ͯ���T�v��k������jʵ�>��� ����x3���2�����Vl2�D�0�^״��8�U��+_�������FR�&f0�M�,�$	��[����?�]#���wǛ��闣�FS�Վp��=���{��㏤�]�pA�g�����6�ݾ�Ah� v�Ab�ȑ�HB>M+8�s��Φ���D�h�8�Ssz8��cC r��o.cn>�����fq���Q��?��*'��?F�N#��,���,��{2���8��Xk��)���8mBv@�    IDATu�6mA��H<%w/��sΉ����A��SV(����x�Lg��!l; ����#��}?;�[|��n��+�-��i�R*N�&["+�Ŗ:S[����ܺrxP�������u�adL�(3"���5Zm�[�S[��пXf�?*aɅ
ж�̮N�'RªZ;�IGәM�l4�8�PM��B�����ܳ��C<�rNEm�~�����qm����v�JD�)��K�=4٠�s"�Ln�f}�iKK�&$ލ���%�Lz#e�Q�0/���V\&�1C�:����R9@D$�X�75�����u\�:��sU��S̢0�d����0��7��կ}�T
�v�Q��~�w�	v7�I𳥬e$�G>C���LXlU0{��G?�/�0���s�F#B�YMH�=������9��5щLd�C?�陚8-8�a:�9c~�P�su����}��D.�'WԽ5'�;'� #@ܿf)Ex*�lv��P!wM?{~jhũp�"G|]��55��S�d���>����S�G�gn���ͤvl�jC��C�У�M3��P�:f����:x��"���x�=����M����q��^}y��t�X{{ml�0��g2��Ȗ��X�_A.g��Q�$��������)�ۏ߹��sﻭ���hH�>��g��f�Ǣ�Q���� �n���Q�t�,�-�Y���.C"/ޥ���ƭ[x���HD#�t1�ߋ��͞nNv�d�����[�2�\���O��~�2�4d{�E��<��vw���o���W�F�P�?�Q�.Vs���^��Q����05*�|B�q��E�n��R.�ɖw��v���H�	���&^|~�|�>��ý(*�G��`��a�%��p6��h�@�2>>d|H�r&�M����Mv��͹�i�as����x�(bT,^V��EB5LssUI>h��]3��=�$֧|�Zei��:h���y�ӿ�I	���'.eqR��lMc;x/�P�:�EE�[dl�2t���l�<��O�$�K� 0u�	��:Vg2Ǩ�D��A�\՟ow;*�6���`�CG��yy�tF�t������w������6qr�=�����P;����?�I�������%l���gc [���OM�d����a�g�ƙP�ZX� ��=�Ѥ�l*@u>�A���Ο�j��b�@�D7�WVљ@���a����uj&)G4�I8:埝��뗐����;�ꭋ�x����.f�KMs8j�%3�z�"^y�e�/�w�OPo���~��C��L'��Y�QƙI{.O�S�-�?���;Op�	D��Y�f$��n� 5���?�rm�]9��)Q�Q�P
^o�Ü]���W��k�XZ���EW�k~��5��w`$��q�4�?�>1�?4���޼��Ĺ{Q�5"$#{&8����YS`@�8"��-/�r�^|�\˙��[6��o�l|Ϛ��&lO)�#$R�X���#i�HL�vpi%�o}����:ַ�����V�|+���*^���+k+")�oֱ�?Fw�D�XUhL>�B9�j6�9fy�:ǳ��߮�V��/M��������7f�b����E$A�]�����8i�qx��6��X
D�j���_����q��M\�x%&aP���y�*�ԠZO������P9cz�ҳ���S�'��^�2�$�3���#|��m|��׵��W�Hfs�����Im"		��#dBm��,.�;SJ�A�-(<K3���0�9$XHX"H�(I�ǭ�/�X���'��R�%���5�H%�Q���#W��v�t���Y�|(Xl�0j��	R"xy8�O���8����>�� �!&�ON�Q�A΅<���k��/�U����y�j/)	D`��@���^:BgG���HJ����eW��'�)R�$�[XCC�Kf��~4� �fS6�y��q�N)>̂��4=�CB��$��{�3'�����C�ny��S��։���ÔN;$�PZD����/B"�H�k�6�A�n7�M=���ߏ�&��وSF�0M��?�����΄�Yl��fQ!��e͇ľV<&�hp�0�wn.����K/.��`�!ݠ��fҸv�P�|�<�)���DFo���?������d4�g�kz���-�ȗ�W��E��>�Ѵ�ͽ=��+��+�����G�?��qm���5:���bQ>t#يm2��'�m,]����O��ُ����,�=�pLCc�[A�f��/*��gv�܅�b�D�gb|�_Eۡig'[��G��d&�m�f@�~p��﫥	�"a�"~��3��ޓ<|��&&j\E"t����"W�z�5�l�h�-K":�F���5�41�/�ۭ`��6kQ�[L;@�|
��	rHRg;��K�|1��j�Dz���#<���D�
�(�.� �c}����!:��BE��t"*{�y ���e=��b���˿�KQl��_~���7NN�̅���!�AA���)���$1�0|<�f{�N/��$���6z�8����0_|��z�E\8wE
�u���yF����&���O�g>VM�Z��2A���ff��r�k2��/�@����z�G�������6�_�,���4����D�DOI<p�W���lJ�|dVw�-��h�d`�\A.�2֣X�}�&���W/"M�����үu��-2�c���4��l:Ԍ�{a��n7Cr�=b6��w2����
��~N$&�9]���_`N�	����}Vl9ٲ�r/|��E���X����E�9F��mZ�r���!��ʩ�חȆ�)�gd����MG��&���u���f��s�Ҋ�D�M��\����U<Lx����ke��vO2���P�rҝJ�����s(0����$HO�C��a�����e���(�zI6XN�-�+7�Z�3��~'�nͱ����b�u�&R�Fc!Ҕ�@�A#�g������Cy=��MS5�a
*W{�¾��p�g��X�½޾L-�\YƓ�w,@`2B>��s��Ԏ�&z�0pN����f����χ�݉�2����o\��d8���q��V��B�Xl��"�k5��������Ulo�Z�:vw�����R��&'H����� F�N�un�aWۓ���D��3��(�1y%�ОE��k�q��ۛ�Mn�#!�<���:p�t��W5��H��ܝ�F�TC�/���s C:i�-�55F��uM�qc��{) ��	X��KR��rj�_�o&xVX�M'6+�|>�<��1��3�2_l��Rs�J�ؚkZ��D��	zT�j��F��)L;d� W�W��1?���"�Ӯ�!�\uZuĢS��U��<xr�͝Fщ�HR$b�,�+��.WLZ(~�\^�O~)��ƃ�����{���E�!b<�E���]�+CM(�h�8;f�x�7��`�x��2�]���n����RI��Y�l�)R��#O�:�}��/��)��z��Zl5��p�3�D?��g�.�tfND��~|�^�-l(
����۷���$ߡ?gtf�� #N]�@{N2��'H�����.V�	C�����l�x��W�q��O6vTl��Z���ӳ��N=�����[���u����9R�D_d�#�T'U��#�T>�u�yD�,�8�T2���
�s
! 	³3���d8�A�wx��LtVj{t���hW�?�����	�ʁ�5Vv3Ā��@S.;·<D���Q�O{t��u1(L���~�~Wqvl��h1�.e���ɿtp�h��@���)�8���-ͦ�!�4<	��'��BD�=�}$��P:ȑϚ�X��ۤ#���{��,/���AƱ��Qy
�t�)��~'O��X02�W����8�$ad5 � "���<A�G����x������l���%5і��nT|�-ڒ���hH�y7��Sݛ,��P;������&�����#W��F�#T�6}/=��B��}�1���n>��{��oՐ��%��*%�O�#��S	2�$HKp��;�iK`dUl'���>7}ήaeQ$t�{���ͬY�xh�B؜�_�L�Cs��H��N���f��X�D��"˜d!ک��YX��N#��qOD��WH�I���
��3��O�QBVT����<v0��~E�r�6>C~�&	�_d�kW��I��e�����f��i�#>Ic��!�R-`::D!,�%�JG0W-I�����Rl��y��Q<zr���1b�,���և�Q�l�\K�
�,����KK��D���K��RM-��GW?��������xl���Xg��$\���D�T>R�G�9�&�|��?�ƥ+_�Wo}7o<��jEnH�By6�zF��3�i?������'��9�q~_龡A͟����������������vK� ���Ǔ�mtt�}��G'1�fPv�h"KFN,��A�t�def�rS��n�b�F�=��)�������ۋ �Y�7r��Ef��L�'>�>�h	�
�%���Qߢ����AJ�������t�L '�u|�S�Uxiޞ����� z3Pjc�G#��H���z}�jYly��y�NSIt4�q�Pf��q;=v�� ��Y\G𠑀|�5)����v���B87�2�C��J��$^�φЦJk�X��~(E��Lg���Ղ$�Y���=�H�d��rK%��H�li�����z,G��9��ݱ�h�����`�����d�u�6��<8%��qgn���hC���&!CΖ���ؒ]�YVlS�������1r� �R��-��^x�">��>���R��?��t�|~��!~^JRv�uM}�xD�ݛ���|�����X\Lbq��1D��P�\A�Ւ=�/�[�������ױ�~��E<�Gt�A">A4�f$�L:�b��3�'�b�H�_�ࣻ�h(�K������y������׉�'[z��m?������a�n^�F��q�Z���p;\Y���~u>�>��:��Va�%�U5o�h���c8Tq��6}����5� c��+'w>��(��z�z�K����u���?�3SN�����gw���~_�s�߳O��`rZl�4�/�}�r)�r1���^n˭���<���Y�����O�٦�BG$�L6�\)'�C�=D	d�E�Y,�Q���j�r�+���ΗXg��2��'��w��w��s
��r�H4`q�����W�]ìC���mC��+��e���+(�K��"j����t��&[s�_����3���)�-�g���t�������s���;��8�`���~��&�c���V�B$^0#�H=�� �Ha�P@1�,&YP"�騅^g��+/�ZM���?A��F����f��6�,���ȵ��=tk��6�;a�ّ�6��07�	C*����h����^?uNs)Dc����<ɜ�k�ŕE�9��mk^\S���m��d7�If�`�P��$���6�Y�9��e�o2+��"(ա�D��ܑ�2;�Tb���13�Vd�
Χ���a��� ZN����I�� ����ͺ��,M;RhS���]&��M��C��<�e�%��"�-�����dИ�f�r5�����̦�wB����<q��f����԰�ز������9�1RR��к�n�g��2D��!R��Mۨ�8=MQ;^G�⅛k��ѻh5��d{��%[�N�6��|��"ｃ#[��0�ɂ&���T^[;�0N/�-�χXẒٚ`8;���54�}�>��5��0�q|���'�bg{�L��H'�H��'�I�8��1">�l3E�����-��1��	 ��pb00Ȋ�?x�iM��{w���&��\�?�5QZ�J��u��'ľ��B�د5��up,�����N)SKXSF�"w��``���*�����WX���O���"�<���hg�&n���AG��\ۘ�����Y���/�g�'!U:�Ҙ���)��D/)�T��	Ʀ�ܔ
�\�s<�	�F���uM ���^7�3��,.T�0���Ҩ34�{�;.̗17_� 3Y�.|=�)��e��/����^|�蓷N�7�"�
r�]�=�����b��W��tJ���Q��H���__y�K�:lH"�����e�p���v�E���U�C�u��/?�:2nw�)�X�\��>�٢�91�`8�ko����>:�����-B+Sۡqҥ�n�T,�h{��3�[XB�P՞�_��a��Z��R���6��9���h�٣F�8��6z�˜M�)�=l�`>�0�@r�`����Cko��������-Y�����hg0���b�*���
*�¤��)4M�ڿ�qi86�)u�� v��f@���MQ�ͻز�-�͓S�`z=��d�hS� /�7Y�⾘Ŗ�$I�.�C#�p�H�dM�
*�Y����L�^�����L�h��m̝��R$�p�JR(9B)t�`q�#��C�v��v�qJ%�95;H��*OlG�& g��sN�(����Zy��}ĝ;=��p'\�AJ�4���#�5�p<2F>$��K�D�.�O6��6��WV���o���HE��Sf1�`n�������[�_��6j'�1����R������cmy1�BN�4��U���o�ީ [����&��I�nWV�t�-<}� �V���HG�6��N�-�'�d�t��>>���f/���q�َ�1��B�C�50�V�L��k�T�u��B�`"Nf��E������.$#dl����Y�؈�i�DPc���p�d>0�=�Y6�DC"����;���Q+�3�]�2�p��L���:4���I��pCn���|vB��.��83l�`0��X���7�T�Y��8��}���{��7�/���;�KƑ�E��������&"2�A,�v��Vӂ9ίTq���v��6�L�)5�<�h��P�bya�,����R7�<�K�l�w��/���b��h�5�!u�3��C��-�����.E�%�����7��W^�����F#qX�;�$�s��Y.�����[Grr��[�״��s��t���䅬m�ܪ���p��C<y��Ǜ��m�� ;���'��0Y�r�T�|e'�:u��\�T0��${�a�Ά�t.^�����!�e*�sܴ�of���أ#�d>@�l��h(�R.�$#�Y���	�{��}���'a~�F�R��%�a�'�"�XV�ș|�J	��z�(g \l�B6U��S�g�2�!�KY�q��8q8�c�1F�,ʧLa�Or�����96��$d�l>֭CIP�l�$��tH0iJ�Ȭ|SK�b���!a�)^7Ncb"3/3m�Al�q��q�����%$�HJ���~��F�DQ�fL,������H��a}?!��瞝�9s۲�zF����f����H�2�M�3M��+N""I�O3�*ϋ0S~616�	��VW���h�����q��
�~�5l�?F1���v����dV0C��D�^�A�m���^7Y��dK�`�D�ay)�R!T�Q��xf���Z�dA��4���q�����S5��k_�m<W�w��L��ҙ�K�pp������Ic0K��-��ͤ�O���t���\,	��3�A`͌��3ř�J>lpEpJ�����x���]��2y}�I�W��1��/�R,��������C�k6�>�Y�Ξ�E[�m7}�V��L93� rE6�SY1�)��״�PN�{���x���5��&�M"N|/�o�|��$�����%���m)���'����9|[��M�d-�t��Wqum��>Z'5L�1������P�Q�!���\e	�KK�W�ߎD�I��Ҿ��b;����^{�����N�ݦ���>�������@�<0��tZ]��\�_��~�/^r�Y�s��<��E>%��{A����U�N�j;3�^}w�w%[�!_雹�p<���>^{�ث�vr�Π�V��v�Q���zKH�?A�PE6W�d��&��R���|�A�N�e��n����n�����:��Ջ�O��9�a%�q�D�[opBO�tR�<p��9�}�
�e� &y��S���Ӝ]!}�%��Eo�"b�
�D�t�=�ܛX��:�����^�K{    IDATHL�!/�����GDZRj�H��9��,�m�"홙F�28���Թ˟�DWl�i:��A_ƪ4M.u�lH3��:b���ힰ铇r:e!�L�������t�=s&�r�>SVz���w��"C3�pӏ��'�|��X���e�'b�M�Z	��;[<1��L�U�]�`��v{��5M�V��ۼ�ݾ1�e�Hϩ�p�^����!�h0F29E�Ȣ�&'�ry�|Z0��.M.�*�4��u�S�p����y&�Q����0���k3��T�8����`<8�{X;_���v;GiT����IEFr
�''ZO����u'�S$cD@�(�Rʯ�Ԯ2��{GJ�bH���o�G�9N)�g#��@�d�S�2C�xh�OC~���c�"t�Ƞ��/c�4�ϖ�y�5�'���̈=�N���U��5���&2$��!d����8O��n�}��0���2BikF�Ԫ( ߠo��l��.n�d��B�-�K��o�ݴ-X�&!����7�H�K �(�A��D�K#� �9��ΐ�A�+�X���X��r�l̕3�/e��s�06����
�YX:/���0"w�L*�s媸0+K����}��Ԑ/�g��b[ۺ�����k�u�����C�b�Ѩ���{������5���x��W��o}[�I��l�V�}y����E�>_l�Vp�������
"qNR?�g�!D���?z�ܿ�V��I�P^�{�t
O7w����1����|^0���!R�$��U\��"�0e!�u�������%���`�K#]XFw�A��H2�n5��
s��)?��<�_%�s	�X4(?Kv�5n<zl�w���i����(�2K�ED��/ ˜�=b��8��6���R���1؝�5������]>ITc�u�1�i`oNH��C5��u�
fW.����jcʞ���!f&!\�<F����O!]A�q��H�J�L �t���&OB��s����zYh�E�\���"fw�Y�g	%&���=��=Y�i��MX}�?�l�l�o�-^�i591�~�9Hy���)MHZ!���E�g�6���d>��A�X\J!�w���P.��j8<�C��p��VW�����0R*l]���dE�YG�}b��}#�̢$��u���e�&���)n\[B1b������9l��sH���v��N���	B�C2S����Ɛ��E�bC.�G"ERY�X&�����`�nA���,�����\�h���ؒ%��͌`c����c1�	_;ƻ/���� �KY��g�@g��:�$�2+K��Ŗ��;Q?m�%rş����"lF9��H;��.�Qz}.
�[i�o�~?^/#�{P�����f���+�>J����E�1�5���b@[���>�(Ⓢ4�����������'Rp7�j5��(�(f�q�*�����kwp��e��"v�"�B�T�J1����ŕ�_����/ZG�ȟ�R���o�������u�v���u���#4�S�jV�+a~�"�(!���w���e��_�<w��C>���+6k�_D��w;K����|�P��9�f?�	�yꌶW/�`���>�w^�.�����ci�ӷ���B���>��O�=F{0Eo,��!�/���H�{˥2n�?�`�C@Ӂi��>�^]ƍ+�x�Ul��9tF1�Z�t��g����d+�|p9�r�᎘�"�'��B_�w�c��(v��:�%Y��Ԡ2f�jk��bU��Z�O�/^�t��a>0�wJ"!F^�b0�p�� ��c^u��|M5b����۔'�:jr]��T����n��Gh�]>��ͭ�lgMl:t���6TR��be�L�hE��N~F�Ÿs�-N�k����S�=&�}�6�kW숀�3���J+�6	��b{k+����v��D;�8�V��K3�E�����dK��>�����8M�N+@������rF�6��![�Q,dQoc4����.]^C����q���
�hQ�%��C����ў���k�g<ʵ�P��4�W���]|�7��;{-l�fW���+�v�Z�w������@ؐec2N#���-l<�"�!�<�d�P�����Үqc��b���Tџ �*4�a|�+����<��"$q�=;����m��n��=���1�g͔��.v�7��=O��!�����ʸ�VM��:gs�����[?-��C��Ho<Wup�1��j�s�y�$.��s3CC�t���<����ͅ����l+�z�b��g��0'w��^1�N���#2S8�	wǌf�O������ϑ薊!W�X[�ô����S,-�C����{N,�/a>��:�������/�g�Ŷ�9\���ۇG[壓<����Q�^���ܳ.V��+T��J&]��IG-���-|�֫��. ���N�,��ߤ	0>W�~�O�O����`�!���ԍ��>��ϊ�Ʈ=�"ǚ��������#|t�Ct�}EV���_�K�;:��_��3H�
��-�yR����9�|�*b�>�̪6����޼�����F��̼&[[rKy6j�&�l�`��K<�l"c�����UWp��=ܿ{�R��>�7��z8�k�E-�'ZF�,�a�|N�-�TB�!5�$?��czb���{��"�4��[q!c�?���:r������|Xw8i%��pph�Kyӭ���z܎����6�^���?�0�n�_�}�r�����0Ⱥ�b���<����it�=c�
zV����YD	��`�u��No)�g�i;Έd|3�(�	�����f�Ab�ɜؒ�d���~y8{����>��W��f�@TA��d�2S�Qʞh4������F2�������6.^<�ã}L�,/����K�Ŷ�-��~�8Q�Ȥ���׏��k�b���}-Ic��Q?�D"���^�!�������Q�����=��r�lO����&�SF�@R<��L�hK���l�L�[:��^;��b&����{?U��U�S��3`1�:�A��<ـqZR�s����mP
�g,j$'���Ӛ>+�~e��"�?���J��v�d�ۿ9٪K^g%NR�q�`zd"H�ٖ�IIƄ8n����%=0f���#7�E�7�wB�jn]�(�)�2��*�d�LqG��ٹ��YU>�!�Y`*�>B��Xl�1mz���'�t���陙�.i��<��c��'X](am��b:��ځ�m�����z��̞�X���-�������%���_x���6�ڇ�o�v7��w��qC��J���0W�J0�P*�%!U;�,`{��d��֯ai�R�����p�?����k���v�È��3]�4��j?�#�M[3�8�����+��G�M������������4���߻~�9������m"W�W%�	#2����I�ֵ+H$��?A���7�ṫ�x�ͷ1꧐�.�=��N?fK�!�dȈ�I�l�X<�J٢�"k<P����C<�{�l�|�&�K�!��w7��mP���6�B.�U��S#W*��RN��EA�C1�Y0mj�0wk�h���A"�p���r�Qg*����˦14�vx�J��z&��Ro��A��yd.�{i�u�*�����`06[ʖu�lm��ih�����3ja��gl>	��n���H4LW��W��,ac�Z	S���K���PD(�2xM��u�'�������lZDH�!�-H��ab'tA�d��u��D1�3#��GX�O ��y����M�"#,/�c{�)�X֖p��%t�m��m�U���a�"�f�~�`�w�g���T֎q\�|��u��|nY2�۟n`c;D�z�׷U ��%��lm�v��ᨥ(�x���!�L�I���Fiilmg�b�ͅ*�L����Z��A^�v���o0�~�O������M�H ���f�b���,;y�xL*f��/�g��02��?�Td�K):�v0�K�M ����G|ʃ(C�u'���9�>N�]o6aܟ���F��L�H��w�ȧ�[H�1���?ϒ�,�B秇�]���C0=���	��g��f4t���?b�q��� A�tI��'�'�XJ��|s�,�1���8>i�3aqa���_&�C�:���+������~����Ï���;����Si�(���͆�ᚯ����E�6fS��#J�2��o�����֭o�����ek�����������A�M}���7�ى��,?iYݷ�E����|Zl	�p5U v��;��ƽ����Qk����
fMgڕ�i�HQ}2�]	��q�`�/_D��<��'hu�p��y<mEŶ�K LΡ5�����\e�)�9a2��a�G	{���áb{�>������c��wc¼F	Lg)�2"r���u��
T+�x��mq�����Р�z\�� �Mh��e��3Ss��{�������_�a9�s��Μ��;~�Vӌ<R|>'� d�������vQ�}��!���PQR��k�)8~0��|�5�r�}Vgɽ'���S�t� �ײs�2(�l��ب(RbH��̘�~�a#�UBҭV[�V�n ��ܞ���&#�[-��Y�-���lĦu�V��l��H��x�t
���|�`�St��XX(JN���!ҙ�]_����N��B�$o�I̤{$�����~0$�7�H�V�1�[M��/��9@>���+�����v�r��W�ѧ����P*
윜ึ�	-�&y '�	�q�j
�����t�#Q��!r�"�$6wZ���]�zy�����f�9V�c,*>f��}�{�߯����d�k�w�n?��b���+�=�7�g��,ɏ1�y]M;m�u�c@Ձ���b�����	�M�k݋Ϊ���e�IR���{N�m�*a���ZxH���3�)3�ǥ�l�:�h'Rb�`�(��<�6�]Ģ3ՎB&���#�[-�霔�9��Z�aׁߓ��t<�r6�J9���B�$s���1]ʦb�/-��3�D^,��rq��ykʟ��~��v6�ſ���������֡겒�Lp�<m�z(d��"�L�tL�ݡ�;�o}�o`i�qo�o�և-�b;s�w?�;��V��g:Cq�a=���Fw7��@6՞��q��u����?��?��x���N}b���H��Nh�0�����`��Ƥ�µ�X,0m��k��j����x�<�����v9�Tl4��6�~g��o�Ⱦ��I�)�2X�X@5Er�8��n<Yǀӓb��m)���9�q"J��r�ep<�m�\B�)sy�T#�@��"-��bˊbݰI>X����>�*N"c|���~��*�JёSؙ� �n<����c�%�Չ��2�bks���d.��];��<X<T�Ʉ�e�ג�J���(�:FF�:M����4��[�!j�;��5R=��m�e��u&R�)�i*�4ݷg&v��������i-��B�'k��!k�Gt�2;A�K�Kٙ���T�!��F��٤����������B
��vdq��E\X#Ԍ���g@�Mj59ݴ����M��%I���k����F�p�ZYٹ��b�(�0s�߾�f��j���$�V��ųE�!2��� �}�'��Q�%�ϥeI�R."�H��扛l�D��0!��;r^�'��Ą��Mr��V���-G�
$���,7}A��+��=���D=�Y6|��,������h�;���4�?Wߘ�u��Xl��p�B5?á�	~�LD���|}|���H�;cUI���B��:��U�L�&@���숯�ރ���ǚn'���k�qnu	[O7������6l����T
� !�|&C6�J��R�%��e�:�ޖ��Y�U�ۦ���dro�.^��U4���9K�O�q��V�_������vwOd(O�Tj��ky\X�`��Ÿw�|J�w��$j�@,�ï��o�tfeqG��ǋ-����w��b�JR�}�կ�q�������L��ق{�3�c`%�D����/������`b�,�~�L^R�F��0�G�T��f���z]u��.����f�z�c�6p��^z~�|�	�}N�Y�'t�1�"N�,�d#��AOtj�V-3C��d#D��qj2�㇏����~��b��0=�U!�.�89�i$�0�F�\D�\@����M@�eJW�/��d;��n�����7v7H�����i�sd���roG��m�l2�(��p{��fl�������,�3i��e� �i��K�M?Y��bgs��1apN�c���s��?��9�N�l"E0S�f0��V���f��y��IC���_ȓ�;��s���;��ڵ*4 nF�|�<L����c#��u��������-�2�d�
�ϐhA�nN�F�'�N�r�47E�,��}������|�.]��"��8쎔��B��bE.B�?4�Z`��1�2lS23��ڥ+(��kky,-g�ֻw�d+D�tY�m��THx6�s�@���0N-/���b�Ꮰ�O(+;�RJ�T�"��I�\\)�ؽ�!��@�$�b_�v"�����bK�(N�BV\���5�I�0�#������/�~��I++_�<����)l�--
��`^���,�2>�V`���X��:��)kb홙�]�����˸Npϖ&K�C����Y��V,?{fHJ�}��
��+'l��!$i6���Ջ�y�V|x��6��@v�#��tb	DcIi�s��X��<W Ӕ�<��h��3�%��rN��d2u�X]����?g����v��q�����ѽ���<L���L�p��"�H<9F0�c�k���H�)�ތ"�?�[_��b%6�`�AR�����@�r��������ݝTu�.���z�nP��E�������s�S:㦛��������~�z�z���I,,��~�t]j�EDC������ʸ]*�p��*b�&�6�O6�����'ҺV��posǭ���8�pz�	wl$%3�z�y˺�d�v�����l�nlbs}�`dA�6��ɖ76#i��J.b!1$�l��l��yB02Fv�|�:]z�����%j�ulZF�
N:ER<�D��;s 9�9V��7����M!���X8֤4��4�'=N�"s�Α�w���q� ��ϒ��	A`"����"��Np��̇U�mͅ�E(Y��=ML�NS���*V�c�g�EU��C�5~��hpB�������f���b�W|��-�Shp�"y?�P�ul����0�G�<$�i����c��B���7'�I������� �/,���sΛ9�v�'��a}N���n���:�5ԋ�7�L�I2�W��"=��J�)���#<X҅˸}�t��*������`�h@����(f��|�뛠�Q.g�	ӈp痍"U(Kg��G�?
1B� 9�GZ2��(��z���`R��[��Dۭ;�L�����R���	ғ�<��� �<Ȥ%f:eޗ2����i,..�\�����!�=��������'�{��?۟B�\���D/��(�;6S��wk[~q��&�5���$�zO"ś޹�<F:P.�qnuQ�~~�p�{5ds}�a�#���~�$J�@&Lj�-eE!�r�U<�#H��J<KF���+�<㇗V׾��U>����O�[��b��w����|��b�R��Ͷn���4�*1���btx�(>��i�!��P�^�_�U�XiR:��v�z�����9߁/��>E��mY�I���y.E�[����]��g^���4Kl�)���G���}�=�p�k�{�Je������NF�#��Hg�hwprp��?�2��[A���1�-,/f�^��O>E-�\��G;5�Ȝpx �i�9���(�Ŋ��`�h����>��3�Alm>�'��십��)�g.�+����UǤne�-Q,�-���Ȯ�=�c��m�m(���#�C��Skj���������wa��4��/�>$@;�3"�^L�qLH��KسB	��0�0��/'Y�YԢ��
&���&�o1'V�"����MC��pz�9�;?;?]��Z�w.�Y�c���4��gw�u�nٔ��)�����3����$1nwl�9��R�    IDAT�@�c� I��u�� Ȣ�I�H�b����#2��
N#ar�J9�ag[����C��-��Ν_�Ҳ���&Byr��&[�'Gh4X��l��<�A�c����9�<�wP�XXL�O7�d'�X�n�H�w1��D�}|�᠍):c���a>F.E�"J�~���D4�f��LD�/$�-Wq��.~���,"a�X�H��@!q���Cݫ"�e�s��`42�<��~V�]�_x��!�?ˉϯR�}��{:�Ҹ@׏�)�%,�|l�y?����[Ζ�1��(�R:_���F�{�{Zck�~�n�D˝�����uϯ��eJ��'[~/"Dr�RN70t������@��v��TZ�w�>��>��sEE�r�2�İwX�����8�F4��+X\;�gR�ɴVHE�r�(�w?�b���������>���o������G�՘Y�S�)w1���b��)�<�G��ف�7v4�ci�&�]x 4@˿�tU��LFN�������?g�e����;?ә��&�?����� s�Q�}�֛x��7dj��{~��(�|��G���p�)z㩴���<�ɬ�ۻ�[(g�X��Q�M۠�fmKi|��U<�� �	��2�[h�0ۃ�����1��#S�w�$�	J6C|>���666��{�� �_4��n8Q��D�1����RΝ��\��u�3����I2�c������l���40�t89?سSV,~,.�F�NG�R��w	S{�(M��D�[M���Y�MǚV�����3�E�)C�$˽��4���~>?1OH�d��A-�,O���$FKg;�c3T�d>"��󛺿�]������n��_#�����4Ȟ��_d�+C~��g�Ό/2�^to�HsJ�KG�5����c����#�1�>���B.�L6Ĺ�e��W��ӹ�<���(��S�p���]�����7�,[�k9	19���y-��u,��P.x�d��y�b��p]�@Hm1��I�~�=���E�����H�@,6=�l�6`�m* �/`s����]G��G4Y�8��-�r��Ŗ������~����������[C�Xlcr�{�\���O�����[;ۘ5�,����Ѷ����@����,b����d���I�N�+'=�ŖϬ�~�#�7G`�{�hJ/�3����=AJ����y?�!�X>+�Sz �z�����5,��nw�l���L�A.P��T2�K��aq�����5||w�HR:��a�U�M%l��z�x,)��\6�b.�B��0����7��s��/|�}������`�o��٩�כ��I�3vE�^Y*��O"F0_-�\.��"�gq��(�W�N1���i1Ӛ���T�����(�v�?�����l'�g2��� ��ĩ}�G�$���7��y����RXM��|Il<����1�4���U�Q(Wu�qwʽm>��b!��b�~͓�U�x���x��&�4R����Nd`!Z�����a�Ύ-���N��v��?��;�a�Gعb�|J��)�Ñɀ��L-���]&��~6�	���R�
�gi�:�1	�B��^��!a�g��f�!v����Ӳ�A�E,p��ܠ9g����^.D�v��:��7�?2��|d��f���m�#��FoN�@vN��c����Ǆ�V>}�y��� tCy49+���~�k�/�I;l@��k��)���L$���.S�;��Ȯ���SB���ז�P:kɘ�bGk��S)�xx��'B�S��q/#WL�ҥ�[����;�0�G��E��X'��w͂r�Ҽ���}v#q\�x�F��^)"�ak��F�i�6��i�M,����79�!%�hf�6Jt��3�I,T
�ZDd� ���������d[F�Mk�����@��F9��e[���l��wk�Ŗ]���⡞E<���Yq�Uǳ�����H;F����CY���y�$dE��y*�lf���f���lG��C F��?�*�^��5ql�=Y�?Ӿq�����I����$q2&T ad�t��˫Y|����������z8<a��x����� �ڷ޻�1�He�jb�y01�ŖLzj�i�A|,��z���b6�b�)h	,�-�͕�����������ޠ��N�fWn:��Vk�䄶m�VR�ٕU+$�ƳR]�7^�KHg*��%�ԉ|�ت�����YkO��}�gE��$�g�R_��?S���	��~����x��7�t$�j��Lżn�N�QSc	OQ\�/�2����C<y�P1ys�<��eT���ho�T��k/]R��l�E���Z{�bKkHA�D���ȲX�t�� s9=$���ݎ(�~�ܹsO=R��Y���u �h<���H��0�Hc���X���veuA���F���T0ha"��� $���ir	o���!�Y����\v0� �.Ϧ3�#w)��VPy�y���󡧦�f<�����{���>�1&��ŕ��4K'��ə:�F�'�1IR�C6����ͳ%}��Zvؚ:	����b�����,΀+�N�X�Z����n5���� ��MQ����Yl-���61���+x��H��HHl������T�I��؜jYlYH���b�M�^]���!.4��F&�T���Ӹ|e�+��灞
�cj�>��ټ������W��O��kR�0í_�C���{x��ET*Q4�{�Es���޾
w��Ĩ���7����$�G<$HhR��"Ld	ȝm.G��35�QG�	~��}4�9 ^�~J6<�D�V'C>��ͫ���qєj*d�Ｋc��Z�����|V�<�c��5Y�����('��o�=K[��׷2~O�zC!RV<�yWl�$>c*�ͨ�3n� ��~w�z�;~�sN���;�H�˵%�I��N�>� ��yB�C ���Y��v���2^�u��Sý�:�jtG	}�|&�VJ��+�Q*��p}����b�լ�}�� J�(rY�1��5�3*d\_�<��4����Z[\��_������9�������pt��d���{��q���ఉz�#!��ɸL%����X^^����C,T�S��c�S��3��+nuQ�P^?�}���Vw6��~��I����ӿ�^�X�F3�΃����{���1j�mK�ʜZ= aR�w�r�*ҙ���w������v�tkK��e�k�P�m!����c��sȗ��D��m��&[���R��39d��r��>����ّ7����L G#�ۦ�a'�HR:�db�h�Xa2�\!��Ŋ�jgFL���p��d���1߻��Xl���ӏ�>*����}-)�V4찲��)9�M�����)E8bh<su��5�_O.�$�bK����b*��A�ݶX��8NZ]��8�o�d���nU���Hd�8k
�=O-X��Q�G���w�����hſ�v+�g��L)RĠ�aψ.|���?jJ-8��B�&��;V?�S��c�������(�O[�f�j�:���B�d��X����{趎���+++�2X][���׌��`�H\��F�Dg�I��P��M�4��Ԫ�L����1�5������ʸq���z����wC���0��w��A���= 6B�Tl��RQ¨Vl���L�bFSN�*��v������s�9�ĕ�D���b�(�Ԗ���=��;[��W�\��4�ld��~j�g�������y�T�"�d`��-B�k9^G�Raj5�Xc*�~�������ʘ�vh�u76�w݃�׽Ζ�)5®��Q����)_�^�+��Dv_|&�16=��5��p�C6�ƫ_Y����"ll��O��w2�4V ´��˙��7.������x������|i#w�//,��ϡɌ�Ns�yD�9���/�N�Ҳb��ϩ�/�OWΝ��~������/���~��{��?xe2nJ@_S>��� �'=eCt�;1�����7�7q��Y��S���4n;A=S�(~�k��O����	N&��������w��>�jl>v��]l5��v�?y�u�����8i�Б�(��F◈Bt{��d
e�>p?>��#�� 5��a<h㨶�B>�n��9<觐+.�3���LojN\,��^tC'��d�H�3�+u �iu;*
��''X__��b��-�Nc�Ftg�^J�$��<�ʵ-�X��T* _H#�5�pD�8���T�¨}���A;s�n�S�o��C|:�JI�i�L�u���ƂM)�WT����0����;XA���2iKy�z]�#��-��Vt|M#i�iy�h�{��VR1��r���t�[VN�hŖi'�0qw�v\cs�g�)]�m�G�'6.���l�qFv4�RNVl��&�l6��g�҄A���)��_�I�BvV���,'/:G"���9��N12=o��G�xG;Ѫ��r��-��J����������f�����N���#L���o����)��wo�&��_��q�{��by)�W���^w��Fh��=!"�t�ð�A�ݔ	���m(��L�"�L�)����4��l#�%g��G���x�N�$�@+��Dޔ"�H�d���?km��V�����4��u!�����Rg���P�'��?�x/s��$��;ڤ+ܞ����Xl��	�a��۩�ݎ�ʑ���Y��E�r0�4��ϟOg)��R"(��imYl=�2�ri�!��s�҄��G':��c��������+K�z�F�<z����}��V�h	��0��QH�s\9��B|rw=E"M����^�y+K��������Ve]�lv�NeQ��S�f1�dٕ�17ws3�=����ܷ����b�I6���$P�P҇����@��>�SЯ�}�CF�8ͨ�ӭ�=;�2�r��3c��}7_�s���&��"�ʁDfFF�[�����{�����Z����ų��ӯI���mq�+���o���_~ލ��}H��>Àr0C�;C�6@�C����|l�#�%�����~�wTӐ]�{j���˫2,�{��d��`�wQ�������f���$%��D-��i2��7�8j������W�&3礏�M��a*�t&P�������V�Xs��l��;�:��{��ӸzeO=F��B����,�F�'� B>d� EbI$T���[ُ�Ȍ����c{{[��>�z��n9��L�4���b#�'�A-��_���;m�D�����Ǡ�J�X�bܘ��Sq�::�\��1uB81�m��g�Y�����)2%���(Ş���9�fj
o2B!g��<xI�R��IѨ��Xe����D	����r.<�f�>IM1ݬhg:����sy�;�Ȅ���P?�c#~�C/�c�2g�y(J�6N��Y�&~�6�/R�o�'*�݆��[�sK��Qp?m?���Y�$�?�7aGA�Nq��{�����CU�/"Q+��a:õUG6MY�'h���1e����XZ]���*Μ;�{���A��Z͚�<&/GG���`>�9pB�\�YJ���KW�{]|~�X���w�{ln����b︅�=~��AcsJB���%(�Y�|H�y�s)�m˅<���LĹ�<�)�}�Ǎ,�̜F�w�J�F
ZD�
��L��_�{��78��Qc�Jp%������B�81}r# �}Iu(%3i��C�$�Ǎ�G�֖���Fmh�'�&*wa���hl
P|ޯ�T�x2^��C���P��\���Z4�(pI,Mxv��=d!��ul%�4���7W��
�GΧ�85����4�C�Zu<yQÇ7�PD�sr^��Ҩ��b0��3+XZ;��z���9�ꕗ����KgN���3x����ӛ�dzS;��_���S�bI�������/������7��8��ƾ���?��Q��0>�#q�[�}��]2����ץ"�T8�x!�}��c,�l�����@�
�!�΃��,�	1%��}�kL���b=yO�]�B�L�o1�'�f�����	[���Kޏg*%'�A��_~�	���?�}V�����'ì��+_�˕�$��ϟ<E��=�t�W��X*�ש��<F>\����[���BT�khvf�&��2���(E"(V�D�	!��w7;�=�Vvst��� uttd�,dS��J�}S�a1��0�d�_D��cqy+�VD~�����4Ly<&ӡ��&�}�=�
�����Kf�Svb��N�N��M�Y�pg��Z��0�M#�Iژf:\�cr��p+�j5��7���Bd�$��\���b)��:�}�$�Lԏ7�GK�$�AG�/�E��3�/T,`�-�!j���),a�e�t$3�V=����$Pp5��a޻lU�T������3���{��+�Z�@���3͠�#\c� x�D���6�i�u6�JW�R�S�Vqjc]ϹVob4 t��ς�Ҭ��3��3=V��b��c�<_���i���/���+Kx�����a�a��#��kf�=�i�Vu��8	�t�*�	�(�\D'�!
yZэ�˥�8_F����L*�C�5ç��5�a8�3��*'������Vq�[���$����x;�x=� �uƗ�ގ���$�[��}Ȝ@	�u&!|�	T�:�~&E�o��(�q2L�1�ڕ����{�0v0��:dB�R�WA2k��<'���D[t�$�e�M,����5�f$%���X� d����9�����{W��1'r�g����V�i	#/�v/F6㡐�QL��9����b����1<����YY���o���nyKF0��U,��i�|��a��(_T�e2]ɗ���KW��WP�-���w����>�<�/൑�cA%c��X��m�(K���g��t�I�����c���k�`m㼬���Nt��hċq�5��-�w܀H���4 ��)}my#��eMcgO��[���/�\�q;���V���37��̧��H�C:_,)h<{���#�'SD�/���bI3iq��(l�^��'[��o�q|<D�;����C��1P<D�@m�,����H�Y72$��9����
~9>>6-]�oɔ�D�I�+,H�ћ~�#�������{|�<�D�VLa�$(��F���T���>�^�|�*H��bIj�fKE���{��aEi�I�DB���d���1��lU�R"�a&dR�/{�|�i6�:�X�%c��8��j�lb�4�'61PD0J��<;�d�F��U���6�� -�oSql,H�U;��.�jT�%��eF`{��(ߣ;���D�LUjS��	���9K�����Uq3���L�,QK|�ɮ�~�XH��j�=y�׍14���>�Y~�D�	���V����t:�$��Q�!D�2���ٻ&$��	��T/Of�?��I�����p���yc	�N����{8����ϲO�1f0���Y�!�y,�B�ii!3�)�s4!�P-��F*
Kצ���4�F���͹�BL94�u���,2[���p��kh���rXK�ص���d4���HG����Bͮ����:X5k��#�{I
tg ���1�M����k�g2��%�},$���L2!���,�P{9�� ���B��s����QI�Ff��3��~�ͲZ�G�{],����w/`u�,��_}���Ec���`�4��i:����mbu}�>�����8�SKkx��&�^8�/n�����++X[�@!�x� Q�(62��R�ϯ�����`��Ώ��n���y��md�>�|���.+&�񈋋�a�,����$�^?�\~����b��!r���@2؝���t�7���Y?��4f�z��c��mquR�P�U��G�&z� e�k2 R����٧��Ge���H��/�>C��@H ���+X�T���h7�b�Z����d����+g�m���ѐ\X0�,u�3+�}'͞�GfYg�g�[BJ��Uf�a��6��b�+ ��!W����N��.%[V��|����T�:A� ,�$� i���]N��x��jc���R3�]M��os�X$�'��CK�5�F����nyOX�x�R�����.�Y��WSU,�o���u=S�%5z��$@�#�wK�׮t��X�p!����HV!d��F4aR�$D���Br&D�D��$�s��d"�ե#	    IDAT�2{���=1}wS�
�W�*g(�}+v��6{���"Y��΀���'`O�/7���-��tD�:>��\\^R"B�q
�æX��E��*{�L�Tq��	��}��\���ӧw���p�l^����.�=l`�1ad�uӧ�Ϥm�֟)�f��Ŋ��շ�(}�K�W)�$��7W�C����_m�э0�"L)�/$�W����=[�"���3.'����]��z����ƒ�t�[����LyC��H�3��SA�[P.���Ҏ�y�'��
��a�������<Z*�sZ���-5���Q��s��i�5�]B̽��
lm�=Z�{N_;��I�.�$�
�%���?��Y��V�#����n�Ⱅ��+�a���(�=D����:6�,�7�ν�x�h�6pisW.]�g7o�����"VVV����Z�)�El�,������������~���[�������F��������gP���R�2fʸY6�Md<Q�g��ӈ'9|��?A�z�ER�R_���*���6l��k���6!����%�753��h��n��|�_~�):��)ڃ���܈m����bd�$��('^����l�P�X�/c�T�O9�G&
��{�1��*�1����N��wDF"�&�X��G!�3�A�)1*��s`ܬ��n|���g�N>�%	}����O���|����d�t"���*�a�ʑRz�\�BA�����$JE#W��f6R��oi�f�����4l���f	m[_3I�l���~���y�
���~Tv�X��� {�6�:����[��8����n��l�T�2P$,nͩ������d�($)� �
��I� �I]�}�8��?ڲyh'��A��2ee�ǛlI#䘦T!5�CZ���@ո�;hy8��������4��`�)DϞ�ʺX_)������3U����������y�ӿ�ȗ��z�����6����g#�hx`��V5����o~��o�
��Z�v�vv��f�'��}�3�Ar̄r����ɗ�`;WM+�F��!�|�^\��z'DL�l���<�̛��fL�X1�2i�>�x�D,,iH��h$�dR�*IW_�Ɇ%>�7[��������8��$�2��|�g�BI+�Ml���b�2�cr���S�����)����_1��糿,���!'��u(���_A�B�DJlUa�@�o�*�h#�ʊR�|J����rz�������K�;|��[����C����ϋ<�V�l��r)�Ba��/�an�g_G�n|�X��o���g��ڍ;�;l��Z������768�G1_I�R(��W��Я�}�h��}��?j<�i6C�HRQ��N}��=�=9wi�J��JS�U��y�9,/_ťK?D6�(*e��ył',Ȳ?��4�u~hۈ��F�ӿQ�&��w
!��Hh�?�����|�����_�_���=l����L����M�#0�~-�F9�9��N�-�(o�E8����R��p��sl96��P<`�No$�3}s�4��*s(��(�"ɺ��Bכ��jP�Eu|y�KU�Χ]�6���&Ǚ��e&K���$ز�]Y[�
��L�\�Ԉ����L��VV����욌l�[�1��tlY1���p,�����)73�I�	l�J�Bf��50�P�G�7+�j"rBv2�����Lo���$�0��c/�
[��$%�@�w�>	�ڸ�~W� ǂ!���4Ǡ��C�Y�k�*�$�&о�[��2W����I~��I�Z�5�qV�fM��۩�CX�ql�g�d3P�~0ؒk���~����"ܠ��������>QV�@�SS�]ZYRCFr6��"C4�A,�@�����YO�yJht�Ź<�q��q��"^�D�m[���G��b{��8�!���M�8%�MR<ǪlǱ��J���$�(�sJR�T��g����l��l�L�&$A/�U�+���)cBcɴk�9g-A�J*����6��D�r=Q�K�?�E&b,ҿN1˗�M�F���3�Ȥ}���p�|i���}@���ɟ2��lL֟cJ3IY+�OdI���j�Of����~���65$���K�-���6�%LQL{(3���&�|m��>��K|��c��D�M�b&��g\93��+!V�SD�N,0�<x|��[���w���ͳ����t��(�x���c�|!���"��ʵ�\~�ݯO������^�s����=o�:�md�
%��Y6$�aL̟�WBsC�Ӯ6�l�C��� B���7�/}�)�N��sV{r=ݿ�O����M$y>؟L�8�7�?���/�
�fK���Vm���>�rv�4�eP�ϲ�Gqz��Q�5��c,��X[�<b'#�mc:驲;
���5��w���4��mƒ�*|T��.��̓��D���nJ�y�>��S��^��
h�aH�(v�a�NM��<��ױ��$&�@�Sh���u���rY�IV!�c3\g��>�#:�^/�*;#�F8E���c����dF�V�%yP'�6�z���8��\�N�<�͆U�|�2�7�|xisJa�����!)�����c���:z=���"LL�	�!*������1h�G�_����K�Âb@�(eD���*'#�$կ�$*e���V�����x�)ΐx�R�D�'R��8=E�yx���(�%�z�F�r�}�)���|���^�OQ���u�/T����{B�{�|a�>_$6w��M��R����q	���s��I[b.���|��l.ă�6~��g�x���VO�1ip}�:�Iq�*]��"���	P.汸8�6B�ٚ�k[h�B�@RTF�-�-�yL�y}�l%���a�Z|i��g�Sd7˪J�U|����a����Z���^��L���N�l�Q�������|�+�T	wT��j�#�q�ްJ�4�e�"�<|�DA.����D�xI�%�,$ʙ�'I���W��F^$��`+�`�Cf6C!�A�!^?���\=����l���㨕B6��p�^���Jo_Z�����@��8��G��c��z��E��o����x��B&����޸x�n5���ǒ�6@5_�����y�ϯ�=�P���lv+x|���ao��{�T��J��	7��C,�1����h8�h��O��v�o�G?�S�͛x9}	\�T�Z�F���@�I�=�w��﫯d��7*[����`Baq��G#��-|������֓'��N���ͣW�'�92G9������rs4�#�Q4`��B+�U�#2c��:���X^2��A��S�����.���t\_�Pi
s�T�7T���\!��"v�F����Mf�՜!V9Ζ���* �s���by^B˫:,Ɏ�j�ȓX>�����\"����dLR�9a����b�����"!�����,@�n������fr�`+x{6s�(�}��T�
&%)cΰ�)���^dp!���("1��p��iFk]��L�x�}r��U�b.�r�aa��9z�f3F�K�-+[GP���{>����4�?u���	�8"�!FwB���{yj��3�)}Ǡ�G���a�'��/Ip˰�)����1��X��q�5��(�S�����
��N]��D!����l�a@&p��M�Yي%���'�,T���CK9�鴣`K�Ϋ�Kȗ
�{�^{�Z�}����|��QW�d
WH�1E�����l_�z�2�F���S�T�`��q-�ǟ=F{@��P��l'3�P��Q�$�FN*[��~nB�J�m�X����/gmyݔC���o����@���;����
���#�X�+�a�}�ޭ,�ȶ�$�f�W���ZP;�������s�1��Y݉|�h����M9d�-,&.����*BB�bl��fv�(�"d1���Ο)��2��>�v��0^F<4r��jﾵ�S�i�:{�}��yLS<��&�:"�{O�sЁ�^B����s��w%�R��O��p���������|�7l��O���a�w��] �\�1F6��L�`Kb�0Na4��<����ZN���:��"��?�3��d\d�ʸu�:���`KT�y�"����1v�q����ǟ(ж�}I0�4^��N��̌�\(Z,(3��:�^lo+P�&;�SX.�X-�(��᠇V��9��[�!Ν��t���O^���g�m�(�i���`�cEL?�}��)�S��/�����_ȲL��rV�!MK:���u���C�ba�ʂ�����Zݎ�,6�Uvn���4��X�S�Ȳy>e�q�ͫ��͙XZoS�3W��0ac�[�<4�W���hA�D.�
�����}�{O�1z)��u0^+ߟ��`hOc!�jA�3�7�Ɯcv��Vm�
`�M�-k�6����2�aN��^���/Sz�b��.2-��X��-IH*"k�����[sSc���l�_��>f�K��!ǳhtNIK��cB���aƶI���vk�Y�M�8�:�7e#I�������=)ȉ`(���3W����Bs��6�Q)��k��{���~���������<���;9���Fq�:|�~qV�M���E1.�k�F(WR����Ffp�
&pX�q��t�U��᥻^lI�IDyH�bɂ���+��3#A�/�3)�͐"���xZ����є��6?W��F����*d���bdz��a�̔Jc�$*��P��m��=!i��
7!�%�2n��[טl����-���%r��mҳ=�ݾL0�}�i�����Y�ty��Z%��J［?���k����,�L�8�XM�O��*V�}4�^�Q�)��RB�E��)�b>zv�f�����)��?���y	�e��7W�C>,ܸx���_%x~���ƃ��ӏ��ݝ���h��\8D�Js�`�4�[SU]�a�a�Q��J�bo���,P����S�6@U��.`:�!boBN:����\�1Y�g��;$V%�Q�m�7!��zu�
β����3���Zw�ݑ$omm�_��?�ͻ��#)V�"�Ni���B,��7+�c«��GR�j�[xBҬ��P���+�Q.�(V�;��(�3�Sv�F>?���
��`(����0�]�x2�N�Y
�Ls�rCR�L;�w����� 0qe�h�g�ʖ��W�+���Eyc7� !M&[��E� ��k �[V��\e���T�a���oM&]I���ib��Y�p�k:�X2��*�2o��y ��H����[��\�U-��c}��^��ԩ)L�Z/@7�(x,;�/o��fS�������[��pSeIƖ���gm+�A��d�z�V�����"��ꖇ�#�)�-!k��^P=D}ƬXs�铙jltދ^��� r-�C��7{�:d�ɛ'���4ߧ6s)t�MY�f���T=�0b8F���Q�F�~A�2��X����+��,�#��+��l�`���X?�����,�V���;��޿�`Ds��%l�1��e��������IN+��FU)&'��-��s�;���!�,Ʃ������3��dePgB�_Iϖm����M1&IL��γ�������
b_�r�K��	w9��_#,�����>f���C	�{�2��s�׎E�
2Y�)Cʽ�f�i�*9�H���r.?TGS��\�FR�>��O�'������<�Lɫ�M��������&�i<bBG�TsQ�y&?���A��c��.~��h7"�K��.�g��Q��������G��V0�i^��+P-X�~��3�`e,�h~����4�9]�J���!�?=�y齯H�����v���j��;�@&�A�Qțl��;=2ڲ8<b�x���1=;�'\Һ�&T�Sx���O��Op��Yp���S�T�`#�Ghэ�$��d%�տ�k���ފ�[���M��7�NP~����ƒ�|]��޼��G�Qo��e2�i�̓�P>7M `����b�>88�����xM��H�l)
P�B�O�w]�l�R����zQT���y�۸}�.z���D[���.R���#E%/2��j7;��Ɔ��7�"$���$��d!��F�>rK�k��d�%<D��V�$8:�D�B�YO��
6a�`Ul��u��H�T��֯\:s0o�kgOH�eL���bX���R'�e��%i�YS���3�݁�!F#�[�M'��"+
BAH��)/�Ԝ�\3�gB��&��#��`c�W�0�Ӏ>{v���DHٌ���;��o�/{r�_�iUA���rQw��a�6���P~�'�Y��Ϟjb�&]^j���֤�gfGU�0�i�6� ��2MZ�l�!p��-E�(
5���ͱ��SnHDs��"
rd�k6�,��l�x8�7+0��<�"~��(UKx򬇟�����y�S�^��Y<T�6H�bb9F�3)�d�9���\4S�˪V��t$��k7���ssRj
�>��_�F1Q��_�FֺuĢ�*2a#'A�U����#VI6Ǒ���ǂ���5��Z^g�i��<�S3��3�<ësԏk��jb��̓?-fs4}�:��ku�P�:�A�6���u�֐�b�e��78\�_��eI�9��o������@g]z�C��1�P.���?8��װ��9~���0�����sc�����P,Lq����>�3��RuMc�K8{�,���G�x�׆-#ȗ��P�S8�?T넣�KK+dS_�x����J����������l�v_ 巐B�(�B1��$%v_�5���G���)��&�������Jκ��mQ������w�_z�<�H �Y��~��Y
L��k�IIX�&Vvq�J�������Add��D�d+��x���_���O+��f-�9x"%�&+5�d�b��C���~%j���q����}��I��=���ʹ �|�Lcn�A_}�j5��ag��i�je�~��M}d��Q7u4�8W))0��̌��&����g��&a��I�e ��f�1�z�c#s�'��rj]�6�YDH�ߏ�ΰL8�*4���)�7�3щ��tQq��Ó'���.<�d�2W��@c� E$�"�nտ���̟j�6��a�@�i�\SO��G�v��ӜAl,#�Ɂg�J�$h4�b��	�
��;�lZ��
h�
����4x��ph�%�+�㎽���AT���LT�R�b�a026+��4�����
��}MI�т�	X��Q�.5|��8�g�K�11k��Q$A�O
�{b��mds��a8E���Q�.�p�pG����&۞2��ۖY����.Y�=􇝓`��2�v�1B�x�im���*^�:'�������M�hF^�=���ynΣ��'�9��O&��Ϭ )�X,�4o[�$ G���|�\��9�2�9:�*�N5~B8�������B�t���Z�h��s�=M�术�dd��b��ugS���Z�JTˮ1{�Dh�6����1�j��O�\)�4|����f�@����O2߈��㠼��K�LȊcE�4�%"���|�	e�®3im�#��k5���J�7��⪐����^�)�R:�R4�w�^ś�\�Q������J�F.g8�9��_�����~��QoͰ�|Zm�j!�Q[f������҅e�p�/�p��i���س�`��n\ܼ�퀑[��Z;x���3`ڄ�6�Ԅ��Cg����n|�;{mt�����{�F��4��,��m�.�������&ݑH$3�m�5	����_a�%���9j�k������_\gӈD�l��f��:n���?��}���;�h2���m6�G�!�C=N:q$� I29�xb�a%H�&��b�z��XѓQ9Q�-DU��dZ\�'}T+�W�8د���*hu)���6�=2b"//.8r����+�@�mZV���u���a�6{G.���B�	g�<�T�Rqk���Ӂ�|��t(�5;�G�-��F���-P�Ҁ��}�0�m�Z�P�ʑF�`;�Y���9ִ/�K�I�p��u�y�Y�,�����v_3�w��k-�9���{y`6Nȩ��    IDAT�V��b5�˄��+�Ҟ������KQ�r���j��F}��B9��3�Mi6Z#�՜������-�c�DY��Pw�5.P�f�1�
�t":�S	���ȓ�p�*,�O������4��.�DBܜhfpfX�R�LH��6�� ���ɰ�vc��ֱt��8/�Z��Ң*�Z�.X�=Y*�)������
��n�F����(���v�]�o�λ���+��zT�_��3ԛ$EV�H��gB�a�� �L��&Vp��H�L�~�ʖ�o&'������),ͤaLT�a�r�]��|�h=K�̄�k�IKl��fy8⡑H�3���ͱ�3�Cc='�;SDK�8�*�c��#�8Km�FJ-!���/�����\�$��]bC;�����:�#�����901#��#�*n3P낤D�Yg��@��O�����F$jQ�|�E�J��I��p�l.�Biaw�?ŵO���#�͋�{�]���kh֎q��/�b����]�˦���3XZ�ãǇ��p 8@ǿ��
Rt;[�����hZACyyi���[gO]�v�z��?�?���|�I\Cj�3Ȑ=�I�������C��T�.���1Zݱ�����Y:�15���_��?���2[�t����E�B&�1���`�,���UT�C*y?��"�b�3�����|w�o�§ׯ��ľ	3v�e�����-�/J���$Fr"l+��:O&�k���C��1G"Bք�C��a�B��w1dY}v�T)t�C��7l�Fo�����:�-`mek+��`�6QGR/��-��$�ep�s �HN��A�^S�^�Y�����<���y�'
�R&�e��d�g�11	#�sX\X6��8�kg\%���U�)�� �Q$'Q��;�D�68BR���}��UP�\�*��g�̵dD���%�&�dc�6�`@Z���Lh�$
`�Z�{h܆A$0!	V�Pj6Q�P,�hy���D����
�d/��C�P|�|Č]�s�Vu��j���of�牨��Oށ1�=�9*�%�eF�R<Dy�jL�Vv�	3�%��:(	uj�}��Oa�6����QG<�aW��Sg6���"�N�ݖ�ǯ��kdr0�9��RO�/E��1����饅<�zs���i<y��O~�+�\�D��A�Ȁ3�3a�C�ƈ	I@�|8C��F�Ĺ��X�	�����.jmۜi�3�M�-���i�F]^^A�k#p#@��\w��xҶS���);�P�rs�d'�_�3Kz�I�dւ-��C�"2��"��4�`E��+�혼(Y�S���M pd�ۄ��^-_�a�O�v�E �MZ�d�x�Ѿ��0B��S���$�7�jҒg�e�lk�ǛE.�觐�NQ�ϰ�T��g���ɵ���;F��a�o㻯��ݷ/"㏱����6��3�Z���[WQ.U���n��AnnS���Jή�~@���b�`�x�����^F�o�O�8��>��9~~��x���K�����ut�t����r�g�l�ɳ=��{�;nc4��
ʺ	w�L0�`�R��3�U1�.-�w������8�pE��(�_�N�02f�A��$H�D��ĳ	z�Ϸ_���>�:ԓ�=�Ze�\���Ԇrs�I�0zL��_��E��h�U\>�w�쭐��kfo���h�B��\1B�*D���8�`�����i����UA	�u�(hAUE�w<sE��,-�H=Y/�HD"�C-[?�=����_��AѨ|�`����-��W�q�*gV;�J%�8�#d��q	�d<3[&k����ܜ�ѥR��q~YA��k�cs󞈵�~�/j���F���9�e�d%Q�J�NN,"C�pl�R�b�8�
����`�Z������)��/^c��K��U�#�GC���O��
� O�D���7��% q2������<��c��]�'��4,�� Tu��8�$��I�d��$d�)eL�Y>����X�ݞ#�X�e��V�pg0�b6�p�C�Do�6��C���aԫ#&qo�Srw��Y�//�գ��e�hL�a���*�U ����V�����m�Y?B!Jae����,�b�ϕpp<ƿ��k8�qv�ƚx��������1�,E-�\Y!U��
/�r��\y��1>��}��<����Y�FT�"�n$��e�����р�z�
&�T��`�?�JB`\P�s��K�7�k- "%/�b#;%4Ω�	M�EV��i=3O���7��d�ˢ`�u�yig�����Hp4���q�V��`˯1زZֹF�����'�'ҫ���̟ϓ~�\w1[e�|c�G4�"LM�X	�/ȕM�k���&u%_����4^�����5S���n���s�/�qjyQd����:@y�,F���8����aWk��w�6[�u���d�g0xz���c��z��d����{�[w��է�r�5,�Q�uĤ�>���g�q��.�n�1�He)��(r��KMf(�K�z�<���k��Z�.1k*��I��~���2K9�$�R}Y9��WAI6�϶_�Ͽį>�����4=d���N�#��	:�Q��m������[(�2��u�b���;g�M�
��0-V6�R�H	6"_��gZ��p�ƃ'�E��Vs��Q.V������~6�j=�XJ6V	�S�0�=|�;w�����wr���_qR�yT�
�"��y%�|퐕����PvO`;c�ud�r����ER����w��	r��$#��D�GF��:oc~:��	�K�f��3Y�%��NDT2cJm��<��6�t����5�5:�q�矐�N��(GJX���,՜�{�3�Yf��Ȍ�L�'�o�=�^��;�)�7��M�(�#�*�I�Z�HC(19�U�yM��}�
�U��d��B�Ct긱-�ذb6E C�7&�B5�Ij�0��Pv�L�ȑ�4�ߩa�m�xt��X�8�F�=�&*����l��L_նX�T��"[:B��ٳ)�C�W"�����8sz�Q����qp�� 6���O*њ���c�[&�#��*�\��I}c��Ks�;�_=�~}�7�-���y��흟W�U	c>�W'�H��Ԟ������`U'jc��$0Y`k�Z�k_�3��ҧJ��L#튴�8�75�}z�f|�f��b��V�6{���Ϛ��I�ı���D��e�`�������<�4�*tN�/�C�:���SxѾ�F
�q� �"��i�;��$2F'��8�b6@5�`s)�Q��X  �
����$���{j5TOkT��z���E4�{��cU��Fśg7����ճ/���l{����û��v��k�� ����������
�6.��+X_��Q�V�-��^�>{��;C��4�L�|s$�v;�~rA�9��)|�7��wߓ��$�m9��jr��{^=�5]rb�.��S|�i��b�����[x�l��|Et	�JZ=	,0�v��2X����U_�Ys�՜�z���5x�������(�@�[n�0Pp%�.G����R��ўf<G���.��J�

�y4[cܺ��nK#>�..<ΒI:oaQA?Q�QO8�%��B��Ǐ����[�g���8�W�p!*�S�<++�r���>��4n4K����� ż��~�F�L*rqqQ�H�g2hӰ���
�r�~�3�VOQ�76�ȃ@Pdh�P�0T��(�vɱ�	:���Q�g~g�h�y0��4��9�řc^��;=V}�l�J�m��in�d��|%D4���	/S���8�C
A���L���Z�����<I�h�b"�8�&�e�����������U�f���A����e��`�k�t��L&i�:�J~xX��b�>h@���l�����/��t��6�Q[��KW������=88�\���٥�|`*I�$I���픎M6��ʶT
����|>F���׮^@*[Ə�������T��L�
�	;�KV����}l�/3(9�l=w��B���e%����ḕE��mP�`d�jy)�Z�I|�l���߬+�cw(��LLnI�cK&1�����V��99��
Wv�rl�Yc���Y�b�����E���)��t9�竲UM(שK�z�0�����L� Kق��5[�ܒ��)�w�ѧD܂���fsERk����6�<��%�\3���r>;�`½`��5�t�>�<S�S�/D�\�by1B>���"�-9K���>=F�zJ����"֖p|@���5����\���oE��v�����[q�Qe����x������j$�8�y���{�/ �c�ع��UC_��?}��^n����z��f���￉0 Z�l=�������Oo����8����'47f���p��J�X,�̦��u�"��Cu�&<������#*�����ht&�.���*�qS0�s��%$��9J.�0鰫T�X�������9{\��Q�+��Pd�A�(CEB`�9�SD>�Qb���t��3]`:D*�D4��-�۝���n��":���$���P)Ve��>�2O/-��N��*��:�iB�������*~�aH�d��a~
pC����Ņ%7�3�0�Py��L:�66#TX��MJ%���U�j3{O�dY�9�&��w9�A��!G}q7��CL�!�଍���.I*ķu(Q���~� �B��	Lԟ�l/M����˔�s�..�X޼�t3"9����C60F;h���������qlÑ�d�c^�I0M��N�B�F^�ϙY]A{�!�l,EcBd��]*PE��Ƣ������nS����,z���&߃��l|eP�`0�d�����i�A0E�����3�)�h��� ܷ�~˫+��Ĝ,d��H�����;j�(9��D�o�k�R.��勨>�t�o�}Q��緞a{8�����d$�c�]	8Q���t*
�1*��R�|��������JYD�
�mw�FnvK�	�Fs�\�>�-l-S��U?[D�m]�1�O�bW�����߭�5m���E_���8�A���,D$��Q{Y�Z	�̑!͑�W�7ڇ�ny}�e#?J��{�`��cλ9`��L\Ʈi*�[�_��>٫���u�J?���ČCdH	$�d~�ӈ枑��$��)9�#��D^��:���D#��T-�L�`��J��%�Ì��CJ����O�P�VrX^1��N�w��9����;�뗿=�v���$��+������t��a�N�v:[ �lV����W��t{/D�������;������	���f(�H�b,UB��w�@>�8�?�:�o�P^@��������8���Џ���(�y�qt��fE�1�g��y贚h��j֐I�Q.e��͍�������K���Sl�P��cϰw@�,3WF�?;�)��Pd?_��m�
�d9��2�v$i�^��Ó�|7{�iVG�)�$!��
|T�D ��C�c��5�^o�[_�G�e}ƌ͈��;w�<*�9sk���E��w�꯲�-iw���nbkk˄}TEQ�F�d�<�� {�Y�˗��(��4����(5�E��l#7֚s�X��X]]>	�S��IH�!#_��U`eR��rO�Uf�"d04(�q�F�/��(�/̘b�鐥��?9��7W����Y+%#	��v��tGh�X!���L�)9�rOr諗�����d�c_��g����脄���3W�X`��4yA|��ST�d�xH��(�'	1�&cj��g��(9Ba??�O>�3�x�/.a>i%OF�:���@� ��#L�&�f�Tð�l8D��$D��7�xC�?�X(#�t�:ݶD48�� ��>+A��?l$�n��b��׮^F��s�VW��so�z���[u%���1Iꕣ?YΤ҃7��2F)�h��JAz�*P=�b�\{G#\���f����r�9P���Y�����	�7+��UU��U��m�Q�uaH�)�im;�cc�����-'�vd�d#�������D���d'�C~��v���c)H1kJ�j��ю����Z;;=���(Y�rH������v��N�B��d(-r"{	�$8YDC�B�%8���.I*`�ܚ5�OP�IH���Y,Us��K��=�����b��\sK�2�uǘ�*�*���nl\����lg��B�q��d�:O(����nw�حu�l�iH��f�&���i�R�)����%E�Z��s��D~�t,� ��S���9�Z+�����^( �o�Z�a�ɠ�+�3t��!k�bGs(���(v}"fa��g|rY,̗��</;��h�&	P���"n��ţg5ĩ(��h�EYO�S�1���޹�Eۄ�����AjFR� ���F��n����uk�OۀR�J�|}"�cB+�`�͇YbF1�'���C�pn�5T�%�V�p�� �`K2S�XC���A�4�Ӻ�|��c\�q���uC��Ɉ84�e$@2��6��L@��a�¾�	Jp�Ɗ��#%	7�|/�˥}�Z_��\E?{���ŚTU�z�F��Ϭ\B<��87�.w&�vDmd���j�^5�Y����
��a�,��EƤA�ɨF��A�?B��GC�26�z�eLů��c���Il�Ȥ��������a`�<������	1�>'�����^ҁ�ޏ���d�D�XU�������$8a�V������7sIh����ɐ��cY���f�/	ǩ1�=�B�L۠X:=B���|.��W�
9!�Ą/��ѷ���v���?�ҩ�����n[����=��y����v�ɵ{����h����SUKd�{3��'
��4��W&�=E�.��^̔dK!��Ratl�"S��D��$�9�G�r��ݾ�ȋ���;�?lg8�J&z�{]�e"�j�?�h9A�@�|^�7���J&�ƀ��d�n3"N��¦{�\�$^r���([1����-&la�v���FL���ɽ�*�3
ȸ@�����	ّɥ�`��FI{�	/�-�V���������p�kƙp{�m�x�Y��q�J9_h�o�+��P*�qpp�s�큕5���Xaܝ��Ҽe��D��>}�ʷ$�μ^��/�~��Hݯ�zx~�����=�;�J��.&�
�o\���3K�=��Ǡ�'����{��!}5mN��N-��l6��C|�����'a�/�>?��4rDMa�f޼ro~�<�i�^Ms��T��PU .�Of�H�;/�A?��3 F����x����f�z��~ܗ��+�Jշ����J��<��ND�P#�h";�9�F��H'v��B�k�ˌ5S[̇
��d�%	>�Z�=�+9Ax�Yd���o���M��)G�(��8�<VW64[�`+ȶo=?n<	����ɵ�%3x�ʤф�ؗ Gz¨� �Y� ~&�
�D(�Nkf�H�i1��!I��tc�VVdƤ���`͡Ul�����3��6\��>���T_ɳ�%�a#��x08�v*�R�&���1����Ì#K�Lf0Ѡ��";?��`�F���x��{�T��U5�^f��9Z�Ɏ5�=����ʍ���桫t�pe�=�[P�!e$H��Ȕ��q��Tc�'�]BK���&B��Lf�JV��|ҍ�����+G&�0����F��6e)�x3�\H�L�qAz �fs� ��_]�?�K.�G�Us�^��`6h�U-%��Uc���]|��������Ο_B��Ƈ�F�;�zs��]���BN�"�us��.�)�4�v<9�D+�fD)�c5��Ս8l����L3H�2(�bH�#�;{�"*�r�9���_��a3��^c��ZI�M����$���d>�<�����c~�\wR)�W�"��{�_��������|ȄS�ޭW%�b�'\��.~��VI{��[c�'j{v_����-� �"BĪSA[3�6>���kN�WL��aG��y:ak��Zt��Q�Đ���WeQ�hP�f����9�!O�V�����Y�,�4��?��ܼr�[ly����1�6�Cn��h���Gxv�D�7F��Ro��iʥa:����
֖r�+%
>�b���EԎ�8�Qku�|8�|%@>;F�?�G�^��<��Z�xV[La��Y=�f=�>~������1��	G<�fj    IDAT���b֯��h����(��ʢ3�����襤��⠉�㶂Y}<�2�]���J2$L�e=�Dd�L�����z�i�U���cu^)Dyp��Ii>�I��WV�U2S,�x�}肭�F���PXE�;{A�ӄ�	�H��/�>S۲ט������e�)5�Y�ҽ��q��"�:1��ef�Ԭ��A�}%�s��2s �Q�u�/TP��P����O�*/I1�Ad��Lt�]��*�D+A~N��s&6��5Slnt�w"�el�'����3�	�"��`�eyV���*&��$��u�KZ��1"-��Ĩ4��ıE���q�����u�������ͨ њV�eei�#[����N����kZV$*ڝY���I@?���1�r�$(U�c
�yX���"�������pt�ɨ� �G.������[o����E�y K��&�`���r������~��5q�E�?{�;w��8V�=n���m�;sx���z��`��l[�lY�2�2�R�Q�6�+������2���)��`��gp���د����v�Zl��$��!b[�T2�7� 7p� �"!�m�&i�D�$Bٳ�_H:�؅�`l�W�B	�Uʼ���L�ss-,�ϙn1OGj�9Gͳm�L(x�Ls;I��9�*�h�ڐ.���$���p��O�G���h����
IKY��$	��?��K�cR�&ɫ��4?Ϥ�r��R�������z�z�:+x�.-�iԔ��ڑ��� �եU,�-���>}��&ض�O��A�����g�Umb��Sp�;�co���If4�tQ��2�ǩ�Ν-�P�)�M��8����ė�����3|xg�o�c:���}Q���d� ��dD�� �{�~��U���0�&h �>�G39��P�!Ȑq��	2Q����=`簋��.���'���U�F�T��KOؗ���}�R�R�9�^�mHB���lK�9z]���I�'9A=�Μ=�r%/�_���������cDr���H68s���-�`IN&�lms1s�)в�`��{�e�e��3�#��{�h�4=m9PO�#����C�e�1J<��I�����0��[����|�$�Z߈��f}���Y_gfC���W�i�;i����c=2VmdD�%&�D���>��bJc���$���\`� W�b�����+;i\0F�ˠ����$Gk��@x�R�n�HU���K&cUB���ǪU��F̬7�$cg\�'O8bp[�?��k=C�V93��̭�B�d�'����eP\���}'��P%�4#�<e���&��B�@0�1*�"���w�����:tŢ>��L��R���l��M�&��C\	�h ������wO��������Ol���pӕ�#K��t$I�M���G���T/��4樍�I���0��qT��/vT��2�D�`��!gŝ��˞��x_�/�*���f���]�<I���6	nI�d��i{�l4/�5�����i
M���8�PQu��t��Ś�$9	U���Enū܀�Nzɚ�8��n�E樣�5�z$Cr:�e����K�s� �$|D���0�;'��%Ϯw��Τ?����=1�e�HT��M���Z2��<�I�P)��>��Ά=�2i� ��Q)���/��ܷ&ضO��^��ϩ���q��9��=�^�����}t{}�[C	���r���p��67K(WCm<���8(������G������?����%1�PX�sY]e۬^��=�9�3��/Q�q�Xl�0_�E+!�2{]#��PV��la6��=V�����4;$���$�g���,1��,��Q��tkٿN�أ#�;�p��8��qKQZ�@��`�6
5tO[В`{�ܺ�3�����٩��/�I�A�.����8���ӂ��ջ�f3T������;wo	6c5HC�7
:�>ӄ ��#�Sʐ�Ŭ\iL��D�(#�m͌
������Ã�+���R�;���V�&��"�lv�'^���8MǠ�/+$&P#mt���)N�����zU�}l�)AE=c��L���<P�Bf���Y��/H�
K����o�r9"��. �W�`�+�?��HM�Ȕ����%�I��0c�OU������"fdE
E��
�� %N�3WO��]�̜/� ?�*7.���c.������'�u2���Eш`71��e��j�Z.�w~�]�-.��5���|U� 8{��~O{�Ӷ9�ilP"LVU��t�v��bua�`{�8�/޿�f���(D��F�~$3�'�J�1�`KB!	S����m>"ҕB����}����I���EĔ1���#�[��I���Y�X���t�8��,�N�|�_�޷���bK,�w;?�(��\�I0�{*%��"5T���V��zc/�yCW�]�)�9Vpl��v��Hޫ�V$;J�:��ݍCʜ@._�qc?B���3�Y�9IB,�Zk��j6I��J��B�a�P񀐰Ia�w])V@�Z^�c�x�`\.��Ő�j&�Q҅�Eݧ�<�|��ߞ`�|�_��G����'5ۨ�cLGqVj����3��b������w�F�`q����2�����Q��X���o �M����������k��ٍt�9��Yvh�r�򰜌�(�C`���b���;.�|�(،��}7B<�Y���l�x�c������a���4eR}N�b�p�p��0��#�>��#���?�U��'��<c�:�)�{�o�?�a����r� ���H�@�Io���k25�������Ff/�U63jT�b�=w7���
6�*�T�<�͕�������۪�`;�9��d�,d�e�7���2�0�X�V'��ܔ<�%��C�����[ll�a�LT����Ɍ'bi��ş�z�v����u��櫆�-�&�e��ʨ%�h�X"��j���W�-a)4�#u��5�$R�k$��q�ȥ��/3*T	6�5N��m�j�=��fM���l�����|���S;q���_�����h�����0�T#.QL3���<��{ٟK�GV���J�
��������|��P���RNN�X$=��>�b<l`8�!�P̧�j�/����ͳ�L�~:��Ң֦z��!��9w�߳ic��Ƶʭ���$(�у�pzm����� ~|�F�YQ���^��L�fB�yIs�L�TT.UaN�`�-�J�$�Rk��?{GYx�yY���-��xb뛣?�ؓ`kd��~6�2����S�duN8��dM�l�493�lc5�Zk��"D�ڈ�b<(�!��L��!�h���QG�P�ZM�;!{
}�x��^��|r�9q�툤����[#�q�۾���􃵇`���0�$*\k	��*:���$[�D9�}�����/�"��$�@OK�q<B1��Z�圊a`���� u��<=w���^��`���E-xm�����/uokYv��{n���ŋ>�����L��T�(�U�쑇��O�Úؓ��˪*ðQeY�J)�)��d23��̈�����}{α��}_P6��I���@D��{��{������x $�����3�@?�6���Q�n?<������
�M;8>�ds�c�m�E���v�l��If��=+�gVi��xnv8.ٿ��ڋ��fY�R��Z��8{���mU�� `�:%J��X|�҅ù��� ���'��3ze�T�TT��@�xѶ����ԃYFw"t�"%�g&W��Td�@�A��{')���w�Du���!<�y/�^/�Ι�7m�r�5��;��?�L�VH�aDܗ"������cak�1#ڝ��z-����>��S��FK�-��U+ IW�b�)&2N;�j[΁V�R�f�}D�G��+�{�:,�y����M�p�<FUɩ�c�'���9|w8���9�.��6?r�A��������Nb��P�@<Qֵ
�M�̊dh�k"�U*@��橏d�Jhp���x]���pd(�糆0�=K���T�nL�йf�^7���3RF�^� �� �5�cU��F�$���u�?8�E�
*�7<�d\�`>���	�'#�q��"x�NT�
S7���m9?�Z� �w��z�����u����B�sC�����J��$MN��땦V��5����]���k
�g�f���돆�ޏ?��C�:�1��@<<V�Qe��ljd�LH�%sk֋��b���D�����u��=�{�2[%h����T��.���k�蒒��W�H�U�8gb_4V�q=��������V}Q"V|�=<Y�mDd��B*�(CP5�T��0!�BN��Z�1�9��V�P�Aw�t�"5|l�Pǐ�'�x��
aoݧ�û�]���~����u ����{y_�*��kU>ȍjŊ9=ݺ�[�N굲e&;��e�Q�?�����^(N}GI�Wlǃ{��|t��Y�R<���M�q,,[���b���|e��߶��Zju�̏��+Wv�l���v��v�Z�������I����w���}[�Vn�m�#3���B��rQ��uW��q.I8�i���D�E�����3 �:i@�1$�4O�����Tkh�%틍q��j̿�C���kG�oD�7[ͦ�[����*/juT��J,x����fUޅ�v�n9���a��_�;w��>��Gn �@�����˗/��
�yp=��X����Ū�t���Gr��z��O��+�'�-��� �L2u<=���n���=�c `d���m��
Ҝ% �SR�Q��;@�<#�'�M;II�0����0�`{
;y���;䷲�p� x���9�=��Y���A<Y4���;A1D8��m4�wԍ8N. �$ '��Hk�b���d>O���80�5AK�B�o���Q�:� ��>��>h��	R����qzB��$��V2�#0㑏� 7 ����k�_����F��Fl�lb�bj[[�
�g/������ݎ>�0������)΍�^��$���ܲ��4`�'>�����z뜝O���؞?/����9�c/����/�U� ���
yi�&�#�<p$˭�@b������NժMҚ��O�)��I�Ve��`o#mɽ#�Ft�d�^[	Wl)qݫ<XC�y|����m�އ=����<�H<9�LR;$j��<C���#z���:��4( WLi�N����b��I�&�s:��7������[�\�Be��#�Xm��>����U����Y�X��3)V������(���qO�w\o)�`�h�$Qܓ_1��<J��[���nm�{[����׾B�=%���:؞������y:+P�ALfꍢsi�Բ���RÖInO�ݱ/�޳�#`����f]�D���6:�^��m�ٝ�u����ڴR�g�o~d��~*Z~��e��Ś��Id<�5X��}�|j'�#����5"˹�9�	n,��#ӉMfSUf��D#��km�ջ�dP�ĎL�#e�\���l DX8��O5̢f�Q�m�_�X���
T����srK{�Ջ�sf�5Z7��Gݲ�~��C��!9I�[|��E���8�d��qcl�Z+F�y�6���4l<��P[�6�%�(z�T�@��i�=�r�5�A ��C��	i�(�LAͻR9V��>*B�H[�P��1p,�u7���,^	S��5�������e��^���ƅQ$�w$�����3��#�Qe��85ƹ�.�d�9:m.�A%��j�(�m6�T	����;`m��\@�3u)�w&�A�Lծ[�sK�9@{�G��-]͖r��X��#�%+��͞F�tg�D������Yi�gg�I<��B���X�n��kL�33�N �=}�tdY��c��S�m5W`}����{��Á�Ȍ�eh1��]�%��L�Xy��5փK����u�F��L�+�����o���=-�;o����o��=y�ľ��i{{�$��t��"��JR��*��u��@9
��[��5�=ϫ������Ԭ�a+|�i�P�26%d�h�RU��6�d�*��1܂��L�r�$¶�?"q�=����]��Z����������[X�[�Q�zCH	�0���m }�矙��^/LD�Z�w���-���\!�'��]����}A얚1(s|�
�4��V�i5|�wx9��}D�86�Y-x/i�`|��5k̈k�j�v66l;�Γ���K�u��/��WSَ?�WӮ��|�`�%�ꖯ&6���+�[V�$6�N$N�bo"�ۇ��A��� ������d�F�Z޹�작�ǟ<����&P荔`��7��8��Ru0gA��-cg���*[���Y�Y��NG��[�v��I�=}�Dd��\^��V��Z����÷U�
��ң��8X\���Rsqާ2��K�f�TV���l"�2���2
��PS{��+���	�~x�<xly�Y�2���MU��*O[[;�l�\m�A^=�t�`������ٝ;w|4�� 8�?�*�B��k#?V��Eo�E+����+�A�m"����®\�`/�Qb��s�'YS��?*.'�9�ĩ�N�i(i�������}*ώ}Ii�]��r}��t2�����s�L����Y�U����B%q+-���믬�/��p���	^��&$w	в*���+ �m<�K��;s�P����O����[��y�� &p� j�Yc7$�}�x�~I	��������۔�5�%�0,b���j��rl��uz]���;v���%�[�#U���K��^+�T�~"�x��0�[�k׮Z�:��W�v�LUJn��5���������
��h���dHJL��Va$���͒ժ�����k������tm2���F�K=[�س��=_��`�8��=��C�A^��2��%�}$��yPu� �T�s�ˇt�KY�n"��p!�8a�-�Yй&�E�G#g&"�ÂF����w�w�����~�\�B) ?q��U�.�9_%Ù{,��!E<���X���rКƈ�ڏ�`�$J4ė�Q�6t~r�@�R�:��U��ش:�~�����}�K#�Gw�ǋ����*�4�Cz�3��=�~�X���Fs�i��en��S{��؞<�K�Y�j�+R��s���pM\tb�����r���'�-�N+���
�B�
N3�Y�.qciTs�Fd=���H�`��k���];�ߓ��+�^Qvp��Ƴ�z<�}���S{z8��ܵB�ci�H }J�J��X����w���S�[p[0�7��=���nZ���-��el�>4F�T���y����;��ɾ�yo�B�\LN`�͍��ٖ�l_4�S��m4l<��O���fαb����h��2jQ��tN��J�`��BV�na���Q��T�]�l.�����a��*|}LE)�+�.��jB5�u��̼�z�B8���r�:B��g�|<����v��q��2�8��{r�RE��d�|oV4���E���W^���W�%y���^>P�_t����{]^�{��V��x+d֨�CD�)(H��_H�aMjlT���C�����G#��He ��P}B�A13�d��gC[�'���pa�&8@g�U��ʯ��_��6
�aw����c����g� �=M��s_\$����^}�+�о���mm$��`����?��u��W����������h_ܾi�*�l%��-ld�m��Z�a֪#l��f�n�ڝ��ju;%��Ǐ��S2��#���;1&�
0�� SqGQ!a��:�	�
#61�
�Q��
w���B�{�1��$�5!e��v�2�J�J)���G����T�Z�U��,�s�$�AŻL��P���_c� ����^|��A(
XD����|��pj��r�9B�POg�cP�k_�f�_�W�V�y� Om�:K��\�d�3��D��èf�bgpAc���z��U�_9�Տ�o��K"W���_[��Y��o'�{^�V��~�� px2�g{#{��������˶������	nO�"����r,"�*��r�Z�ܱ|U��<�    IDAT�V}	�c � R�����v�{b�Nf�=����N�LG�kg{K�,�@M�d,Hz��ڏ?�o�NVj�X��V ��f���:8��jA>�Pҥ�����>�
�h�%�?G�xriB���]�t�vH��-{�	�-�f�
��W^�3gvmskG�y��ؒ��~�kNL#L�o~�Y�ѣ"`�˒�m� ��-O��p�
�!Yα�}$��|N�`+X����K���f�Οݖ6q����4����S��E|�����J���"U�����Xc�Y��_����Q%����ݩE�Z8
�9Vm�vdR4!©�u���lY�7���o�b�h5�|!ש�p��c��I+8�+w��C`�1����� �)�KhK��V�N�Cu���aM;C�UQH*�?V2(w&O^�\��y��j�δ	�9����
�Ȗ�c���1:UǠ��8�`{�ʥ`DP��NO��x�N?�^��	��/�l�|���8]�xޒ�oo�޴Kܼ����7���j�/߰����͟��= 9@ƿz���ВK���A)����5�Ӭ��ݪ��F���Ǚ}��c{�`�`L	R_��$�.9���E�_9Ĺn�^�=D$��0R�-�U�&�Lx�5�_��($N9Ly@���_���f������ �"�Ҩ�be�ɨjjX]�|�F����h}��WR4�	���I��뾻�#낵��LN���"��X�ƹ�3�D�e9�Q�GA�#$����5�\Q��̂��F�(�7	�z�jG�D(��.<�j�v��X�\�v�����y�Kl����ǷV�ūX"M�����6�0�mu& �6����@��ş��2����}th?��Ͳ�O!5�"�F������,3�-=��e���O�`���u��U�� y���Uc�u:m��mZ�-t8�P'��@��bJN\��Ӷ�[V^���}r8�����}z�ЖŎ�xG�T��2-pA���UQ�3V����Ϝ E�����4���Ha	W���m�%#M�\"���G{�N�̀	9�6�z�k��E�
��?�o����[��3g�ѣ�� +4F<�X�Z�u��5c��>OSӽY9��,�K��}7�F� ��$`���j0����~�6�5*�h�pfӑ�b����OpA��ak��6(N�jؘ
���@�̕ۊ'^�r�D�T�T����F�Z�L_T�H~pRp�~���e��T���8ʡ��
F��Sqg�?�ONap��%wTb}�c�Q,T�B u�Z����""��Q��������S�<ز�U٢%�&����9 �lw-O�\�c=����]x�%a��n��k�snW�DUպ*��d,�(�Ub/|`k�ʩ�U�Q.���6?�s�꯽�������Q|��]8����U�%fj�@T@,��Ԫ���&^Z�f�ٶ5k1�*JAj�j:��$�����`m��%��E��^osmD�}WАZ�[M�����0��G��c���Z�l�
� t92oi;��g=뜩�����:ЫlX`�K)ʡd�Ϣ^-k���o�����A��-bU ��&�RD؜#�>r�	FU/���l�+}zR���A��a���a����j�e��/ElJ.���U�ɞ���G�W�Y���foKn��|��[7�~iz�y��_|r3����F���Sߖ��[MC�N;:|b���%�붱+�\�LrI�N�f�����5{�`ǣ��34Uk"p0^�c�t>����6�qߚ@f�2��m�j����-Z�<Fs�%w��7��HV����Y���ut�˙�6Z��w޴s���̓Qn?�����v0�leM�����[�%��3k��R��@[�
���!��4UOҐ���d�7�׉�#��:��@
�A�G�_X�d�@�U���z{����l��Œ��:��?U���W^Q���o}�4zA5�s�2�m�nI��X�LrEU-AWjTA�C��X��3a�3�D��<#���^�G�RiAؐ�[ � ���s��H+�l�6&�ScL^�EF�8t�`�k3���
� ���c�!��*��[�$��?A˟#��C�ÍĬ�h�|1S��ć��*Gl�&��DBX��5j�{�c"ܛp�r��Y��a���ձ��>�i�"����x`B?�]�HP�z���8��`��T	Da6�2M���rGah�%�p'V,�����4S�(��4�7޼fݍ�F�@a����=g��Ԏ�to��e��0<Z��U�sZ+W�\���?#��o�#�����;9i[����% �y �*��h0�S��@�
��0q{N&ؖ!;%������*x�E��,��- x!P���6r���y����7����L�Q�|�?PU�,�j��Qg�]�
܏U#���A��t��X�*ac���$t!��`m��TnE��`�B�G�-k����ـ�iv6�ђ�F(Ys��n�%U|��#+[�,|�J�S��%�6�7�����ѯ�4(�-&��v����0=F	[�<\�x�l��U��h��s�m*�/�������?+d�u�$�u��O�A��Jn����%��ڝ��:T2��{|B�^��4��z�}{�����3���lA_�U ��y��L�J�����ƶYַ��P��ika�ΖͣT� 8? c%�P1��D˧^.���}K��}�׮ٕKg���&ne�f�����G6^��
Y�\��	�����d�Q��D�� �-K={�6�d�S6pYTp�p�[�gFP�|B���sV�֌�Y�O>��#Y㱨���)��"�Hp���0�7��M��cV���9��g��cG �L�K���V��ܱ$ih��dG2#?
�lcfK���XD
���"��۽��"˒��^��[��.��1�9����Bҗ"v��6D�Ħ`9������	��Ke�1�q�9�~11e��Lj���]���-���99m Y�9���� Ea�W�����R�f"@,+8���S�:Yə��&��"O�4c�T���{��
%Q i�P��D�х�ܥ +7��[�E��0����{�+LЗr��;ć`+Y�׉Qȉ-W2 ���T@�mlO�H��iao�$������Aᨌ��@ɞ����e�I��4�΅7._�d�Oo*�~��oت����oڣ�TL?	�U����h!�E��Y�!�l{�V���t�z�ht���ܲ��h���M{��`���t�a���1����i����\iI�����~:�C��ƺ���5�9�`�Xɬ'�rjf�Ps�p_�2_0����-��'��Q���r�!7���ɬ3���(�#*|��fz>
�����U��Xʼ/ݟ�XBW0�e��8ER_�B#'�׫�m��5X|�����)���Y�[9L&�ؓbyZ���ZU�8~�۱��r��o�K��o����ӿ%ld��������喇����de��R��P��I)�zy!�t�����塵:���z��/ �4~�cзg�G��|bO�m�Um�*؄QHt�ಒU�u*�ݸ�ko�ֶ��Mf��I�;��aj�ζ�3�y����.��fqa�N�#�\w�%K��vJ���s�l6�p0����~��-{~0��
-b�B5�s� ��Ct��}a䩳a����	�O�	)2Kzu�k�sA�z8�	�ͦ]�tY���Z�~���5�鐩�U6�6E�:�sV��%}%�t���T��٭3
��n���o�b�fD(P^j[R�Eﵮ�-=�,����E:�����M٢�iխ�,	2����~4$0��(b����
H[�!px��`R�X����^I�M2�� Sͫb1��]1�!1a�(2�U�h5B^Q�_��T�۬F2�{$��S*��X����,fK2���'5Wf��3pQq�#V���X����ߐ\�s�x�u�xU^�<�#�;:b��K��_d���	�$�`E(���\@�	�d��s�;1jq`��A�IBE�\���f��W.)�\wv�֖p$&��h�+��W"v�C�R�z��=}������;����������S�{��ҙ@j[
��b8�`K�P.'
�H5�m��A56��͞%�knl�pZ����L����V�X��<��bj���g����"��hA8¯�G����g-���E�Uu����B%K"�6�V� �]V`D�#�l�2�@��`˺��n���~~ݐ�bam��@�M.�Ar�$/�Q=~'�N���^h���v�'V���5�c��&$��z�H��3�v����	�T��Ld�Y,���^����6z�5���`A���_�ǯ,��}�/���?\"����Ǚ����E�@}fa��B3��RC��I�o��K���>�
�Dޯ��4�0:3��#����j6]�m$���28؜��j̿���׮��W�6�=�<��d<������ϭֹl��"H��#��ΨsSa�=P�k��V)�v�®m�Z� 1����#��h�V��$�R^��|X��\���A�0��0	]-AP���+Z�1Jf�Q�QM��!I��lԤu,����7ok>����|ލ��ܹs��uF$ �K����x�@��ٰ��}��Y[��t��W�Ҽe�P;�J���F�hC��^g��ph�΃m�G�()���g��&:�@��$"���+rS�@5�Y�F���Q�`+��P�r�}�g:�ь��W���TL_�C�,r���;�3I��<!��7%���� Ʋd9�������K��1�2�8�!,����0S�=����#q�V�Aj�P��çw�Oy�分+k�!<֕*�����@^/[A�Ҧ�<�j�N���B����f��#[,-]-m���A������^ѭ���Z��%������ߚ�%�U"ָ�Rro�Ү���=��3+�3����W,����_���i_�3fO�O�-O��`�I��U��Wr����m�)�h�n�f�����wU�.[���ٓ�<[��� �dv=������{��~�<o����s=��DbU�U���P�g'k'���	9ױ�����/��R.��Fr��`�%����b�������)ϙɬ1�;��:�0� y@�,�Oy��!'��l#�JN����:�>��q��h �VD�<��9���j�G���\��Ҳo4���u�1������~y������|��P�V�:��rwґ�>�@M�vcSڥ��AvRs[LS;:Xؠ?a��Q�N�`�N]��7�ط;�6��9K�i�Vn>�&3�����[���W�VM�G:�x��c{�dh��e[��M��0��.���ۨ��2���[�3\��UHX{����'?��C+�:6�ZV�Ïv8&
fÄ���2X�-N�N�ߠ"��(ܸ���K�)�`Q�I
:P�pgϞ�Ku�~p��`8MU͙à�������s��Z�E�.Mb��l������l<:	PfA�6+���#����pEF?ڡX`d��#���MM����a�ڱt ���������ł� y�;�͂~0*�<�W`�}k�����Fuy:���E�H,����� W����&F��P�e��Xt��t�"�B��
b��]
��J�9bU˕*�
D�2.�H��HG<]�����`;1������< &R7���c�ut�ۉ)28/��Y�d&�sX3��v�\ki6��߂��7P ���嫾�R�dO�p���������]�~Mp�+q�\`��t�F�_��?9	l�~��[v��Ƕ�޳��'_ў�W��6�w��rr����=K����x e��*}���+�٪o�Hls�c�fɚ�����qj?������V��JA[�U��s�"-	��1��gx1�c�%���\�
w�YN���ˤ"�<�_̓�\�!��.�b���ps��K�b%�"nKh �%=�3�NX�~>��D��X�a��u��u/�P��`���z�gP[�J=O�b �ńcG��{�eN�/�X��^�f����X�ʦ1������f�r�k������������=9�蟭�
�����!=ە̓LZZ�x��bӅJ��c��Ԏ�����ck6Sk4綽�R�doj����l��Jn+��bw6�Z�h��`g��v�\�Z���-�bП���-����8�a��3���:A�7�
-f��3>���;v�Y��H�̤��"��Y2/��<��Z�;B;|o�$B:T*�H84�9��\-���^$���0���'��	]��A��� )F'�7���՘f���2߰G��|`�I_U������͒�W�9s�h�2�L��g�C�7� �$��4��=�?؝�ԏ�X��;�x֯M)���g%��� 7��TUO��`�����+`@G#j$�#ʦW��s1�cͽG!W^W�� {��!i�g�1�y����U����~o�
�&o]gNG��� �G��ǜ���	�5	I4�K��O��������`K���Я���8��G�� �-�,�Y��:����<��[��������oKj�Y�/ǍD-\'������qT�	�1�2�J���g6߱o��W�ٟ֬|�;v|���V`�.�|h���X��B� UoB0�t곲J9�v�j�.T^�>1�?}l'M[%�_� M斑���l�9��Gg�~XÁ<Gf�D�Z��_opHՓk*MO�H����E���e-�:$�"���B����������)e��-XW�!/ֱ�[ĶS4B q��e�a�Qg;�Jљ�p3��W���sv�s�sq��d$�<b�a�X�F�I	k�?����[&�����K]��l���Pٲ[��*U)m9�\��o����Ue����.��9L���pi'�T��>&�3
���6�e��R*qPN��L�32����j5 G�b�ԫv<H��_����RK�`;�	*�2�_��/�.J)�TZH��Vm�r���%���/'�E\��ݪf��g��K;�u�E��J����6�5P�l#~�A|"`S��̘��ժ/��>�3������������'���[b�GZ]��v�თ�i�k���ҕ�bs���SM&�y!|Tj�lѕ�����r>V�����'F�6���Xݬ��jF`���% �!�뺱6�(�*�׏�~Tp	���A�|Q�Y�S&�����`Wܳ6s�Z%F����"�؍"��|k�F��
9z��W�T�T{
��S�I;����̟C�Q�`t�����������d���%���Nm�ꅬ��.�v�*���b�^!�g�L�u�1��3B��^+s��@y��Qa0k++6��4�U_�K���/�g�W�v�i�5�B��O�B¼Z�X�<��S!jwe�,9l����[����7^�q ��@U���aa'''
��N��ЦOH_���k���g6޳���;Vm��O���v���ȋ,��[� �N��XBz�a�r	q�[�<��ulw'	0�f�xϞT,-uѨz�������σ�F���lc@�ǲ�I���$�ZX|���L�U_=h"�z���X�]�@��Yk� _�ڄ��D�S�9��fR�������"+�X}�ޢ\���H�D�`뭰Pه��X�ƹ�l�ѫ��9������u?Z��{:�*b�+3˱g��[��oS�r��oY��#�j<�Z���w޽�˪f_�=��������?S�]ev�_��pa���WTw�ҦK浨֪>�� 6��9�/�%ib�v�ڭ�Z�`N�Tb��`�an��M��3�=K�����Җlr�5lC�g
���z[���w["" ��I�k�����V��P�P�,��;�K����6��m��E����#A�_a@l�@�ID�����jc2qD�O��>{�`|'Ɉ=�������f�>s�����}�(���~��j�9E6�j�F0�$
@v��v6���g�������f����u�XR�Te(�ʖ`Ke��S��X�3g��t�uiJc��
.@ޏr�������U`��QbGB$�ŠƤ`B���`Io�W�    IDAT�D��
T��+jS��^��>��mG0<	r���BN(�S��p}�LƘC#A��6 �ཐp �>}�\,��@�� �D՜�QA 8l#��^k`wƤ�=�I�d�J5�1@��|�ة5�2ZF ���W��:#5�#׈��b#���U��g���\��C���bHu=������|�*�3�ۖr���ٽ��
�|O��I�tgK�C����w�`�s�����5�u�?��7vt��DGI(�}$�)�� 6r�sB�dPP���f�j� 0f�6,�-��~n�g��{��<�7O2�Z�D/k�х6ld�G�\*�p?_���9��;6���g��z���kM��D"�y	.0��S�T�F���U9<<��>�:�i�z�9�2�A�����=pZ�`�9)�Ft��	��>N�z��}��������1��w�w�j��ǉ�}�^L��zT�Z���b�����K�m0�\�}��m����4[��+ش�`����"���A��д���5KɄ�n80rY�t��Ҫ5k�uZ���K�������s�w�o�ꆈN'4�Ԏhe���G}[-�A�����O��j�r���Mt9aQ@�M�uˬ��&N��Q�Anp�9�����n�{(E��
Y��~�K-�vy�Ƞ��T_洚q�%o�y:FT��R|$f��H�7Tt�/^~U�맟�tvk8�y]4�����s��s����D�9ن��ܙ�
�����٨�͎�KJ!�U!޴MY�1?A���~��p�.�y��c�$�>%�oa�R��kT�����"T�Ő�(��P�d��������=[��xf0�%�����93��K��E�i�O#�S�K�s�3t��A@���~����a�Ղ���b$ N�8�{^���?�L�S�f�{Z:��,P����aU	k?�@မ�����ޞ��N�/��'��5�ly~w�?A��?��W��B�?FC����)H��/��"#�"H��������{���~�w����e�Zw�$y��2_�T�!+���Ņ�K�0,޺��=�G?��o���:u��?����iOl����3$�R��RT*���lY":��b���j[��Y5�������ݾ77�nZ�ְ�L����sx|p��`����9�8���C���/
��G��)9�PO������cqF�q�Lœ@�>�[�$+��'s� @��`�0Fa�u��ɬ_䙐�g�T�gA��s���26����X�эs�����gm��ݙNu�u����=�hX��&_��
�l�-Ux��� ׌`KeA�ʶS�}�*����<���{ 'R�In'c��/�0AU��1Ė�",:t�Cu�b\΀J��VJ(Mͭ^g�$�n�4��ᄊ1N�����4k�k�H�yL�a1Z�!������sV�T�Z�H�i>dCc."��r�rԋ��I��8�}nG#�r�bU=_�>�H�x�����I_C\� �8\��U#*|}���9�B�ς&kS��ʫoسg����u`	޽l�/0"x�W�/A|�\�f+��\�[+W���=�����U�;�ڡ>^�,A=�kyFeְZ��DF����Ҝ�om����l��-����j՘�c���P�E��$T���DR�&�&��щ?��r� ��/ʭ?9�L�j'���O�;�>�Ku�^	�Zfv2xu�׳A�6�Gx{4tK�j�H1 $elA!6w����Сj$�5��P�7+9>�"�8��{ذ���#(n���1�j�Q)�p�]��4�J.�Kg�=���=�y�KvC�mG�NN�φV*�#8ё~m�����땢ƅx=d4y=`�W_���@�6j	��r�y�[�TbE����~h�W_{��������ճv���������@�.>OB>�m��Z9��M��b�P�ehk\�������-/.d��l�޻ew�#'p?Kab�t��+�,U��eHR"�II���bc���d	7#�W"!ًATb'�*1�6�fJ���g%Β��8�Cr�}����ע�8��ƀ�gh4�(:�S�F��g+�r؃�G����k��&�j��.��բ���aooO��Q$OP(�<�)��?�9
f��:(�T9�^K)��hb�UŐ��V���7;��Lg�۝έw���fD�~���`�����`1>�������4���l4�m:�-���6��Ќi���qI�G���L�	�����2�WƆL��T �����X
yQ����Hb�Jj�ɉ�[�t��ڠ���C��{:X��l" ���ryl
m4���B*���*��O�ݶ� Z<�s�U��X���BV0P	�*й�\C$�E#:H���D���-y��UkO0�g����=�\�Z�X��!�\�xή\��jW"��JL� �f��ݵ�~�#��届�h�S�c���_�Ě2��v�z��F�������SBx��B��p��C�x:*'i#�]��{@a,�����q�}� �a�bY
X^ҷ�y���0lJzQ��n�CS3wh᠈� f��H���" �"�À@�f3��:8��*�8�7}b~3�
���[�X���"���+��e������0YAgP�&����s���� �1�?�?x"����!�*ImUk\�:{l�-�ELבKd��Au�%�aCK��Wǖ.-O=c-�,Rf���o���v�5]?\��ˣ��>��:\��Ϩ7^��R����@�{���G�����������NN�A�m69QM����"hy��j�R���W�NR`�:m���
啵z�&���w������m�zM�?��`�XL����'��5�N^�T#��z�
00�^H�9D{�$�99�t����?m
*}��V��T֑���=SO!��8�b/TO�Ǽ���Պ����@#�N����=1����G���pc��߱JV-s%1)~gDs�o�����N�}�t)g��s(z����*VQ�lYۜe�)�c	��J�`ۮ5l����ݷ�~�d����ۓ/������X�MK�2c�s�0�LSU�n��,S�\��1	620�f�Ԝ�>�m@� 3zm�|i3tY!,dd�.W��]rhn�fѶ7f��dxd�<��F�*��]�O	�f�bU�(�k�#19� �����xH���nf2Q8���֝���͇6]���rŦ���tQ�����<��1��E�ߘ���\㴲�T<�B8�a\[�ѡ͊����sd�9`*����Rb����!�r�-�F^�K�6_�f���c���M���B�#�Y��Fް���Q�*A�K���ӯհ�����>ǉ����_Y,�p|OAʐ��!�#6B"����ܨʂ����%�~�r��ޗq"$3gUN!�2v��OЂ�a��mHD��T"�>a��b\�� �;����0Z]�����xy�3{*M�0߫��X�޻�wX�IP����7s89���׀zW|���_�B���v�d�[�ל�J���KW�lQ`Jӡ�k�X��T�R�ש�^����V��m7n\W �7Ѵ�đ������H�R��	�������=�����ڎ����v҇�H��cC2Z���V��v��-��rj�݊u[ʐf 9f��C�<��/�6����Qt]���]�-������<C��2�p�V=��O�}W��������h���j`&�L��\s�#�Ą���,��9EI��D!
)��U��G��[1<�8�� ύ������{�e�mA�B?7
{����woߨg�>��[�A�"Lf ���"�"Bʞ�x�� ��/���0J��H!l����שlw:��o�y�+_�`;>������=Kg�E��x��p�ԻX%���&SU���8Ԡ�3.�^.������RD� �`eaK+����/ Y�؏Iٖә�Kfv��ɭ^�[���x x��ّ+�|��7ZƸ�xoe8~έ?8��ڹs�b�B����u��������'G�cZRW�P�90JB����;m #�j�j��&���LR�.!��JW�UVb�m�U3������v��-�4#��/x�<�nG�v���:�Rq",�
�%h"�Ѳ��޻�9L��K���$�/7�Rݰ�#F�A=�����-kw��r���Y�s"G���/�&�71'w]A"����Ke�#�d����W~��-CV�{�ڈ�Kz����{�^�D_#A�=i�(8��U���SՃMl�yzF$R�+ t�^�k�Ȧ�qv��j�0[�PS���z��G<��<�HO� =A0��C�s�|�@RT�k H�ߥ>�<���|�d��bƀ(@��������f�n��,�����,)L�}�#~�`%c�����ݯ�#�W�+��gP)!1aJ��X����!�P�l�=�Ԯ��mg/l+�Wl>��G?��1�7�1Lk�ϋ���f��ܶzT>���mk�i5���5{�|j}��N��6�0��G����^S��lyQ�1[�l���d�,�|_x���[�&��L�X�uiB��_Z$�9l���e/�A
 B�ާA)�ޥ�$/�\�ڑ��y���ft�bb���IR2h'�������yO7B�T�Pp�Ǌ^�Ԗ�PW�,z-~�N��3G��5<�z��d��3�Y�>k��I}Z�5T�8�(؆���o����_�`;=�{�?8�Y�����S;ҿ5+U����P}<D��d�1腘K:��C`2* U�d=�@0ue�mУ��Rj��銾����3kTgV-d�?�9<ˋ6��`�@g��\B�#+��|,���g�h*c�a2�to��<ٳ� ��$�R**#�;$�㐹�/�/!K�2MX��DN��{�gt5�S0�,�^h�ݶz�!��ٴ�w(��s]F-ݍ�z�[-v�P���U��Lv߶�����\!1[��-�v6�TٲjeG��Y�BxU���;i�vZ5��X*3ň�R)3$ý�e�(���pZ���,vv�7�/�m���fCB��Z'ArQȯt��� Ar��Ug����\�vz�=�Z�$X��SP��$%�&��KQ��#�@�����\�'O�ĒY�-�xIBR>��,�����O�%	P���N�*~�đ�����E<�4�ɜ�l$n�q*Z��au"ǉ�������MF��ex�-E�by�W� Y�-�k�u?�^�5[ޗ�J0���ǵ 1ar�JE��3���M��������+W�l�\���[ߵ��Ħ�5d91d^?S���U��x��eY�FICЪ�mo���Aj�`i���=�/Y�v�X��Y;*P,�w�,�YA%�l�<6m��!���b=2�DX��U�����Ց*��Z�D����*U�/�t�\�z��V�T��q�`�s�$�Z\�Ο�u����#@�g	�o�������j�l�x��C+�{�^Ism�
����;s�8V򲲎L}�FQ4$�d1at���:���nT)LX��p��E�\��Un�;����y�Kl���t������,�;R�/N"1vSc3]I
��x:���[z�E�F@j����꒢��C`d�񥚕�[��Irv��S*�ls#��NjMQ��t���pn���la�y$��U�U��̶w��Lm:����b�b
��õdG'c{��=y�\3Ĝ}�X����y8�=�zE����bpǉp1�ez��@E�p�yBH��{���.�7� ���g���(�R�+�x^ockC�(�m�ӕĭ9&�R��ۧl�~��eT_�f��ٮ�la}���M�-Ǌ��mH��l�~w���P�B�����R��z�3uV~�lL6i��S/��`e7�w�g�3���RP���ٷ��`>K��dQc,QQ���<�޷��ҏ�ʃU�j:��2��D�D���˼GE�$�}�l��~�p2�I�q���PF^C�T3v9w4� ����R�	���m����������	cT����
���0YpC��r�^�Wȅ(~QM-m8x.�x�kWR�:����s�e�R��T���~�W_�����ZE��`�����`�3�"枸�~p$B��Z��.�6<~d��~ƶv;���-{�u0�C��̓B[��@r���-gV���Ɍ.�:%�h׭ݪ�s[��w������̞�W,�nل~8s1��9Sٲ�X�be)����YnK8q��c�/A�������'��ȭRP�	6ҏ$zb'W�G_e"c�2�$R���ɍ��B��W̰�z$)� �[��cm���/���$�U9=A��T�z�K^8%Ϝ`*r ��0��>W1Fc�,"��^ˮޅ��*���<�1<���j�P�7[贇`+�����7�|�KU�����ç���j�J���bn�'�è������P�3�	$	*6zQ��l��w�B�B�	�%���G����g�"����K%��F�n/�Vk$�Zh�l���~�Rqp( 7�|㙳;���h6xo���6��QdϞ�ٳ��b�����~��&<0g����M�}�E��*,�͗�����T��
D�Ytڛ�|�О?�w/����������-��N�m�=�F?X���/�>q�n��}q��6s�[`�e�T��T6Q��ա:�yb�M��w�Q涒�%g �W�A���/���^;p1 �vL,��$XQR�V�I�����XK�y�ah
�H��C��՝8�csRޓ��G����г')��>�E/��^�eBH���Y(�^r�E��L_g#����P����6��Fk�v9��e�DT����θ��%b�{=���{B�uQ�`'�V��RU��!�魈 Z��ǫ4c.�bW��^�']Ml<�9�o�-͎lQc�!xLɹ/��޼j׮_��ft�`�Kң�02����Ib7
*�S������vrx׮_�h��7쏿�W��1��:�S�J��VX(�B�B��V/X��qa�V"�^����jf�̬�3�я���my�g'�(�"�~�E[�!~9<Jo�?|d��y*�ٿ1�bR1�-�rx�Tf�T��������}^#�Y��L�V�G01�b������5�-��H|lY����kFQ��i!N�n`K��.��^.ō x''�)���D"KB[����v�=\�֠0�ďJ5$�}�&W�V����qKȋ�WĹ_WwSV�n�uT���_��olII~;��UkB��5q{)���z^�z�k_�`���?���t5��<b������Ȉ L���{�g��[c�g0Z��x��n�8��_6���%��%�ڀ-�:��-�;��/�R�Qh�,?�B:�n�fۛ���,|��Z�1�����m�j�����s�n���&��+�/��* ���`��ߗQ����SU��f�K�!�W�D����Ρ�e�I >��"�ܯ�/��8L�*ؙ�K��������T\Sq��ͭ�x�����Joon�GAy���84~�����?����8�t��ͤ�U+�5�@M o7z&@�(������n���}��=z����-�|�/&s`1x+�g��6�*���iK$}�vZTZ$	NHsWe��:�ټ�sӳu��,�#����'��T�\����#T�@ty�7���(���.F��a�Pc�NN\2l{G�����I���~��9 �%%��
��az�Q_���˛tА p� �* �5��@�$we��T<	��{b����Q��i:�l9�l5�4�oK�uH�Tě8��=6����ץ �����܃{������Z������+/�|޷������+v�ʶ��7�<A/����CW��Rby�ąS��XF��������/R+�m��"Me����[v�O��ɨ��v�`I2���~	��W�"�zz]���F/Vu�Yb�,���G��u�Z�Jƣ�MP��6�3\��jKV��P�6a[�@]I�FU�r��*2�By���տa�9�"B���1[Y N}��(#wb+�P�`�^.0;����(�����e�    IDAT8�V�,�"˚�O�at���9��iD�@���gl=A-�E�N��Q��P���	�`�m�l����Ƶ7�|��>($��	�Kv4���`*� ���n��l:a��e� x�Ɛ]
6����8��
��\�o5O��Bu(�!�:*�s��V��6������ll�~`�:�M�N��[�6um��L����H���G�d�M��:k��� ��,������N��]�'*m��Z�_T��LE*-7h�����@��sx�,6!s����w��IZm|3�=���������������ST�:A
�ҥKlggW�������&CU^2���oݲ��﹬�lŨz`6�-I��ݰ<iZ��q�58��@�rq��4��[��uͼ��o�D&b��D�&N�����C?�~ �ϕ�D��`U ��/Bw�9e��A�<�"\����d�0�A�	�q�qxp_�_���za]�2r5��<���}���H?�Dj��o:! �\.=Q��3{���Dq��a|���W�)���p<r	I�����INt@�2�u�`�q](��A��J%�}� 6@ɿz���r5�HRH�ѯ��f>�����˱z��t`��P$� sG̒��r7nܰ�W_*��L��S�"��U������P)rxVo����'����'�����zm���[g_��|ް)����&�+�ǰ�C���(%9P�*����ZU�q%�Q���۰ái����
R
-�-pȚZ��2�<W ��OrØ�dH�l9�sUp�q��Y�Q���g���D�-�-Y�浔��`��n�G�c�T?�odYc���5(� Zͦ�����Ǹ��'�L-��"��%[�4<_)�'��ޕF��s�&I�ѵ���MErL�f��%I���.���%��	�����[=�^E�U~.�{�����Ұf����}٨���	�*׌&2D1Ё��Ƈo��%�lo�����j��@F�<�s�ݪ��/�Z\Y��Jeh���r�����'4�]�b8�ق��t,H6)4�D��ק�(d�m�4+r����ҙu��̤!<�/l<�[	vZ��b�J�ة5��q�����nY�ճ��M&�����_���yO�l�e0O`��q=**�J�̢ -]-��{�r��?�3���{��Ⱦ�d�Ξ۶�rd�[mU�$��e�{牌2ƤJjp[������Φ]�pN#@lbƅ��`��]��������}d�>v�~ym��}�6I6-)v�LƷ�����2�u���a�L#��ҡ��rY����@J�`��C3jY�^-fF��"���e�@a�!4G4��_dL�l^w�i��׉��r�-��ĕuf@�w
s�u�iĈ 0$� �\���h��쎏�l0�#�L�Cz�Ԉ�d�{��{-�P��>B����D 񶂣T�y���G�J�gX��^gF$�� �_W�NbA _F 6S�U靺r�ˋ I���T��IJ�eɚ"j1����X�6˙#瞎CoiG�wn�� �K���mwT��FV"p�/�̣.g���?�����C���v�e��ݻ�����+v嵞}��߳w�m�Lc7AymnE�~�(2_�Z�b���YͭE�V�kb�&�?/k��ߵ�~�Ҥ�=��PS����	B���BM�����C�$�x�Ցk�A���Z���:�BL<���tlc�e]��y])|	>��b
"����$A�NILy����U���z�����Q�4�|�kEBNU�jy�p����g��b���k�f%_���[�0��(ơD&�����'D�%a�7<�U�k�x�Ǔ�޶��lA\Ԣ���w�~����H��J����F���&�6_L�]�����Ǝ��h?#4T������S��Ð�6�T����"K�E�M@-�v�Z��M�G6���]��C����3;�uxb��P�C�0/�-EI�!�h��X��é=�;��޳��?>a�����>R`I����d2b��e��b%�ƫ��k��b�L���s��g�j3�<U/y�����ⱂm��t�-������ �`^�↍�bn{6L�~l���pg�
�\;V,n�:�{R�b���a�3�U �Md"^��+Eyh��
�ed���$���ѧ���2u�-x��zCd`{�qr�`1����o	�5���:����sU�I�;�
�%�#}S!0�ɝH6�Fmze͆����NX�#H/4�ZW�^���0k?@�1Kƞ�� ��Ҡ� �G	� �g�l�h�7:�p��W� ����\�D�q�g.��,��,�S��*�!4��c�͹�H��g���`�ҩ����.c6�7�<�Sx�1�M�bckS�X�ޜ;G����=��\8L��>e)W����]����Դo}�;��.�Ŏ�Ǿ�4C\`��T�H|�dV�fV���Jj�d�џn�%&r�U�j�c�����=;�t,M:6�F�=̽���M �D���W��>��vd���S�E=G�&���aݩ�;�g����1��h�/*B���Bb'Ғ4�Z�*R�n1ⷷ�w�ێ�v�>V;!���:y/z� 1�Ai��P��������%k�2m&��}�P	�K���(i�	�?>
�{�+�Vα��-�-1�� ��>��f��{D����~z���__��_�?~e�\�Ç����`�?�'���P'�T}�����>J���F,})':%$� `�;K��؋�c�"fY����h��'��]dTa!z_1�4 ǘM6Z�^����+�Z���X�������/�n0�](lI^ck�{��ר�ы=�(�0��@�Ǻ������XAI�{��
0 ��l0��Pb3I�W�Ԫ�ҭn�zu���{�W�������3v˜�bZ�U��ސ�
U�U�%�C�V���~���=~�!4�ZV@9ٲ��|ݶl�"�%)����1����#�T	�y���`~�4/t�T�hS��E�X蟒�/pb|�|_��������N�䕠��*|��n�k �0�C�3]����Z, a�H�jv\��C��HO�?�b�!�����T�F���Mܝ�_�L�~F�T�̣j��`���y��W��Ș�.�}#8z%��#p�Q^�0��$�t�.X�0vL�@B@EK� ����[i�`+/��q�RkP��
��5Be�����FW	�ܯB����x�X���g��fQ	,|N�U�������kg/5�/��o��ܣ���A�l�I	�E[�4h��`�mf�Rn�v�z-k��Vn6����~��c�7,/y�%c��H��sD�g�A��y�ǕL�,�cn̮$0������XDvm<�i���Q�����b�]D��&�J%T�fl	������y07)��O��ԫvꜼ�3[H�A�$ [׌w�b^G�!�p1��Q���� ē��$[�j�ŭ$�xZ�G��=� #
�[�s�y_��֞T���E�r�7�V�H��`�=�Rۧo���y�?����lA��\&B#�(�r,%�ܸZ!t=a˶r����m����?��þ���k�"���4�4W�YX��U*.m�?�A��5�;�۴+�q�i�x���`lK 7���6�,O��(�/)( J�ϊ��ha�=�{���Eǜ0�N�3`���l�� ���h��m�Fx�lf`���ARp+�}a|��(��ٞ]��+?��xa��e{�6�%TJ!ؖK�ol�$��$|Z�<��ѡ��k�:6�.�������]�!�⤂l�%2l���4{����d���fϝ�Y���gϾ���{����B�������aA����4B)�^T BM�;U�}-w�qO�Xe�GɈF`g�@a.(�4�B��}X�-�!g$�
�z�I�y&V�Ι3�#
�s��VWBL�R�pJ�u�ݫXaB.'�q�as�H9Mmx�w([�G;i�9OV�����Կ'��!��鷡|��^�}���a`�15Q�	�|�E�0`h��H2JZr�`+)r}Y�������:t�Z�^�u)Hai���^q�{� N�.8��r"��IZbR�۽�(Z�ط�߹h�^�)�޻��٬fh�g,�[�$r�F��
�i��.X���R>U��L#��v�J�������}�zb#C��y�����j���p&��菷,
r���l��`�~DYJu={�턙Z'/e�&Be�r�+��\V ���M���Rϑe�хoX���Z�2b��`hds��f(��}�zJ�p�
,d�b9!��力u#�s�ڋb% O��#V�Jf?PT����1;[�b����/�D�$:�`bt��p�k;b�ly)E�]�Q=Z[�l�OT��\�B�mw?������7��<������s������zbWds%S��h@v(O~�[��H^��?�� ْlI�(��p�n��f�ǚo����|���s;~i�/P�U��=����~��k����KA�q��[�{f5��F���#�6��l
�(Q�$ifv�FE�x�=���e�A�k�62����aw0��*�`L��E'�L]J?�u��y�jLl�k���e�c�z�j/=�e7n\��`d��޷�,�ě٠?��틉��0G���p�O/�E�;
��n;y��=�� �dq�-�F��G����`�𣳑E��̝��6Z�h�zޞ~�����ު߰{�����Gn.�	Y6��]��gW�\�j��|�-�?�:=�v���Éݿ���~x��~R���\�q|>�2�=����8��\�`f��N�����V�PE�S�/wz���$�x��K�A���\�]���#Q#H�j�ReF���墔��sA�X�4Q.�Uo�c�hR�� @�S�0Ǒf�?��\sg��5���8�֥*�r��!J�P�8����bBw')�H���! �g��
�]�+�dҸ�٩>���Qu�3QA�k6��9ZC`,l���ji�y�I���࢛���w�0	#=�%vrKrq��E*�C��q�	{�[����s�
Q��2ש�v蒔�&����C̵m��6�ۋ/]�'�ޱ��ڷ��w�� �mv)����Է�f�V��6�Y�����ʹ�U�k֪����V���џ�>��~�V�-����#㾤}�	�5\
���<A��%�����Fp%㞱�=Y�
[PI��W��t}k���}�~D4k��t��vw��������W��[̵go)iJs�<���%��<�s6<ɞ���(��i�_�u�Lу� ��Gos�8K��yz�l3%��b'���M'�C\����������I�1���xo�ZH+9���zS�-�wjh#�㥍�&�����Z�W�%�h;]�+�yY������%� �2���׹ϩ��k�T�la�3�^.sѦ3��R'rP�0RPJL�d�<��%��M�wvd'G��_-칛���s5�v�a��X�(�'�r���ߛ�N��ÞCp?V���������V(���9����u�r�S�OS�x&�:�P�,�|�:l�Ԓ�AB	�>�R���F�`��S�Q���3O?f����Ù�m=mw���{l�Y������r�R��vw�T������v���z�������{��J�{��:�N2M	y��+awR��m08�ٸ%Gj��f���4m$�W���gk=	z8T��� <��5�fnV��\W*C	~��9�g�_'<Iu2��h`�w�7�z�Jh0�i0\KF*�W����aμ�z���}FP�=��5j5��L�yThX����ɸ�>_��U$�G�W^�WB�+�=��
�I0r��F5�.v����/����J����wɓ\��ֱ���P&�*������� �=�%&3ȼ��p)�)�w��UY�]��J�YYUY29@fs�,�������&B����Y�>�n]�Ǟl�_�o���f
����b�\�D���#U��e�\�[�<�z�@��F�=�W��4����P��5��2Ke�HQ$�p�b}�(���֮����}K�G[�4Y�I�E(W�h�w������($ԻLm�h#��m@eI��9��-�^W�%�l�>/p�Kz�.���e0zr�Dh{�(���4�d��`����T�jMb����!Vu���5$bn�'�YflK87y�8':��s�IG\Z�ް��&c�R\��agk�8�Hd���,?Fީ�?x�����8�9�B{�G���dr���Ei�? w��P3dzv����N؍���!9x?rR�3�(�h;4g�}\zN�2�'��� �z��N��:>���}I~���孱|r�>mu��Y<�@����\ۙ`�"��Z"L�K�pj�q��� ��?z�Y6|��0�!���ޠ��
ST��|�T�J ��+��Cw��
ykԋ���={��E������ݹ��n�y �r�b���}]ӌ����T�����n��?Y�MvvұG����e�����Ӵ\q�
���lK/mz��Ҷ���[ڸ����Z>;�j9#r��N�]x���^,`Q�C�q�l���3�J�XC�A3A���X�;Q�͹��7�8JpUrrs����d��?C��W'�`�!������<���_D�af;3S��y�#���䙤�D�`+Ͻ���mR�A@����؅�]�z�����ݮ#��j�����\��j}��SHT��d��"�$ssAk|�x9.�l��j� ���e��Τ]�C�26�5�>�B����b,:$�ϻB���(�������˗܊.��`�$r�z�wY:9=�}���T���b�dv��m{���v���}�߶�w �ԭ��2>7�ȏ-�b[S��FTAТ+�䐉��m�7�$��J=o��=;l���oܳ���`�80�d0q�Z�T����Κ|�N
�毒̹����:�w��s�s�I�\b"�H�:Q�^)�t蔽0��	p�
6�?HĻn�m�^w;���`�>P+&���5((���!��珱����}~�d4�iG�3����T�En���?�\[��F�ux�{�$�ѣ��)$'%�$�>��ﯜs�x[9�7B&��9۝Z��+�^x6�I���1��B�m�������o�Rd.�ӝY�3��<2s��d�Bb�9�J
6���~.�6�1{y���xZ�;�!�2h�~���"D�J��eb�|6��{�cW.ڭ���N�yݩ�{t|bC��H��C+�D�>�?�Y�D�K8��ЫE7f�ݫi�p��������N-W�h�x
d�>M�c�%�8�a�!���y���s{I�0͢j�����o^���/X�s��_._��۷�$غF,U)���7#7�5�"�e�XY1�?2
R��������v|r�Uؔ�ٖ�,�ٱŪn��'�*�����f���V�����׊V�#ߖ�:D�\A*�S>_�rի]Դ3e鵻�;c+0J]�	B\o��Hd��H��A��$�v���������9'�`3����!����^n֪���@�s����{�~@��Ęa���G�ZS�sDߘ�.�T�������n�3&P]�xI�-��1 >��Ր:���Y���~����F	���cu�d2~�9$������>>��>�iJ��a_����JCY��hb�j]�?D�C*ps{��O�g>�II9�7-bL^��ؓZ.zZ'�'12HJj�������G��'_}��.�+_������a�	ab��$e���i!k�:�^lk��mղ֬�k/ɜ��U�B�a������k'ݪ��UL�%��ytL r��ry�ۍ�5��=�_��\��d���Ԭ+���6D��绯�5b�Z��TeZ3�iO���O00��`���xe�Ιu%Jk(#B����,JW�2O#>J*��.3��6���U�äN0S�M�FɖRo�\����'���\26Ic>⌤y{΄��y_�_������DX��/Ir�@�x��ʺf���y�sϫU�j���3�����0���׽�6��dP���Z��ffa�RيU)�=�����7�3#��)3�@EI��bӠ7T��3��*�s����g�����ՌtZO�އ�ۓׯ��/ܴ�bdg�Gd�    IDAT:�����c��ﰸ���`k�{>U��՚ɜ�+Ws�����{vt<���]�B�"1�q�2˂K0.&�Q{Q�����*Y±����(�i$���瞹jOݼf�Ή�F�&�� ut|*�*�O���p7�.��=��������N�G�ְ��C{���t�)xi/��G]�\v�t���2����Y1?�|v =���̊���a��2H	I*�ԃ��>A�x�jT��B4:��K@K����"��H���x	��刯W*u$ -%/nc�z�e'A����d�LU��F���C>��^U��H��^ӡ���a�MA{���CBA-'I�1ZCB�u"��~��oi�rU�'(��T�d��u� �Cu)z�\d�Թ�s˺���Z'RL�TA@�k!4���W69�}o�:Id`*������q/���O?i�z�%k�+��`c�#b�Yh�l�`K��{ i�/��K�v�&	:g؋/_��K�P�.�Jf9c �@��e`��L��Zw���k�0rye�RN0r�Y�j� �(R�}�Ck
��|N�VN^\7+
Ff?�y6�m���V���=['��$�r�7I�?(9��x�� '0�����ʄ�K5ҷ�>p�[���B޴�HTY_)�r���GPM� ~޿��f��~�"�v �%���j�@
��P����r:�b��眓�*��h��	T�+���m^�5A
O�������L�A�լm�Ӯ��V+l�����O���3�L�g#�ϡ��EW�{����٠������,D,�E�����*���ŭ$9�,9��k�����Y	G�?�N$��6nF@�re^�TrV�ߚ_Z���>x�-�x�i�<q����:]--�ݳ���U2�'�?�>"��J��e7"�mWȔ�6Y�^����m��՛[&�P�;�����{���P��T�Y�gs! ���bd�[���^��^�i�.�0Զ����*�KzN�.�p��E{��v�+Z�n��|�C������<�w�}w]-E��L�r�=����e9�ҝ�9�ul>=�lvh��Y}�W`BP�4�f:(��$Xj��7Pd�l('��SV��*}�X�'�xV6� e�i���G0�����D�N�Ƽ�4v#7��S�w33���\��g4�ﱳ����s��Чù�9�F"e1Id�a̡�ߩP�9�|ͧV+�TY������M��R
�i�P,XPdR�xW�$'�W��D{`�.i��0Z0>���-�H�4��b����zP\��u������S7�O~�%!+>҃���3�+p
��0}��dȞ,�������}��ߴ��I^<�"x"�`�����
9�T*�u��V)8Ajk�j�ZΖ��u�����;A����F�T�gTqy�jR:S�H�W8a9�օ'"Y���5%؆*�fo6T�"���|�%��'�qF�%�#��bQޗ�'rY�t�
�YPͲ�"Qd,(*K�����;��R�-e.^��V�N��U�D�+��l����N�B�-���E΋���@���p�+��C�&����!By��Y��ǰ���S�mV�
��`%oUj$9,Q~a֟�l�������A�U����GK����@=[.nΖ��΂�!���Ol��W:I�SPN=ي�����x@4RlI�[X�E/�v��U�̤Vl2��K�|zv&z���k�e&}��7pX��kY�jٜe�-�n���Z�B�0�7�|��{��Fӂ-�5@���j�or������bkE��h�z�p[E����g���?���{gvxԶѠb������2yl��,ɽ�m�l	�R�� <4Z^n8%{x���bs�W"3l���`kp*�Z�F�#��ZY��w5/�5Ո�{̀���Os��B��;�83	���@@R]Jڿꇖ}�_�;�00\T��*8LRE��-��e]�=�V�{/h]U�����O���O�!��&�zK�-�]d�wy�( o�ê�W���#0&@tҔ��;�Y�\��c�G�T0�QD?� �=�L��&�q�z恨�A(����O D����g-*;,��q�>��� ?3�X.���瞲�|�Sb��:�ږ�U,93�$3$l}mx��*k>�'��!��׾m/޺b��/��-��9ۺ�'$�Ɏ� �Α�:Ѝ�����F�E�ʖ9[����?��?z�`�-s�h���60�m΍#��_�`,d	��o�����(�#���x0r�F(GZ�QHzB&F�ؠ�DD��q�=ͭ�7	W;;F�Xw���Re��UYs]��=Qt�T%̜'[P%\�Ua�7p�x 7�6G4Bl�q�'I�n���8��M�����b�Ϣ�K���
`��3�9�����+!�x����K��y����:ؖ��^y��͏Aj��_99<�7�v.����:+���[�p:�E��C4�7w����9�<>�D�ٿP�Nլ̭ɤ��M�gd�<	X�Q-��v�vje�N����D�g�H#T#�nGR�����c ��=k�l���p�h{HN���]��Ձg�o�����Ƈ�X�$�?��l�	&�S!!S��
~������CPf�l��sl�?e�~ˎ�{6��ûG��%W��C��ꎲ�ݝ���\���6#��&iiNEҴ����w��@��
��<r��+*�G�Q��xpd;;{��ǥړ�����	"�\�C����e��8�@�>��$]�w�U��K�P��@��^�M�T�|�O�h�~R�P���=�}3*UHH�&HMϭ�_��H�0z� 3_��H��MTD���UQ����;��q�9��!)�g�`�� H�� ����Dz���$�B�ѻ�Z���G��c�)*� j�=��H�B$�HrK,8cya-���	<�#���g��������5P�"�^҂��6S��(���d>���q��M�6�ܱO~�q�x�d�m��'iD�.�ٱ��� �����z��f�*�5�f��Y)�dcٶ�kb#/sy����lǋ�z����� �$[F�$.�DY(Δt����+Hg�ܔDG6adB�hs]s=F^Z��!�t���G���6�=C+�k��){$�/��1Ҙ8/��BV�/����R�'�ɮȞ<6��C���VhNR�ڄ�Q`��К�n��<o$�R�Ӽ{HW�:����8�I3>���i�s`/X9_�w�M��"�`d���b��_y�����Z�2���>M:OlÙ����額;���L
J�EE������\�v)H��z^y����y�H�T�Y@�=6��:�+S�1��i�@N�`pz|b���JŹ��U��g,���Y������aϦӊ]ػl;��m5r����/�o?��|�'�XTl0^Ʉ(B�M$�yI�k�@0����n�.Ҥ���/|�g��T��^�/��g�����Ά6����Y�;E�4_���3^�ۖ�~�b��|	x�*�˗�Z�ݳ�|���:��[vݳ-�,�%(���l�pxh�yך[Y{�OY1�����T9t�9��$X��<�?،.l�p�y��`˦�p�U�a���$\v/Gp"��<.`&e勥��IG���B�F�uD*��vD�����xD����\bL&B��z�N�
(4޻��Qlr�&`_HC�QQ�j}F�M5"�->gf����d����� �b�,c��ق ��� �J)���d���I{��2���c���N�e����u6f�\L��@��3����?c�ۍT�;�N�&�R�r�����m�'f���=!���Znvd���M۾��?�ӿ�`;��h��X�1��1�t�W�1�Қ������YcܼR,Xs��m�2Œ=:���^�m�іͬ�e�O`�'Q���l�wR�D14�z��?��
�DFk���FN�6X��F�5q
t��JF�M�_�iU��³V�@�⚞��4��VCҤV.FJ�D$q��uOq�3潎��%g���V�c��Ո#��7�7�m�OEZ��۰	'��P2Ȥ����EG H�G�Ȑ�Re+"W���-�����S��O�֛�?ǯ_(���l����h�~u������uzx�.��΀(�g���WbJ�:��?P�{u���$/O��F0ܬ9����G�dZ<���*��|h���(8��0�,���Y��T�����.^��+/>��Y�T��m?|���pܱ��+�,m{+o{�V,9	���{���m6/Zo8�r�d���&Ӿ�>9�=ࢃ�g�FV?�WK���j����l��-f�v������i�}m!����ڝ� Q��}�	׮^���-�taWD(Fo���AW�\[��i۾�Ϳ�~�oFl�-+�Ի"�p8�g=���2}���S{���ը���#m��ɘ���p��7�`9'�8d�^�<px�J/�: &����zpR��8���
j���x
	���S��Y��6�����lyX�av>�a�����uR?�{�^�a�$���"jC>CK0`�+UA�$��u��咍�r[��7���u��σx����%�K��""Zp^���4R�a�DyŢ'-��l�Ȑa�tڶ��a��I�� 	����5"ؾ��O��VC���a-x��{0e�@�^���E->'{���<󬝝<����~���[cwi�����5�K��X�~����H`��} ��3xn͆��5�ڌ�3�Ƞ�+U[�l�k\b��G���jQ2��E�umm�����h;�ƥ@��	��rYc8�ra(*vn��"�7��L�)��>l�o'�ƚӍ����u7� A `l��^�Yߥ�E9����V"��׮�b){k3z���)�&��A����?�C�9��B�p��G�"%>�?�?�)֪
�Td��$�x|���p���^��-�E-���O��"0�ǋ �`{�ï�'�_����j-����ye�EV"ܯL��<��[���"娠����dt�SC%���d>�)
7S<pS���:����4�d4�j)g���F#)0y�+/]�$f�ȡ=���}����dֵz�i����޷�cf�v�RnZ����5�6��dC����Gv��r�X�0���y�ơ�@;N79US���һXT���0�p	>� ,X&3�W^�b��+��O�yώN��lܰ;w���*؆v/=&�N��t���*����D׶R�k�0c����X�!#��;V,�X�@��Nkn�'V)S}���37�ۅ�;vvr�ୂ�E�����v�+.X�J�:�J�
�C@���N��O=Rشk�X2Q�n���E6.�.Vl>��~�bS��@Y��J�иKb�9Ni��gF�H�F��Z=�N��8Tc,	�
G3����x�)�H��`�.l�6�Wū*6��RHj��J0��BA��=f$��Db�p����v���<QI���.��ʥ��n���c��'� ͈�3�<c/���Z.�J���O����Ѡo�N[���Lz���^<��svzxǦ����_�e��?�������Z�L(�e�x�z� D�f[y�UWV.έZXY���E����n�XmhΖ�v8۳e~��٬`X�&�ک��.�O��u��qi� g*k��Q2�� �ڮ��		��Y$=T����O��j���^[������XFI��ֶ�Iz�h$S�p>�,�R1�	Y�gރ���8�$y�����}�j
R����M
(����!�#�D���xl�E �Hh��8|��P�K�ت#T$B�}JX�XQ�w���s�{�mۮ����'���d�:w�{��_�����E���Ӷuzl���&Y�3�M%P!�KzםU�bh�B�uiC
^�X��df��26� ���M����1�Q�,�Z�p�����8����q�A|1]J"ϖ3��*Y������b�;x���������};>���$�V(Y�^��+lK\Tx��p���b&�F|��Y'����C��Hp	)ewS�m�L.`�bab�ܺ`_���ۻܳ{�Vo>f���aK}%Rz�X,h�h�ٻxUd�~�1���&l�m{�w�o��r�=b���lZ��4����ss U9�M���涻]��;>������h(�P�Rj1fX���(6B�A�	S��n��k4h9Ӻ!��=s=#����\�GE����*V��TEG�{ ^���R�Y��1_;2��z�:\R*�u��601��4�7��8�^>�*PQRy@���� @y��J7 Ii\J9��v��"�[:�J�}>l��S.^�믠�;�.�t�X��Z�"q��3�}��:���Ǔ������3� �I�1���!�8��14ر:XAR�l�I���=c�ᙵ�~j��³v����?���}on�p=h����Bx��Hg��E��ӊ�V�2NE6��VU���l����Go�`�k�eY~�c��Y� �eqFH�0G����u��s4���@=Ҥ	�+�=`�VYr� GU�W$*B0R0������T̎RQR�ˮ��d�~�իW����p�2�ŵ&�ܜ�� )�jZ�ީ��D1�~���j�$A*z�alA��vm������B(��dA-�X{)G��
Uh��E��^��+Hye�	�:���
.H�mc�X�FͶjuۭ5�r�ŏg�m���g��7���;��Y����'9�LQ�qat�r�'����`'`���+��`��ߛ�'n6?�8lۈ�,�߃���C	��wxHљ|e�u�WE��m�p��(Ӟ�j=�`���l��z=2:��N`iԪV�1I���p +�-cw�� x�?����Ön�N����H��_+K�4��M��k���U�n��\,_�w޹o��d���$� �ԕ+�lo��m�]����|�f��̬X*��۷���߷A������`��-_��(�j�U�V2��/�=Cv���o4j������8+;��x��?�����O� }��
Z�j$��a%��������L����w�Z��Z�>|����<V���*������POwcH_�/���!/���p��O(��6䁜�����%}.�Ъb�L�|䳽��+eEu�x�8�:mUҳ�lO��d!��㚭{�I�k�����R�Z����I�k&�D,�J���v��M��n&x����4�Rg�ReQݒ������\�#lf�x�9N�}����nڍ�.ڟ�v�ݹ�:���Ҩl��DT[���Z���3�X1���-��1g���������~��}� U��zN&P�BH��yVf���r�k�g��
4�E,\8EP��X���%��D
�$�Q������y���bһEj��Ju)��&��/_��`K'�#���;!*ؤY���s��h|m��0��H�xz�J�  �^���<6�ɑ K)0���/N�N�H
��gҾ���Y�g7=! +�O��D��qA�B�N(M"\�<Rx`R��$hA���E�ݩ6��­'?��m����m4m���eK��)z�4���J�]3�@��I/vI�q���g�����jex���CF�̩%�A杤�"#�4+�+����.�L�02X���[��סU�XV6w�^U��m�vm�t�)X)e�R��iUT{���l:�rf�W[�=$�r�J��d����!�{$�Ƥ �,V��ˬ:��/<a���/(�޾wj���}��#k��ww.b�K�_������֎2���Gm�8���Lʕ���ӷ��?��MF��8��,�+'#y:�=[����t��/��p��v��%��`�a��Y/��"�%}SH-!���ȃ�g��3����+Y�9��=	ED��6�~2R�Ҏ ��׉@���Qo+��l�>��Mx�{�^1o̨��Ɩԃy�$�ϓcp�Yt<;�8�`/'��{|��É�Z�쉨ڣ2�ʛ�3t|>���8��D��DTR������N�Q(�������|�){���P��v�u��I��n�"����
��4��X�{�����p���W����l_��w��{{�?�ш(��N.�i<�SG��t@B�RC�Ń-޸�f�bEt�wjV�V���;ڲѼ��V��le9�|��eg�?�~%q+W��m�4T\���V-0A\\�N��휏{;XU[�8%��    IDATlK�U�%�U�K�O�%1�i�PP���u���x��'jeŽ'Ъ���j���K�3�K *`БXo�I&��	n"'�=I$��oP����3%^��~�}�׈��=������O�A����m���C�w�/������������!�R��ʭ?������8���U[7��xb�mD*�ƫ[�՗	<�s�2�h�t�px!���Zmv$�Y��q�*
OGƀt�7zk�}��,ln(��Tl,$�4'��u;=����0i%d���Z��d�� >��<W��Q��� }c�]���[G6v]���,����1�p>�F�YJ�T�@��F�Ez���.:�3=��?�i���bo����'w-_ܳ�c\Z�]zI�!Q{��x��1�O����`��C0cS����{�	V�a�>t�ƪ�Kz�lRz����袸�ӿ�Y�b�sp2r�&w��M@���Nm ��F6�ڨ�7�+6�/2���|'�i�X���C�n��/��D�;���F�4���L[�fx�VP_x@ż	}yO��sw��s+�S|&���
�8f�Dx�α�-?$Aʟ�p���
e�G�4y� �1<�#I��Q��_z������ 2@Ϳ������a�J�� B���ޅ��l_}�U�t邳��: �R��x"�y���{��!	-\��=�\��O>i��[���=��{�ƞ}�kk>4;>f�-,_�ʏI�����Y	BT�����-����n����d�V��\����D�m���l'��%M(�"mW�"xl7���@�� �b�"��i.hj=[�v�^��QiCh?��B[��/�����I�zD%��iT�hl�;'�q0��p�ji�e��F2�I9�}��8��������z��H�%n��j"#�<��ZGIfQC\i*@�*dá3��>b�������{���>K�b������(9��}��RNe�%T�}Q��}�֋727m쇿�_�=�����MN�p��h`��xd�g�T�Rk��\n�ግQR�P.!Hq� ��L�������9�������b�2�;�()��.�I�Z�t.ъA�%e��<n.vQr�(����O�E�Hv�bG����C���2<@�YF�lR*�P(*�0R�p/�Вʑ^g��حtyO���~�מ��k_��~����OX�~��������߶jK�����]�v�._�*&2��p�U`b�i�n�siw�ܱ�wokJ� �̹���[)�z��1��=��9ؚ�g�"D���A�z�X���$����r�����5Â��lV�Q�������rBVW�"h+���N�Mil(��h
�M�ʂ�8�\6�\�蟁���2k��S��8\b'��97__-��ٕ�&�/�-�1l7�_��I,�H`�q��`�����*����r�rh1����>�Ip>��W/ۭ[���Wo:�PR��nL�dڳvK}�`�:�=���7�.��>�'onٕkM����5ۿC�.*آ����m.�d#�+I!�6���uIƂ�/^�+�;��y+T*
���#��bY�[��l�t�}π@�l�L��sOAJ���D��(�2��� ���a�,�y}!B�^��YP����R����g"۱��$%�	�T��	jgY�ӜF��4�`�N���c���V�y�3��E�S�T\<F���Ť�s�w$|$
��,��{64�#و ��\�כ��:�>J���Q�wmA����P>1�����*��^�ĭ'>��v�z��`t��t�R�;=���)�$��#�,� '����㹪\�@�����F0��9���S	��<�٨:$U����~tx��Y�geHh�p�NwwFq��@��[d#a.��.إ�%�L����?�N��j��1���GOփ�̚cZl�9�փ��Jy��݉G�O�����Vg�;��I���_�������3�o=f��[����B�� ���(ؒW�<����c���ޏLJ+o�����'?;[�8#T�9d��I����r��)к�'9�k�{�	�w��R�A Q|m��`��.�mT��9S��U&f��rT�#�ǡ�2�	H7`����A/�`=6!&PY�"�%�[��&�M�=�u KyT�!	���2`ۀqׯ�`<�;B����6�uV!��x�
h\�/�oSB���>:pI���f\S�����2SJ��4�! ��6�����r9���k|��k"�*XG
����H	x�p���x=�8	�O>��]�-۰��=�TӮ\�����؃;t{3�-�.�E&�R�so������lw;o[��5�̧.����+������[�T�䍖��g+�doep��ٺی��	��hp]�n�
�ĕ�bLAo;��]�����S�%��<>��TV-�'l�H����&�f�Tt�>��6�H�2yֆ\f��Ba��H�����ۙ} ��V�(��Ԏq��+\����IK��F�2놿�ِ	�u��M�@J�^��G9�"����LF��\�j�,�Q)+�
F�6�_��T������{��^ٮF�7���g�
z���E��,�\�|�]y�B�O�=�d'S�2�w�jV�����2��
���0�+��R��SE�(���)k��_b�֪e�P��T�}exP0	s�R��% 8땀K%G{֭zA����\��I��e@7@��3I::�B��#׏�K��M�b���D�K�Z�>f�����~�>i������o~���o��|��DCP��U?5��z�j;;{v��'4������Ml�����Oj�����slK�dZ����-�@Jc[NJq�6�g�n���M���g2�ؠ��4����ͪ�*A7ؾ��ϿR�!�,xe�i|���L�}Y��&6n(&�(�g��^Id�4���T#�J΀�O$i/'���^���d�W��*����ϣG����g�`{�5Hh�־�ㄈDB���Ä?#o���C�:��N������
iI��E���nؕ+W�`v��uL�tq��0��!G�%�!�$�Ik	~��]�ݭ��zwl�]o����P�*��uK,�at��F�,��
�%�8+�g�v�bE�{������,�.^�U϶�Y��?~`m�%2p���*ۜ��ng?���F��+���wiu�|G0DmGU���x�$^�� �|�S$J�����`��ኄ�Q�d�a]��T�,�����L�Tek�y���k����\��n��:z��z�Ȑ��l#*�H�z�N����y�D��G�k���h�Jv$� ��H	��;�oL�wh#'���Z�-0r�\��[$��>�`��<�YY��q�h�+Z�T�ח�5�lג� ��fC���Rd��d��H�p
��X3�s]єI�&t�r!��?�Q�H֭�9բ#��,D@�g+���y��m4�Eh �oѦ���j[V)"������w߳^�c�{M��Se��鰣��N�W�Ju$w�dF@�;����R�7	t�hE�~�7^�/��/����kv������Ö�ޣ!���1S�L��;�,�a2��z�J?�ʒEL�}��m���fX]�g��0V���+�))��JvX`��Ѭ�#7���=��&����L�f0��Q�� rN�ʋ����}S{bЯ��$��	G��4��0|�����9��Q�-�s^����Z��G
X��So��a���u�%�?>O�u �0և���g=gl��?�É�_�Pr����q����&�e�!8�A�;)�	����<	�3ͬnb�ƾ�^smw������U-����̴r8���eL({ѻ6�[��X����d_���;���۬�+Y��h]�m�|Q��°�(k����k�V��,�l�[-eD�wi������62�-0r�l#ز^8�Q_�0lS 	IN�(8a�t��DB�� �)9�0Q�����f�(78�Q�����$����n��A����U!�6`��s�
|��*8۵	A 9i+إћh��gդB�L���#�^���B$0��:r",_�o��#��ZF9J�<��qŉQ�ne�A*`d�Sm<z��[T�?Q>h����Z�;�VظE�v�vrJO��z���"�����n��X��K��aF6�t:��l"d��X���+"��Q`����Y��u�Zp�N'�nW\a�s�q"vc�?tj�*g�BM
8�h��2u�R���ۥ�<zt,����KV)׭���E�Df����l�4�Ch�)�������a$������^��L#�����������Z3+V.���-Ic* CH@x!O�v���6간3���Q���ټo������?���̴���tf�z�Ǘ�H�eNX�sl�|�GHE:���O��>Ġ$��_6�*�oI�8�Q[h�:r}���7k@M1��g��9�'^�����Q�T��Cʑ�'#�zP�U;st��Հ�t l@���UU��
���7�r���D�bIT2�^���U�f������A��҈�)�x%���60�g���j���.;�c�E�y��^�Y��U��y)IAлpyϫe�h�}�N�NG�����ؤ9�JX�g�wl4<���}��+��K���}��S[�M9�2�ĥ(I
��J��=��Z^X����?x�l���U�M�s�eo���F�f�-����}fl4�k^����,[�3�7@Z�i�FmͰ�Q�W=�#�>�ʍ��Fף���[19����]��Q�V�� u:�����(=�X�u"���S�ae�ceD��O��c=�\�
Ɠ�Wṃ�<J3����zžY��	78qFFu�8^�Ϧ�5�B�(��)��Q�y��(ʹ�b$�^c�� ��a��\�~�02�}�ot��,��bg���;>G�������"0.�L�, �	Y�o~W�X�׳��Ve�e�6�S�!�<���sF&s�􇏎��+Za�J�����g#�d���oc���F�x����|$դRaa�[%�~�f�B��ΔM�껖ɢ�۷ã-`���t� *iA㈓T^�������p�멪o��CD�L�LX���;/�o��?����w�����s�P0=�+���$� ��{A��^kj�˞�Ѩ��q���~�އ��9]�j���)��|<�2��$T���%��d��R2b0��ϗ���on�8hT�=�e�p���ܵՆ��:P���+`�Ș7�r�0C�{��}�zM�Б��s7�1A��"��{V�K#k�L
r�=�z���F�^UG��A�P:̸�
"���A&*��ێJ_�-cA����h����#~-��&�4Sc��Z�6�%����7n��������!�	ctz=�Zp�l��O��$&�._�բg����ŗ�٧>������}�?�ˈ`:AH��Dv1��"�e3V�Q�ac8�Ra�Q z���V�y������FF�b�k؈���(�ȠPH��%�Xfm��ו`J�"��_Eb
r��õ�FKDgEJ�6!�8�)Ur�9��m��9����IIP&'�To4^�F %���TǺV�9[F!C�����s�ƺu$$�?�����0��7�Xk�}�3�XS�Ұ�"��ux|����^�����y3��T�I������`�9��W�ã��{��4���7�v���iuu�o5��Rv�voر�l��2�f��y2<h�>8��a�s 㱬��)N���l3r���Z\�:f�3k�;��-Z~���0�m��K�Q]W�T�3���c97�H糡��Y{��5��W�F���%�ە�/ٽ����P�V0[6�C���r䉓 `�q����ɉ�N��5K��`bvS�󂫎�W�����oپ���4�3_����퍍�"�7�O�V����v��%�5��k咕�%��;�l��4j?x���B�Eչ\��`�'��-\e��RI�%�Y����m"��W�-k2���D��1	�c^6��f;�w�ԝ�����w�ff�բ��Kso��(-��1�U��{��\��ѯ�k�y?�Y�a��D��B2�^n�A&��"��w#�����!?�	Iǵ��C���@���`=���Q�ǡHG����E<7�(D-���^��]��$ؒ@��#'H.j��HRСF�+ނx��ǭT����[�����?�˯۷�u��H����l��U��b~���G����WV֬a�9�Jɬ\Z�ҩՋ
��b�Gb#G����`��y���{���6� ޻���WC�=��#=N0���A�
GpX�|��պ/�:Qe�y�G��Lĥ�ϱ�&��uD��{�[�K�/U�!�ļ *�g����\ģ���.)�${3�r��{W0sI�����:��5����N�^Y�I�;�E���6ׄ��-9�ە��n=}%������`�:��[�e�� �L���,�Js�+�<<��pj�,�U�%˗���mnC[,GR&���V)l2���i�n��7��5�L�&8W��T��(;(f_�9��FîF��*s����9�H�%�2���5
@
z����.�ј�/m0�`����g��Y��O�!�+����b���`_']Z�/��ac��S�nf|2S_���������_�o~���o�e��>8�Vg�`�C�er�Z���.J&�B��R�R���ٱ��m�5궿�o��޷����#R�����wEbZ%��P��N����Б�s@��ҁ�س1�ϴi�*H�Q��I�#�eH>4;�������p2�+ض��R�oR��+�~�s���A(i�F`T��F9>l���DB�M��_M=ڀ�";"�D��DD�)X��)��рK���$'���' ���� =���3F�/��	���$�����.�H������]�7~�OFV��NT=�F�����ao1�R\X��={�ً��7������{�޷�aӉ�.3T�3+P8�kr�( q��iT�l��i�`[�l��#O��l�o�fp1�)MM0c{n�N:�\w�	k@3�)�ֵM���$���,jT�Z)IO����9������]��V�`ez�\ͦڛ<?A�X�H�J+Y	O�2&�����ґ���KK�I5��H����Er%�֫'���/�$�������������	�o����Q%�'�l�hg���S%�H&��rTbmla#k��<�����l?~����[���A�4)�h���-�9+�J�-���<9l[�����=}6�p�X���Ҳ�ѠC�9Z������f24�Jեls���y�Q��� �1F�SI4.�VdF�p )ʵD�2���Z����z_�&�Ž=�T����ӴF%�q愻��G�|'�j��h��߼6�FHc:S@�X�a�h!�"�h�����%���G��/����_���?�Y��k�{v��F���M)恷�H&�2�D�-��v�:�n�k���F0��۽����xBSTo���є�6��H�'A�Q��ro�G��؜mȹ��)����z6י��s`	�\xo5L"h�&1�5��^s���A�8_�0UT$*+@'���|�S�B久L�yY�W|�P�Y��#�l�F9t�(��k3	�j|z�I�%����*A�h�"Z'I��4z�:���-�'w���K����3�և_�ܢ������#y��U�"%N�B~�mr<B��F��,��lbׯ^�Bvb��=��%{���7�o���Y�p��3`޹�i%��A�K��X��|f�V��l���C���z�����:�f��Fe�lWF/�>�(�Ě��A.��R�$D��1rNx`)W�tA&,��>#Ye���+e��:�O$� Q�F�¦rL[*U��'�.���`K���fo)ˣ��g�\H*R��Y�m�!�5�u���v"�z��na0�e P*�/k?t$,q׬��^G�`@;��2����ȩgQv����vw��+W�|�*��ß��:��w�-W�N�vt�Q�)款-��Z#��6���u<�I@^��*լ�T�<d��ee������=:��Y��I�hV���
6�b��L�}yV^�kZ�Q��j(8�n    IDATn�։ժ>����=-����PV���� �����m�0H�-���#�N��2�����C`;�����P�2����;I�1G6Y��c����`_���տ��=xԵJ튵Z;:�h�`����-}�����.r
�'`k���c;:8Qe�:j�l
���f@#0���[JHHL���D2�<%}�f�މ�5�y�6Pl^�6.��u6���4�L�X$�t�Gp���G��7�B(H�\�6���Ħ%Y����8Tx\T����U-p�f��^�_P
�FFε�]T�q8�w��Z�:z�8�f5�%��p$$|�P���5+6����.ir+����ꩴ���G(��YY��̛O=�q�K����I�h�Wط=L�|n|&`}���+�,��|r`��z�n<�g��_�+{���V�^�芤=1-Y��1[ %�go��}�!��[����fѫ�j~l5g�����vY�� �1t#�iq�:0��Q"�i���ɍ��t�`�}.�]*�������F���'���W�bk)*E��$����.H�������[�"��h�f���SA��$S)�ʍ�:�m$����Jӥ#���P���Ík� *��ss��
�I/@~�I�QD�jM�Ý�r�����h�V�v�ĵǞ���i�e�s���������m��Lr�i�����ܚ{%���6�m2��0D�6�����m��.�Vo�c	xi%ڠ@�㕝vv��Igdg��ʳ\Q6~(")�M1[�������e[��<�Z��4��.\�S ���"&02Cp%��F�C%��v��{�:]#�џj�*M��0Yb�vEc����Ŋ<�FcP`2Y���h��D1��|�%�Wev˶����엿�)��_��=h[�~U~��GT��<ز�Պ��y_����+A&����&T��zvvڶ�IONE��W)d�ʕK���v�����|+�[�<�e��lÄ���k�F������O�	M���=*j~�I`��a��Q����uhs�b�5G�B���x���~����1ؚ��s[�A/z`�k�`D�8�t!&vz�>��*���B
HC�� Չ���S#U�X���!b#IQ1D�)sUo��M�!� y:��%�Į�������uϞz�i�E>nAT�x*[�m��*ZF��Ү=�����k�Y���]�����o���������ک���4��^2��Z��%� YŌ���m�kDA�V�*�bD��T�T���k?�/62���V�?$����0�����1N}�f���
7�6�sor�����ծ�ߘ����>��r"�2fw�V��������/�ҨKRR1�5��عc[��_��T��L#�	�i1����hڡ쭤D�����϶Eb=�"�F�\B�:��<�����Yμ�`���q� #�~�5�}k"�lC�"*ۭr����?���u�s���~�����/�~��o5��ǌ�Y�2���7S�u#���<(� B],[�PR��t��9�R�ʎApAt3�5i%�>��mw��O�*Tl���8�A�@e�����׊��U��p�9���kiF�,5H�?��h��A���J�cziy��R)���f6���C)d�dS��&ػL�*�<D!�Du- @gȲ�S8?���ǿd_��쯿���m�z�:ݹ��ŀ���d�d�[��.�����l>+ry:��t4�Ng`3���w�c��̃� :�8�w��t�h��9xe��d肙���,)��VT�1��X�b�1.��;�x?ڙ��0sT�����t����mR|"ea��i4!*M�%x.�^
�i�gS�BզQ;���C[�3���#ٹ�N�8�p��,k�+��
yN>��O].� 1MU� D��o�Q�=!���<�4) QY:k�Rkፔ,�E�fl��T����*?*�p�}�'Hm1����O
��]*&�ܳG��s��q_�R���d.��eWC;x���?�m�������{V,\�^?�ZH�I����3�V���Z]Z!?�62$*��v�V����;:IԂ�m��kc�ir@��g�<�j��Q�=�l#Iad) X��`DNWħ�{ ��gL���ֲ>#�r.K�m"ݗi�3�o��'z��#1U+g�2�-�%$`,��'���y�pY�<��
bi-�|��$�n�}�w��( &R{;�z��87���Y�����x_�F\k��1$�T'"uK�9U�0��g�U��o>q�F�q���ggo���{�����]�t�V��(k����a�@9u� �|{6���m�a˚M'=:u���g���$���U,Kv_�[4����Pҏ�m��[�<0x�#z�(ݣ5<���
���Ԅ��+wB�E�L��x���4�"IQE0��h�@���0YX��0ˠ�ڵ�d)��N&H�$�F
2皰�YJ�0ز�m��k?��h8H�#+��O��W�s���}�[g�6j��=<�^�Ì>��&x��v�1���!����h]e+��`y�͆]�>d���琏Ô��j�����d�׎`+����O�������D!CNp��:�e�6�R�IM
�MN�e���s��\�
@ٌ����`SN ��t��*%���L�@��T�D��=v�8x�3��<���<D��	I������S�Viu�3�H?v<k����	q�*���p{��@��C�:)Z-�HO6+r�� 2~oQn��'�����5�<Tf1j�k�fByM�3�|�w����	�W�������ף'$g|�H�"�⵸�E�	�C�J��}�>��v��=���忶�~w�J�+��
 \oTҀ��8��ʏ[��,X��d�jުż��b޹�T�=<����MW{6����eq#�έ���f���g����i�3��@����E�c$J	D����賒���$W�����z�iD�׉�DO�U0�	<�0cOG
����B�c] ���Ґ�G�\���k��O�v����AL{0A��(�C1J\�!Grf����k�k���@�����Vv�%���E�Vs����-���$�k�-��g�Y.[�T�f�a�J�v��c/����w�cl�����o�h6<���-��/�xV�G����Yf5�m�免�};9jiCoU)�����3�Vk`�A�f˜Fsc�m�U�H���z��Ck����y䲡�?v5]H��C��*Z�s*#�u#��� �8�s�8��*����_��Ҹ�P��b�q6W�\��Ճm;<�Y�?���D�SU˜s8�,%QA�r��M�ĺz¹'A�0c5�A�z:�rqd��{��W?y˾�7���߶�X�7֘�\�sm��m����yl�r��=��	��g,t'�����G�\��a����We�B��k������U�'k�;\vz�/r�s�9F6H>^1�!�Y�g�C�P�V�����X�/��q?ct�0���H)��R�y@� 3�af����{T���Ò��u�-��`KdM�R��]eIa*}���n��ҐL����M�Lt2��qۋ>'��WoԳL>k�^��ݦ�1�����fpp1	��B��HB�G�|�V��4��a�T]p�2uo�lC����^Y��|����s�n�V�}����K�=Z0��O�
$i�WG��kM����$�m�s�S{�����=����k�;0���'-�G���]�ŘAȬ\�$U*0���V�b���5����^�-s�-SrQ��W�0q��d9��~ib������& /��x� �\��O#���JOIS(��^(�K������I�'��r�uQ���ɏ��5EƓ�+qb߈���	����EX��I�$KΗ���4�@�BAA�N�+PQO&9��xE��/N�QB� u~�kI������:&ؒ`����JY�Iu����<��`[��[��Z���˗_���s�cl~����;ov��X�T��nX��cO���E��KV�`?��ao`���U�Z�����9�{3�s�OZm;>��lU��h*Y��֮�i�h�&*�?Aىe@���S,��RK�]��p\�;,)׎FUL6��m����[��s���gi6X�P�bDne�R�2��=z8a��h��1M�XH�3ym0D$l!c�zI���"��Fb擸�D�lj�����?���������C��l�޿�o��T#=h��ۆmo���K{
�
b��QƆ�a�j��#P���-I�E�@�� Tơ�����%4��)�P���%��{���K��[v��J�V� `7��\z����:��p�oF���V��Z�!Y����H~	�~6�&k3��xo�C�t���m�] )�e#�F3U�T|��Ҝe*J�\^���HpcA��H���kN�`+F)s��E�n��L2�B9NH�a[��tX U�s$�
��0�t��a���HGT�A.8�-©*��J"��ȈX MI������<M�G��cBӸ{���x뒂���?Q��/�l����F��C��(�o�*�Kc��EDƉ�����U��\o������[��
W-Wڵ�rn�9f�����E�H(���'�m�-#�F%���`��$�`-!Eg�W���u�g���E��	9g�I[��`�Xg�H��=�D%�5X�\74���ϽJl(|za7�`+Q�lA��
J=i�	�@p�#�V�d'�J �kWUn̴��0ж��4�D�f�T����9ZO*�:s=���� �?S��6��/_~�cl��u��[�vۗ��u�Ά9{��6�$Q�sY���{�ﴬ�yd{۰R�V.�d�>/����Yg`gݡ��]-�Zs�z��9�2w^ffR�b�#��Ř����W�V� ;T���EhC�@��cBP-�ߝHN�z1C�6$��3��.+i0ͅd:����N[s��2c8� �R;�B��T�.���:*4�����BD��esU�������w�g��~���P�j؝�G����Oa#;a�Q�r�$򘵲��RU�y�t����
�Q7�$<N���<h�!�&����D����'&�� 3'y�蕽�c��x��~�'�n[���l���`�=B��A
_��R)U�^͞�p�����6��$�F��$'�ȩ�r�A8�u���0����8<'x~-�l!�������#��vꛉ�{1�R��dCz#?��PřX��Aߡ΢'Kwb$a����H�R���U���۝���8�T1'���u�$#	υ����ɱ��?����P=l,&�p�c@��Z�/>A�Ǯl���׽�}��������G�Zn����P*�r����9"5Y��8�`����-�d�(Y��V�J՜�Je{pж��os�l�\�`a�����պ�;6%�鐗^ 2�3��EJS�y�tk�E���	���t> }��nC�+f���@ ��@T+=�`�}�>�z7���_���p@c����3';���'�g�-��`�uS�6	p���r�kz��[7ӱ�����XS��MÃ(Z�ټ#"�b� ��Ԋ�� ����>��$a
��8�`{��Տg���ty�����C	�#�W߹l���?�����
%��̩��e�����;����?cU���(��V�8Y�^wh'xa�[6]�����j�y�f���FV�-�����{eM��]�\u�;ߞ��m��`I�%KF")�iɒb$�؉d�%GS�%��$��$�%��"�T$��Hv7�M�po���p�=c��֔��~vU5#�L+h���3U���>{��^ko�jwa�-�0��ǡ6��l70�����&c��M`(l�-%�H�n֑�4�۩[�S�Q6����f��7���s�%f
ޣUPY ���V�J)2�8I�ɨ3y��*�p�a��L4[�<���W?g�l�𚝞aN߰���4�G�1[F��ӊÄT�Tl�<���G/I�x���`�C'�G�����`�v������ܗ�Q8/A�����1R�|T�a0��|=,��l�(��
!�4	m3��RO*nNs�!�3�&J>��"��`ȿ��i�ܝ�V?G&�i��?�̩��nH���d�ƈJ��O'vrT۱A�z\�R��V�
�(р��a�HXV( �	�]R�ZWG��~��P��g+�����$k� � #�%����h"Yн]{���~Xg>*o�-����`��<�����#��F�:t��/_h���/�g?��=��y�g�ۿ�o��#+��4=���b,�8�-���T�l���r%�F�ի�흖U[e�.�v��k�n<���M�w��:=�yΦK7��a�����]P(Zˉ����fzV=Ȅ@ĹE"H�\�i��V7���0�9������\)���%�)��2�'�&R�z��WC�݉�����@�@�;�w�Ԟ�ڳk���z�
��Q�1=3�&l%>���F{G���j��g�ו5���D���@OR������*yg�ZS2���e��VQe+��\��vgt���O\��zo������;y��[��Ɨ�M�v��C��ܲb������`�bæ�:���7�V+��<���LZ���{b��+�{x�����<��`R���`��m8Om>Zn9�FynO]޶g��X�&6���/+�F����"#c�s�T�R�c4�3�e����^@�B�l юnoi�aNU����c��E�=�u	X��ٴ�lyx�Ն�*�����K��{����l��G߶�.��=�?uQ��Ƕ^m��]����!i`��s��7�P�`��B1�Jl�g=�pCI��i%������+��o�G��k>������g�3���V���X �	LE�@�<�S'��7��(�,�؀&W6i+G��*�=�P�	�d�As�a���A�F���6��(�3�^l2�<�G2��cҰ�7%A�����yR礍�jZ�('�Dr%-�ԛ�{a̠*�Q/ڒBT�
0�u���Z��P��K��!�s�=��ӫ�?�ix�d�öڝU���٬r�]�{0^�����v��a�����#/�����?�_}d���Sr+6���$�0�B),��m��e�l����e�dRa��;��ݛ�6[�)ؖjU��s�s�y�tb�u3����HP �J��j2O��<�[ +1GkT�1;/��M��ֳ�\��-׸��v��zDE�sϊ�aJF��AB�x��ܚ�k���K��N��T���d-jK���D�rB��l�zX�W{O0�Ն�{2���)���ؓJO]�7�f�hPa�(V(�j*bp *e]��[
.��V��SO=w���������{���{���o��n}
���R�*[6�7�;jX6�Z�p��JQ�i��PD&��l�������?h���j(X&����ڵw������9�,6+8�o9'`ά����Ŗ=���U
�-3*ޅ=|��1���Y�q�j�4�gC�2#���,����3mJ̱!�8��E��&�dw!�!�ͨ�]�&4}b�D��a��'!z��6;�Y�lCI�^(�>�����1���}p�b��g)f��L��N��>;8/z�QQ��iĊ���2���ӻ�<���5���o|CU���)`G`����{��j3z�|&����D J�t�E�I�9܏4J �n��Q.U+3Ozb+�Sa�kK0�I�.�sUis
X=6����,T��8�X��d>6���6���<	�ʧ� O��}���������b$�Z��mD4�*�5T������{oA�M0"�')�-k���Ȭ5�%��Ǐl�$��-K�e#�u�u�i�ucm#�?�n���U�����}�+m>m��?n[2�ǳX��R�ǼW�%�F�����j��F&ؾ�ޱM�6���k����L�a#1j8�z�p���)4b��mh{����=��O,ީ'��Spq-������(�9s�D	����m�oA�M�w���gU���B�N��$$��sy(��� f���K�.�IDOJ�3�M@�Ţ'Y��'�b��D��f�     IDATȀ��8Z�J@Α��=	kK�3#���ν��)JA���\*	� ��l;[��O>���f�ч2�޼�;�����?W��HD�T�f�ʮ��e����l3�ws9�j�m���쇙��\�$��jan���X�T���{��{vwdGݜeV�!�	+2��ﲡL��fϪEg%ss	h@�Z�b��ڬj�H�̓��Ix9�!#K����d���I'�L1_����`s���;7��6��5���fK�֩!� ��|1�\�E<1�����h7�#���9�ti�>����h�[�62��wm�ܗ6y�����=�D@^���0��
S�c|()��Y9�[�R,;�����n�d���;��{���! nN��Fի�+�F�2����w�f��I��P-J#+�I��5�8,��l_7x@�c-�K����Ub�D'"ɐ2��g=_]��i��70O$�<�E��k-(l�3�~�]�;�Uީ����x�
��{���%*�D�3A�����1�4ju��ED����s�{H\��C@R�/��8��1��g��cZO8�p����"��k$(� ?�Ѱ��r<��-�3����rv���}���/ۿ���o�~c�&Y[֜��|�y/� !@޿�V�Wl6G'}n�vɶk6!�a2⒃yt��k��ڃ�]{�����-�b��cBΣ������j�dF9�|i=ǬsI}[�${Q�Eb�6��%KU����0\� <�g0�u�Hr4��=�l:[���=0�gӄ����a��~/�=�XWkQߛ ���v{��L��ua�璜�`+Y�j�ծȇU�N2�X�Ғ�.yK��>ap="�g����Q`9�8��v��ȋ��[*o��V�G/1bAU��l������]z≏�k4~(���7���0����l�X"���UsM[�/jh��m���W,�V�����li��@:0m��n����lo�c���Nz3{��#{��=:��dY�_���l@��rKk��V/ͭ^%��W�Y9���6{%�M�w{�?H�&��Ӊ>����P���󞘋� ���h�=����;�pFE�ʐ�l���'Ć��=^����3+��X�4�V}b��?�����=x8���l�'��rb��Z�Y}>�:B�@�Q���bz�ꫥBA6�� �T@��'yq�{�z��p�H��ݻ��J"6LxFT�H5F��/�|�r�'ʶO�O2�!��k�$C��͆S�JF/	�5�Ц�g��&�Uu��u���G�6��(���D��>^��x%���*?�ֽB^�a{���Kq�f.��"g!��둵oX�	{�R�^.n2�����5H�Q��� ���6٨��~��=XT��ц����y�&��
���`��fN �ܴ/d��c! x�ٓ
������?o�7����g�텗��|�K
��a�}�!��]n�V�i�<��jռ�m٘_X�U�B�D���5wv��~O0�`Ԓ����8yc�'��.�*�d����ӺJ�b�$ z>d�Y�?/�	�I�j�L���T���K���n���3ㄨ�A�:����ҳ��&�e�U�%���DK^�1�H�$�؂�+q�(6eJ�F3��>��֑nk�}3���c����IYi�K��&�}/��_�KR@�%���eʝ���tq��Y1�a4�J���l�M�zW�~��l����/M���ϣ�C���k6vYhڼ�g��$��,j���	�BJ���IW�S<-����j%�A6�Ѵ`7��;7ۃ����Uc���7y��"�p� �C+Yf�n=,��wl6�S��(-�%��n�bٲ��~�JE�� k��;�����q&I�֥j���F�TA�E���5z˱Ѱ1l�������w���v�����_���2�Kvt<�n+�-I�)!z+3O��3�F�-2�x�	�jz��`q�)Ң����� ƠZT��0s@ir�&<���T"��#k��+Ǩ����4��C�ޣ���FO&f��D�p�s1P%QJF��y�T�i����B�xR*����zČ�y����<U=�J"��˨X���]��&�\�;�f< I�b�]�cuX�+��D)�sm^���_�sT��BI�Bي �1�d����n>f�9��Ϗc�kR�>�=H+l�����`d�#F�X��N�^z�%��gvv��=�ܶ=��s�����%�H�e�^�2}pX�#�L�P)/�Y7k7��g�jeN���}}�j�Ζ���=�q������x
6&��oe����Q�t��D/��T���DTp�h���|Dk2��A@��Խo���1g����Ŕ$A:#�֬-��$o����$Z��K=���y*�ޫ"O����=���ʖ-�Eb*��C��c���)�}_ �z�#�����fR��Z=�����-�4����%k���`|ދ�$w���m'���h�Q8�,"�n5[���}�Žz������)=ۃ�_�[ó��7�޵���n�2�e�nKf�0{�n�rѶټd�oٱ�5Z��H`�<]��N��CY^�A[X9�y����Ɲ���h��-sq�1E��~�&����t$�w��Eт�Mg�7UHX����Ê�ۃ�x2���r6�$�62l�&����#ƒ����}<���#��H�y�@��%�[m�S�)�s�ٶZS�����v�\Ǿ��o����E;>��:��T�|�Wo���X�v�a��$֤���$��CK;z&����/4z�C��wj��v_����xV@�G6�$(�-�2���\6q���QA�Ҧ�%�k�����ί��s�4ʤ�x��N�e��̢*�<.�	��'�W`��4��+tؽ
_ ��
:0�	R=��$��d�QQ����%�]G/u\Re�x��Q��~�*+����*�R��T"�3�[���ͽ������O�KF���&�3�Y��k��3��w65�6Z��^���Z�VF�-ݷ�_ص�
�����p԰��g�y�-7�BH��
y���U+sAѥm+W�����T��j�{���ڻ�4-WٱZЬ�9��¦<����`�|'��s:�)S�o��
�T\I�궦j�u"�#l ޲�5�}DI�y�&���7VPi�J��l8^-S�%1�+����|��g���]��?H�Jb�j�(�V]�
n�W�yqR�)I����b,͟{�[�.Gc��>Ϛ��L��(<jU��L�`\�FC�h����{��Mk�ǢHJ��R�n5ZR�z�駟k�Z߃�����K	�''�}����o��Z6~l��D�?�bU�QՆ�-۹�Dl�^ɌG��ØDYd`���rE����N���KRq0Zw4�����;����ĺ̐�4��,�V�#-�Yq����*��U�Y1�V�>�L(�,����.���L�BȼUma̜��\J�8�L���{�D�R���qasTo,���$�/U"0LCC�4�1�45������o��ު��ѷ��ti�Q�����eyβ��NͲ�,l�[X1ɻ�2�F�����J��o>j"BF���HJ�3�L�^~W�0��YتV64Y��'7:��/�A�9N��y�B���ƈ,	�������`i�ȲU���/�^s��W�k�V� #��٤lP���4G}���X��J�yh�J!�,���1�("[�tD���W�
z
R f������7Ru�H@��JW��U�y���4���nx����*^z�I��,�.]^/��s5���I�`��ooTՑ����	)IoH�r������>����>��y��}�f7ߝ�hP��Ӂ�{P4�0z��*�.��[*�6K�U��Q�Պ'��Q��)y�v�Ў�U˕�l��I��l2_:�d���S�4[j�`4��#18�MW3�����������6�D�Z�V(�'�.Ѐ����V�	�(A��n�ϒHE��MS�kQ.����",����J~&�}�T�7H��3�������|���zt�J���[��h[E�����$x@"s��g�(��|2i���#�����l	�+���6r۝���sO<�l��>�P����۽��<uoW��c���U�]��;항�o�r�1��l���o|ӌhY����w# Yl\|l:�z�b����C;<��G'�/d�%V)4�	�q���fӱ��\���5�=HP�sV���g�!O�5���% ��MGsY뱙�8���U��
6�����Mlɲ� j��,$c�Է�������E=:�~R������~��޶:U��_��^�&Ӫ'������`;�;]?>��D͟{��n
�莦2��#K��a���g�X"̐�J64yY�"� o! /9�4����0C��R����>R@F��4�������?�&�1𳎫�(���v�WKlC�7�	�/*1U�	�c����'��T��Ca&�U9ɡ�s�֏���4��u,)�C�3�ov��x�� Y���u�z^�>���/�-A�TN� �j�'�; �P���A��֦���67|S�{J"ݜ�k��'����"����"��p�oI1K�<���_c�Zg��[�>�_�`��Ծ��W���f�n���˝�k������R�k�0g�:s�S��ђ��r)�V�ݩJ�������C��f�۹�`���p*�����ɥ�Qm�8%�f�	�Tĺ�I�U�g	���.���^̥/|_�á}�W���p�F��L'(��#㇜��$�=[��Lz��u�xP�{�I�b$�2_�8[jC]��T�^��"���S�'�H�A���F��a+VK�<��� �������K�s��h�T��j�c�>��DPc��}�s�T�(lm7ۈZ�>}��3J������·�۟Zd�-˺"9i�:v�-ذ׶y����r�e������.�Wt��sX�<�3m^@���(;<��{7�h��\�l���W�� :[N�¹���تp#}f��`�}��s���Y������1�ˈG��M,gk�+Nl������6#�X�<�tbh '6i2w}�}L�L����Ɋ���vN�j~�`�[����V�n���+
��e�F���b&�Ġ�HE�7�jH� D��R J����!_���?B�~m6^�[���(B�H���a�� +���!D
e�#�^��u���\���P?k���ɰU�W��kv3؋��(����C�~��J�R�f�Ǎ@�5��ڗT���{�Z'2v� ��L��}R�J�][6:�dB;9��ؚi�06#��o�������xp	��Q�6�]s�2��`I;�׋1�hYh��u�ds3����I�+�g�Y����s�"q��U��"#�x^j?>磊|*�����Xvf�?۱g�ٲBeb�|�M����h	�?:����
s�0gI�h1�c�'*ضEkT1#��Y�f�b�z�^{�={�^�F�]+��l��L�`=[�NF$��z!&�j���^i��iL�FP�*��O$���xL���W*s&!^�&��ܚ��
���WJp��t��&$�cW4c��o )k�_����汒(L Sj�e4��3�m)��ł3��~�3]�	��W��(�J�Y1�&Tg����;Y	&� 3�J@ӳ�ݤt�q< E�ݐ��J6�����Q�r$�t.z�����ɓ/>�����PV����/������5��hxh����fGg���,Wڵb�i���T1�% O�l�1#�	,`�`"�bk;w���ЎN�v��}
X� �E\�[6�?[T�T��SWwl���Z>�y�޴��X�:4�}w(��-m�l����:;3��Ͱa�'=��Pi��S�&9���h�i�z�����{���IU��g�.��^�"�7�l�������
���{fG'��;6/la���z]�!i)��X5(�hϬ�#�W�Ie)TfT�%X�& \f�bs�!ɋX�i�M��w0W�[�������;!̓�?����ಒ��	�h-ȷ��a����E �=DJ�{�?�Opu��;�z��/��2�YJ��7���H��>˴a�,;��x_�d����|!����q�;L�~�-Q�
Ip30h[���I���h�x�P?�����^+�yTȫi}?-��!4D)�{��!����49��C�P}$|�?�K���5��	� 0 ��z��*?�����~���պ�����7n�����(�26G��F��)\��Y{�d�&d��5�Ek��֪@��;�麽��M��+��)�f˜/0�и"JU'�qB���^��5*3�l3�M�8rn\���k�'q��1l��#. ���Fi��<)���EH�yo�ٳH�a�#��]򞩪Ŵ����2�&�8���x�&g.!�VB���K}o	�h�`��~��^��0|#�`��O�T�J�9������G�{2G<�y-I7ܟs�(RQ�%ըYd�����@��n�O?r��G���N>���d���;��ϳ1��}I��?�;>1��j�/nY��6j�E��.0B��)��TR��L�;�h��F�a�l6���3��&�����O��)o��@d�"�gnfO=�g�V�ZD��vv��w5���o��j�拜�I��t����j�I&��, ܉�����<q;�m(dV�kK.O��q�	������Hk��=�Z�lQ�B��v��k��9�ޮ�����m������p���u���C���q׳��*F-��q2Ip��3)�A[�35��~�ަ�5|4��o G�y�5�ে)	DU�=� �@ڏ�c/�\Ώkͦ�ۓޯ��6
�s:v��{TmM:9��v"���DkR�Qljlt@O{���:��ͅ�Z�$�OyXxj�t�1V���X���]$<�=��~�$ܵ$���5d��LlbU��|%� ;'���k�d�Q�8V~�[%Ӝg�V��L6x~WjV�T�PI(h�vDTHQ���Eʛ'�ձ91(�Z�@�.�2���x��؞y�n�Wl��[�oۍk�,��QW�8C+��*��M|d���o�]��^�
��UKk׊֬B�)Z��ܴk��ۍ;]�O[��n۔i�Q��Ζg���J� A�8�g�|&�\����Q�ds��T`�n	R$�HvG���2�r?�d�g�L���,*�7Wn��I�� 	�p<߄��漞ǜ^Ľ�3�>
�9�o�Db���L��������l�����8&HR<����/���vb�c%��;�?�Jٶ[M������c����c>��+u+�+B2��DL��Bf-L6�i�W\�X��E�L .X�R�V���.���z����y�C�g�A�{}�{t�V6~��pxh�bݎ��v������s�JՎ5�;R� 
@������&v2Xs��<�C0�9ΰ��X�i���#o��"�)��[ع�]<_����ڸ�[��M�{��r&�Xɱ�"���|�j�+�t��7�.V���i���
\s�����J���(�q�aN��v�=2e���#�_�~��Q�$o������'?oW/��O����W^�r骍26��U[�/�2������|�u6����!���xy8�� ��`��8Pj�g*$-� ���T��u�i�R��j�v�W6Ti�?=+g�'��x"��pT�꺲FԦ

�w���=`e�f����rQ�$l���X��qlb�&M`��R�0���S�j�8Y9�_�G-6{b���B��08_B��[��y0��5�^/�Fө�
�Ғs-[�]d�4��F���S��3IQ,�g	����g�0$���*��k��G�V�0b�)pDEIK���z�%N$|Zs�J=�RU�9ϛ^o�T�ְF�)v/��r9�v�l�Ϸ�T������*���v��]��6y��<�O�"� m#cᲰ���ꭹ�jE�D���������wg`�]{hk[��bg�6�X����Gc�T]����*�5���@9�x����4a'3�#��-���J�/���E�#G�[ίp�	H�,)O%�9�K��=���_���I��/�H�I�B�Q"�T�g#�ٓX�p�<z��ad�o�m$��;�zS����|ʜ����i�C��T�uq�YK�-�    IDAT���'����W.X�E��>��dn���?�b�%]�J�N��N�fY�j����EkX��hRS{B�4��l�M%qi�v~gw|i���/\����F�,����?���B6E;x_����٭{�2<�W�V�����K�D僠2����@O�;���lH��e��<z|f�B�Z� �~)�2#[�a~�hV-��T�+,�b�f�D�0�If�L��|U1��4�z���C6O�;6V0]���,Շ*"ppG�C�bU�p�\]
����Ԓ5&�5�h��^�o����'>vEf��Wm8h�o�έ;)��S	�y+Q9��E�01����;ҩ��x}s�AU�W��%[��I��9�a"�����Ksy<�d�>������P�����I"���*��'��׃�}gyS�F��o���%�+�A��C|��������C>�� b��Io7�4Uˆ�_RY%�`��rµ�$#¹G�W���"3ة≪��$�AM�'p@�>�58?7!G�֡<�7��q����Ծ@@3��:<�B%�g�,2^��^Uo����AЏf�Q�,��EH�2��`�5�0<=�L�L�I����
uT�V����<'�xz��v��v+V+l�5�j!�����}{�ݼuU{��p�gk�F�q%9N�^�Y���zcf���ꥼm�֨�bYZgk��{���}��}˖[V�f�70��$#T�$�����v�7, C�5*T�_9�'s{��@�H�6ѐ$�𹒥4S��x���% O$��{R䞰T��$�b�!������X���9$N�#x0B�6��"X2�Aŭc�MD��Ti�ľ�g^��ჵ�ǢF�="�"�ll��G.��KO_�NӘ�Yqn�gG6�r��pf��>��ӱ�;�ȷl��Ԗ�N�1����R�i�BM>��l�U�9k��Y�,ըcD����w�3.\}}3v}/��/e�'��������ߛϺ6�`8����vt6�����<L�m����5�%C@ �9z�Gݮ���+%'�� �l��h4��b�p,N�ި�� �a�f�[�Eπ�F�A�\j[�\�&;��͊��o�D�g��0T���xB��]03��sj>��WQEG�&�f�0sU�$��tqB����-�Y骚bM�~n�9�_����~䇞��oݴW_�n�\;�ɴn�E�2`�����ͦl�lzTD��3����}_�ydĉW�Y��y���ƻ�.�SO6���2i����u�( ��hC"���:�(F!��U�+[m�e��$��s��iS��= ΀;���HTű��#]���������'#���BU	}ĪWa���fLK�;�*[3}I�V�7)Uy#N�^���7ZJ@ $I�"�6!d*��+��D_4`y�˦��6n�����y*i�v�ё52*�'t��� �:+&>Ji6X,�ef�R�&��L'V+;�聇dk�DB󞥞ɴ�����OB�i�A�Q�L&"�fG��sԐ�U�jU.��^ն��_<T�Os��7o٭[e�f;���H��Ge[,"LC���
�Q64�d�֬m���%�ʹ��B}�޼~lߺ��f��Y�%����-��W�$J@��De{5���H!��.�p]B��J��ֆaE�)12FNB_��p��,�u��<!�NdCÿ|-?4�ӜsXF�����WO�CYJf���E{&�m)c%�� ���-^_|���LQ�����غ�إ�}�'쥧�-7��P'���زEE��*���m;eL�t���PP,D/��P�l�F������Tޚ�m]�.��V�e{��?�ĥ'������l��G�[�\{����G糾=>�ٻw�6^T�7��E������ٲNˮ��jlf��t��?��Űkg@�3�3�rp!^�(�$��u X@}�Y��X3���Tʌb<�{���+� *D|Ӡg���"�V�&�f@�Ǽ��*y)�67����O�BX;٘iS��Zb܅�����i=���h�f�nL���ڧ?yՎO��xj��r���
��#���xn�̉_d�[F����B�gT�)���6&w�A��|�Ϧ6şW���@x��nb�ݕ��(z�z�Te�|�O��F�,�Sa����KE\��
��>3Y���7����IN<�	*n�Xd�8!�B���5����GC�)X�|�D�;`4�x&"#���t��⵸&��k�r����Z߲V�hy��cZ�v@˼��Ʈ�F�Gbn3h1>��Ь�H���K��6���ٙ")���^0�^�y�ȗr��p_"��vѻcJ}p�x�Z���3��܇R�h��1K�.]��1.X�v���
����ŌE���v'����ح�5�ζm��L��i�Gu����C�� #�RF�`n�J�v:�2�,��j[��k��}`o�8�y�sۊU|�A<葻�+�{�y��ҕ4R�d@���8W�X�h,��S��ׯW����'�J�6dUيU�=��i�D�֎�^|V�㊊���pD+�,U���k���!�l���^
�NI����y<C�_�܃A}�8&}d�ut��)�a1?��\nُ~���JȈ��F�����t8�-;�N��wo۷�߶r�����T�֑q���3�Ʊ\���HZ9���+#�v�!�����~��KO�������o��;wn�O����ѩ]�}h�Y������A1�QP����v;u��jh>NRa���Ãǖ�UT�2���m�A4��:5A�Mn:��ɑ-�Sk�k��iX69��Z�M}4&�����#l��傊ȯ�`���N"�d3v��iGe;_��$�M�dM6'���aG��Q0r��	Vskֺ�+������vE(���;g�����L���U0�0t�����RI��!��Ռ`[�|��щ����4��,�p���(�T�s�����76"eʉ ���|3��@�T�U���ryD~N�=��\�� ��%%�b��˭Tk���M#�o��T"�QpIl�Hlb�6��@c~{���׋MD?cx>)�hsJ�G�N��B΂��LNL�q}e[R�1$�2;Α�-�BG	b��+�HW�-�����H�jA����416�6W6q���0vNX�\6w7�`��D<��i�8q����֮?��]�2�H�+�l:��t���US�B�rrz���\[��yvw��ē;��P�"��Y��)1~�߳o�r�޿U�ѨcG'��.7��[��D�`��N�f�:Vks�W��m�a"S�欁�sy۾�־���M�J]��$���Wu� �A�QٲFCv5�I��d$-�Q͊۰1��zNB�1����vz��R���&���������A��@��x�]�+�x�սO��0P f�VCjKD�)�����:���'�i�����H�{i���
�NP蓌��ʹ�=u�l?��/�Nsh�eO	�Ã[��7�s������q�g��yÎ��Y�������
�:]%+S������k�����lIu����?��K�`�?8�x��[���A�����}xl'����(��sd����U�W
K��u��j���"@���Ç��m8�T��w��e1=��Q=���?���0n5*
�˴BQo�+Vc�����<SU�e�dg "�Z����n_��B%�y�β6�<�0�d�_1%�0�:U���R�6�m���AED�l�����y���Y6Y�ÇT�M�w�v����XcF�r�$�d��#s��k4���Nsx|����:ؐ�;A�Q��[����?>Z��D������66��K����l�QS-�
����d����R�/�����ס�������C�9���6}mՃ��%��N
b��]ְ�D�=:U1�������=�I���ͺt����%R��� �Fn�^�X.����F�L�O�7�9`ŨL���`��	/�xԀ b���\T1�����Xޕ��9�����t�_�b�g���Q ΍g��TG��P�� �~�)S��3HO���_%W�U�f�ud2{�/P"�ȋϬ�.��.2�9�+(��V��ν����ݸJְn�.�8�K���-�5�,4T+�u�%k�8n��m��;�ƍc�΍G6Z6l�#Ѯ&w2�p̫{��u�z�I%���_��ҹ'>�������E}U����J���*!n8:���}B���7�=%�|�c�3jm$�$�ꥧ	~WJo�^��S�h��{3_=㔌��HN<�����z�A#تm ����USì�\�ȫ�Za���;f��>kۭ�e�C�w��ݼs`S���㾝�j�'?�qkv�v��#��+7l�똕�Y��blC�d_Сgc��UK�D��T�Ћ��t.����'/?��}e�	�z���������c;8��p2���5/�8YUwa����v��rm������<>�ÓSO)+�6��/�''/H����dؠd:�V�x'��w���lUm<�˩f��#؆ 7���£�BH�:86���C�IA,�'�
��s��D���d��ƭ�*A~+X(=�^8tHe�����g>�	;>�ogg]��M�h9���]�׬Zk�d�=od�l1��|"��l�����!N
Cab�����Q�"��Pǳ��0�±�|lK©=:��ב�G0�����Nl^Q�ש�ub>3����cW�L�t.�z3�x��6e^?`_fN�$�b�/����{�;5N|�?�
��DS�yg��&�ql�ke�y�ղ���xj�	��f.�Sp����D�d�G�k᠓���g�	^t9���5jx�:��w�6X	VIR�zA'�cH<�����n0�RaD.m�$$Pr16���c��ýzw�U�8� M�tu�@���f����m��`9+Ɉ�,DO xvim�Q��w�o�6U�������v��_߷��U�۰�؍��2�\�׹�jyk7qEBeQz��)I����VS�v�h؛��7���~�p7�l#���MlZ�߾r�j��]spF�u�5��'����� �Jk��$�����d4#�q]���^O�nZ��!�}��5��h�8�!��@[d���"�ߥ^�&����U�]��rˡݜ�J��;�Aք�ʔ�s��]����vi�l���ݺ}�n�;����깉��'��瞿�v���e;V,W�hVٶ	��^� �5z����z�:��+�.���<��|_��a�c��Ϋo��<<=�ó�z�G�=�M���Q�-�4jv~��
���Ʃ��D����w��{t�c:<���2�+�C� �xl�sa����gMr��ڪ���G�;뉀��,�����Uj��y��G�d�C�r��R��b�RU�|���~<P�R%��6[]�P����x #����)�;?�	�
Ҽ{����9�R�e���6�f����$Z�Fu>�i6�f�G�U鏸g�H]	��P� ?J���q1����� ��c!Q�\~e�F&��%��<cPEAfrpl�W���N5��T��5������Դ�YEH:@P��#��'I�A�X,i�����:�/U�:N�](Bl�ZM��זs|��yM�^�5��B�z$'�$H����S�-��ɰ�H��g�X�NΎ��jX�Yw�C��=U���\���9�`E�ec�9�k��ؿ`If�g�����n�����3����6���3�H0��P)����uI�8g*jm�02���~O�^"�U�-�s%:�z��^͘ 0����d�3�	֪�$��Y��Cq.�P,�ԇ�l�N'6���杞�����7*vzִ!�I6l�� �Ê^�So ȧ��.�4ɬ-U��N�ꭖ�U���C{��#��۶�׬�� p'E.�"��rέ�.���P 'ı~ث�;��9H`89J�5�|�=��l���-7���Je	���BJ���GeK����� P�������Hz�[��!SzO�gq���E�'�61r�aOb��-�$L���4���[O�L)U9�Y��
�=�d�T��Z����mO_������~�v��I�8����>��gmgo�^y�-����Vj>cխ����dC�_�^������V�5��iv4��p���Ͻ����}l��e�ڵw޿s���g����mo(�d`Ye?���ɉ�_j��Wʶ��c�JAY=�zgg={�w����H3�#P	=��`	��W��=d#=6�o;�r��
�i�<���26���˦����鄝��?:��Ebf�s��Ye=X.�MG�06%��W��^����ԫ����0U�G�˿������M�5��=���QO�i�<.7��ԯ�E87�;A�k[�4%S�.]����dx�d��z���5~����%���6J�|�ɬE�KUGvL��k�%���$'�gz����TWz<d%)�y�2T6/.��b���7��( �,)�uH�q�!'�d%>�1���r�qҋƄ@NR6.���ԍ�� =Ɂ�H�6�t,T�kC�\�Ԟ����y���I#֌�'s����;�V�9*�����-�|$��:�M$4�=�SJ8$&��Y���AJ��'�� VF���,蕖}#�.4��}��$;r��'y�����G��}
B(!5�[��P��[��3��I�n��׾vho�U��Ӧ�quG���}Jr6S�-��Ts�锬�`/�;U�jg{����u��׆����٭�#�X-�U�\�x��	=flc4�
]}�ZS{B��׎{ɚ��$�alM��I/=>������z-:šX�P�����Ǔ�~9_G!�$Pz��ю�3ޏ{����Hld��ȝi��v�5�ٽ���I&�v�Q;����)Tx�$}��) �֩U��M(Z�vxҷ�df��;�*�m���G�۶�~�%{����k��cY�-+��(���ﵛ�7Bnf֨���(J�ZU0Ix�vv��H�����O=���/�-'����_>>9��ǽ#;<;���c;�(Gә����2w���Jo�����zxri�V�r��ݺ��޼F��̪���B�P'A���1D��6!.�t4�iַ|�	��K�-��J���^��R���l4f5n������Y�7�nwh3�B�̰�r+5*���urR�IT��'���/^��*�.�����j?����l���e���T�$3������Њ����/����S��}X�XM�"�<�>��`�@� u�a^G"強o�k�e�M�W�Z6���G־��o*�f��a�"Hb<䚱�WU�*I�-��?".i�F�띎�Fy�`O�[V$nE,�%�5OE��������I�$�@�Q�3��'c��ԧK���))��w�!y�z��7W5��}��ZD�yo���:�P'ËV���	�k4��#T�"%K�.��Ӹ�C��.���F���}���n�ד�M ��*΢WT��͉S�l,�����B��5��9�lvb��4�������}�ώ�ڵ���[6T�{�돭��[���uN,�V;g4��$�Cɸ��4�Q_j����gg�����C{��Ȳe�W+���-ʫ��E��U��R�fO[pP���8�-WC�ƍ
6��N��	�!�%T#�d�a�x��9
�OV�(o븎;�Ʊ����N|:Ml���I����G�(R��c.������?�^�ӳ�D��Y��.E���n��:}.�+��9�`n�,W��'���{���:�}����?�)q ���u��ll5˕����jŊ *���m%v$��*������ٳV�e;[�~�٧�~��&ؾ��w���/��!Hu�?����N�lFe#҅o�A����2u3��gV���ZiZ�?��w�A[�W������ ��3te(������X~��\R�Y"�1B��ŧ�0Z6=���.b��I/�=<�bS��
SY�L0ɴ�� +�١��L���d@��n��#����>����~�����Ye7-g}+,��$>@
k;yiB2�%�@Y~l���^��]A%)81����\c��?��T1ͺ��%)0!���b���4�XՇ^o����$��u� �#%1ZD���Ge&q���H^�5p��*9I��l��d�ڬ�ڮ5�<��;[��<��q�5����8	3H���l��U>    IDAT�N��s�F��_����?@�T��znO�X�1o9�-�XU����J��9�mP�f�y/U�J�(�^�����Fl�u����?�l�5�2�
�7ߵ_+�Y�������3��
�Q˜:cYf�Y_�����r�����{#�ҟ��o7l0ڲ��$#5D�'V�a<�B���D���N�$��R~)_h��jQ�6�d\�W����LV��(s�T���/���<iT���bk#?����>�<��R��'ҡT����m������/���Y%k˥�c�d�f��hK"N&�\c�}3��^�6��t(	(�C��D�^J�8�3B&1gE���jR��H�u��p�˽��%G��M�|Q���%s�5+�v��];����Xy2�Fnd��h�����J���z׾����su[�q<*Zdk>�V�!�� ]��bŶ[{�ll����?�����}l������z��]S`���Nz=M�!Ȯ��c����K�:&�6�Ǝ?k��K'W!��+Y17_Z4R!GIe&(��x|�Q���T �l2V �T٩|N��n� Ŋ��~ C�i����-랍�rx`BN�o��@wB�V�Ez���o�!�\�?[-� ����~�s��/�����M'� &@ٿ�H�AG�PJi(逝���c�%W�&0O�CQ��RI�}��8t,�@ �;t��k�UJT�x���=b�_��C�2zUi�0W�����jP�L�P��ң��rWX���q�Z6�,�!�E�Zߗ�9{Ktm���הH�����5�2�4�D(m>���k�^q���uܣY���nx٢C�h\���*W�?����l�Wv�a�*Z�mT��B�2g��^+G��X����	2�t��"x�s6Ÿ�a����<hs�Φ=�Nl6?���`8��d7��W�|dﾻe�ٞ�K��'�D��Ւ5�@�s��'V�ϭ��Q�J�lg�i�[e+V��+��p`�������L�?�]r�MΊ˪8[�[a��*!��%U����-�
7�w�OʳD��ω*�d\_smT����vX _
�2���	d�E�|* T@陜�< �x��'���{��%�)�:{r���/���͜�'�%S�#�K%���(Sݢ@�XF���X�$~�ӶZ�}�*A�;�6X�_�X1�Ye>�O<S�����(������޸c���Kuiїq[��>nT�_���.��-�۶5j;v�⥿q���/����wo�}p��wN�������0���폼�ņ(�F�=,g�a�l�G+�.�FAR��+��<�7�Q����Or�`���4몺Ն3�=��j�<dш��֠��Jh8����в�S�2�k7�v��%�v��=t����QM�zs�[�Xձ
��k��wmZG<T�&ؗ`[���~���_�i�.߷��t@!=��+�r�d"�j�y�5x`C/u]mFD��������LJb3��d#gc��MN.�9яL
GA:�����Q�*��6�c����ڔ�����V��E��A��J�s���77���W�u�HAd6z�k�sݟ��5z�v
�m���v��Q�H<b��D<x`l�1j�����>�g��#	P N���΁+H������`�	Vo�pJ>��6C8	䜬 cdj�����T�=
A�����e�Q �I�2��k������ b�A�n�;��~��n�ܵl~�Ƴ�e˱�������]t�܋��kx��lg�%9�^� ���4��;�?��{v��ٲ�c�V��K9F��'�z�6�+���v����7�F�zԵ,�V�s�#A�#��Yb\0�[()O�l�(��\y|�E8
��0���42�3��B@"yJ����T9���p֘WÛ���|,N�d��:��hE������F>����!B��^.�
�ff[ͺ��h*��ƶ,Z~���|h/^-�_���v���ݺ`_z�ͫ;��v圛5PH�na�{-�ze�M����[aQ�F}Ǯ\z�G�\����`�������7^��s�s�Uk�զNK_L�lе�hd���Ñ@���I������ҽ+8�p�����g�A�c�l������3�*%�g[L��ݕe>�N�v�Z��5�52�w��zg�������4���vnoK�\�7����2v���l4�>0�+D!���$�yl~l��%x/���\)t��	�ǿ��f�[6ߓ�v�X�ܼ"�Fz�4Ɛj\R��X�b��Kغ�{��� �8�*06���몂I��s	�?)���d���;�Y���^�*��Y��SF���a)��'z5��/ɀf���3��� ����޺�GY,z�nϺd�̓}*^�;�l����mv6���5迮#`F@&�E��BD���}�ji�In&�����GR��w�(¯a">����z$��-Ч�c�i;|�D�"R�̯D'�����d'kT��w ��O9rmgDh��߻��a���Ӽ�}�o/�ܳ;�wm<ݱ�lh����Յz�Q�v�U�'V,��fǔ����Ef`���۲jk���쏾z���U�l�=A�<��l<_�6v�G�@JR�:��VJ.]�6�N���Y����C�
d	����z�2��6���h� b(���܏��͐�\%6�M}]�Dfqc�.P�5R�A�~�0�˃(�;f�]Y��1�#�m���#�%��jW.���s����Q11�<:��Pl�d;߬��K�#�~Ξ�r��>:�?z��u�U�n_T;�<]Z�X6DZ8��Ė]}�Hs���f�\%kT����>{�ʹo~��/��|�߹���N��{A󭰋�3T��7gc;��N\.L�l�>J2G�����F��*[�e~OhH���˾.�& ��˦C��9���d�l���v�B�v�*���e��w�����������TՂ]8�cO]��^���[�?���l�|�D���wHPa4�t���$}c[��n�^.Fi��^�O��y�����n��M+��d�����"i�:;N��Z`���=�E�{67:����P@M�f�'A����L�8 ?�C�Q�y�:�sm������L�T}�C��+U}`�%�]q<���3oWu�3���C�U~D�%�C�kGf��BD"�\5� �+i�GbI�/E�4]O��<��J<���8N�qbwK�{�!�G����C��{�Z7�W�)P��#�ظ��'��{}�|�q�{��'�&���]Y�Q����O�'�-=��D(�eg�{�������ӿC�-��?�I�Ɠ�fg:��xiGGf��ڷ^ۃm�ر�ldV`�#`C��P�өɿ�\��VٖӉ�"_�s��[;m+�;���3��˷=����l�r�Z�˒�{	KXω�TE$��z]�XJ�f�~}�H@�+3G5���w�w����-�a*��e��F0�a��n8k*�tH"6��~�}V\շ�ax�3��S�@�� ��%NCb���w������h�o���5��+r`q'����C�_<��"f�y��s��KO�Ž�=~x���ݷ��Nm^���@�][�s�r�C��]��V���o�o�Y�*;�-o+�r�(䭞�Y�Y���?g��5�;{��i�):�[�ē�ԅ>�F�����o���{�z������Jk7�v��aHlCT�Ύ����1o�z`�L!�H2/�"2�%st6uԙ�2[*[J��x���&UmĪ[L����&�q�E��.]ڲ����۲�`������������
�F?���tl�Od1\���w`j^f�-���o��,9����RQ��_������V�ܴv�ge`��R��)B"^A��QيҒ*x��[R�o������z�럄��cAH��h�s�"	BA�PE�z�^�A�*�����2�y3pF��?��2�zO�d�]�lu>����0���!=1���R��vEZGR��J<6������ùJ� �F�@j��M^�������*_��ݐF@�r��6Bt�Q7���R�l��3�u�����sN:���ֽNs����6��>D�g��������q���xg!�Z���}I6�M��VbݰF\�8����a{9�lܵl�S�%�^.+�hno_ڷ^ڃ{6���-W`-��1T�{`n�n���Jmf��u+�i)�\B4�(���Ζ��;������W޶�^�
�][��%X��QU[��>"�'��VvQ���f�Dh�$��в�g�2�Ǯ����'��y�~8�����ֹ#�iW����
��$S��{����'k�E��	�*H}��!��Xz7���>�����:�{���ĈVa$������ ��u*���fs�3����~�{����߿mǧ#{�����l�,[�V��E{f��/\�v�nw۷�=��f�ڎ^��,j>g���.�o�3��I��p��Jź5j���TKm�r���|��+x��_|�j�=x���K������|��޾sf��MsH����4k��C|a4>���h����Ke��A�dN�IG+��BRߖ
`�� }�o�I-��g�4���L�)X�;��������=;::�� A�<s��F��gg���ƀ {9� �,^m�i�M��Sӆ�LU��Wy��B�(�V�g?�m�����UoZ�������C��fV��e.�Hv:�)���7>
&ZUA�t��L�o�P#�)�ġ���0<���a��N�z�� �ɾ�^�,���
�:����9�W�!`y�q��Hl&�>؟���ʊ�(Z�ASK�C�ꏖ�z�ZO=Z��S���u�^�����:���sl�l����z-�Ii�`���D��n$4���x塻7�����������;b��2���@gV&���+���*M^�������y�(20r���w	h�A|�)�β��L6�ٽ�{�;C�qcnG��67%��� ���A1?��V�*ՙ���.��,�E�� ᛫o�H��-����폿~�z��M�a�2������V��%>�I*Q&�iԇkE`EH���;��{%��d�@ϛ��O��Y\֗���h����SR�|�a�;"�vk
�9� 繓�"�%��
���W�)a��xMx���,�/i}��Zi���),�p�RPOEEM�T]�uH`FP{]c=�񙍲3M`�>͖��𠥺=�O}��������Gv���v��c�w׬޸�r��c/��ɫ��sW�0��WX�z���bC	ђ���c@�.����6�z���&Y.�]�{��ٓW��k/>���h,�����/�v�\������׮�y꽇��>��ɨ���
�~��V���T����J��\��Q_@�(����9	�K�����q��lɳD���:uyCH%���V�٨i���Ce�̨�L�ҒE�93��y��3B���� ��74�=°�}Ro����<�:�6�bޚձ��t�~����~`�܁U�&�$ �0���&җ��ȉe9�ȇ�
���a� �3���V��+%1�Ŧ
/�w�4�*�ƻ�C�^�jC�  ��>�fp39��*�w�����=ˏ�`1���j�Ĝi
:��G�&���$��6�\T�`8H������=^�)҄��r����X'��=py�C�ʇ���IkJ��\��#�����Иב��%�9%XF74��?)R2��$�_���}OI`$� �&9�	rO�v:�b69�7��݇�����n�7��Ӷ�5c�>[�v�Y�r}���Ejn�����Z�.�5E�B.HCӇ�-�-��;�\�lQs'�B]Vm���I͊����$>�Sp==я{!fvb�k�'��"�&S�v��N��H<]���2�_N�T�kJ�"q���	�s�=��<��Q��'ף\�v������W�+�XPz�@����Q��}Y�V\�9���T�S�˲-'��Nmxv�>��]����+����n\߷���������'y�c{��s{v���v��C��+,_:o�ƞ�3t����m7Z����ǮX���A�
��]�p٪���쫗��ؕO}��{�]��o��]^�����������o�����=���k�2;7vg�C�5�i u�3y���b�-n�ʈ�1|Sq �>�UcT��	�>`��ك��#_�&����	��̭���� �����'iFf�R�%�b���$V�N`m}&q�ѹɸo�!
���TN��`��o�:�K��������U�e�-���ǁ������,�뒰��� %<����~�4�`���VA+���1��5+�)��WS���2A�Y��6�K���p�r��������#Rծ+�5]9`\m���?8��6�m��ڍ�J�`Ǣ �*��@p:�P�Zl�}p�"�76����Jړ�������M��'!d�F/w�h�ae���=؄W�XC� ��e3u\l�)��)�䘻����`��\ m䞀����B�!l�c�a�����̮�m���s;<m(�N2�FO�UJC����Ǭ�t��q��EؠB�ۑ�R�m�r�^��M{����FsF}��X�Ҳzظa3�O����b$K�,����&mUVe��M�I6��4�����HV�����=�A�� �Y���GzYhwv�Cr�&9$�Mv7�U���J�އp��qo&{VM,�d#�2#o\���=�9�e?��\@&�������<�t+`�Ky��g�ҹ����|�9C�����w�|���.�ij��g�"	>�SM�Nn���Z��$�#�lF���#d��b�Qs��$6�_��jY#By1��/~��	U�J	˺�5¨���5��_{O?�D�{��v���	�z�!Ƴn޼�������Jx�s���=�`XD����X�爳@�PB%>����Խ�3LfY\�r���Z��6�~��W��;��?�x�#<8�=	+C�b��fî2�B���1�}�ܜ��9�936uq�W/#����ͣd[�b�r�p�TC�'�6*�0"u�0*$�v0���9�����<�	�[^�9aM_;BɆף^q�ô��27�+�r����^���k������x�f��d'C#_'w.�m%(]��#�c#��Ŝ�5T��	Dg��=^ߘ���x��@������`�������7\�Gw�7���Jڡ������7`�q��=�+�I��)���Zv.���+UfY+���z ���˜���}��֝����^�1�����18y���2[���%bw�~<'I>;W� �p͟�����ri��u6�j��*'F�A�jc��Q�tf�0�9���M�l;�QR���f�� �[��}o����J�YKpT�����M��Q�R*�H�<�%:��*W��nK� ^��^{W�6W���4�4���*��"�Gt�V�;�e��`K4��z� �ZI|��3�"�'�����y�'S�_&�(�M��2W�䓧��ЋT�`�m��=��}��.�_���$%h��l?!�%�0't�|޼�@9��/�RѸ�A������q���ed�Ed�3�
D�3|��:>��-�+��4���t�3<��'�E<��ӳ��h�d0�Ĉ+i*F�[�s����`m��G�p�b{kk���."\���ڕ�ߓ9[:�����s�p��{C�?���}�XLƘ�)#6So%�!�1��y�VY0��q�l=�Kz���1�S�rB���-7�zD���w��lÙD�(FMh�PSl/�S�ƊFD�.�*J�,����Cd�"��6��6�rYnS�+qu�k���$�(�M1�	V*g����x�����#�z�� ~�ڜT��g�XLC	�}�P���d����c����Z���uԨ�tf�e���i�ʴz0��g��Rs��3M����t�ꡆq;���ZY?}�fT\iɳɐy��W�0}`�=WG1�ߣ�� JI�h��*n��|�v�iy��^|�_C:�5�����ř���L�����K���x�y�NWlaA�6��^X�`)����@{��a�4׷���z�IH�h�َn�(�����?X��[�}���1`5G��E�j>�	��V���JI\��go���̾˵:�B�L���x����e��    IDATL�5d�U���k<eF�%�w��2���fj/)h�3�}J;T��`�[*��h�55s. ����>{��bՃ�γb������$�1��|m(�K̮O��c�N�����`�ݭ��6��1S�P�0{j}|��>����6"�k��ʕr��mf��

�a�\D17�Zc�^\�sϬ"�!��{{{�Lc��\A����ޭ;wqx�B�_A���ETBo2"�*��l��|�o\��ׯcww��X_����e���\��Ս���?t����w������[�ٳ�t�GLgk0��d�A�9������pAR�2E���H�K�/����D�mq[�c�Ҕ��CI����S(JI�Ef�%ͷ�Y�XX#���"����M���[�0.Bxq���o���&wG�(9�\�b�D�F��rr1�Q:�?����'�B�C�����g"��lb����5d�!���^��'��#���6������jU���`C�zٝ�&I��;�e ����ЗA��V/�B��8����'G�⥳�v����(a�2�n�-�&��'�j���$�|�9Y��X�D�?_el˚��e&����s̿Y�5g�xs7��l�������ۙ@�3M����?D�|nD(�gf��|��� ��5�ߥʟ���`4�D}b`���Y�@�I�3I�1u1�|���NO��_(���8=+�3�i�cD�2���X[e�v��f�f���%�9"���.��+�u��L?��[x��1��M�r9�zs]d2(1`ۀ�)���ٺn-���Cб�k�Y[ig��MkJ�4.�P}��0�=gA�>V�`5�Pa&���� $^��r��v�y��N��r���۪���=_�&9]��=�P! ��w�9/�N^"�Ty� 妲U,9ǹJ�
jq��_�ň2ml�f��a}��gr2��Y�Q������ν{(����F\�a���ְ�qv�����x��^|�)t�m���R�aue�bm��}���ٶZ��������{��7���ߙ�K�SPMcL�a��ZL�Ȏ��M��E���-�����Q�8���hC��Г����RB�d�f��^l�# f�!J~тI���9V녱��$5pZ;g�	hU�'�фRf	LI�v'1�M279(�g�A�ѻ*?�Hhg.�cs$U���������#B��"#�� s9��\yX�'ɼЛ b�����jI$�Ϩ��;�$��ʑ��]1��')���Xa0���'8��0��w�0����֎e3�V)`�nQ�e\�az�4ɪu�!���(�g�P'z�^Dfx�8$����8}���~��ȯ����"��3�e�).�D�+;~��=iw��gٳu�Gɵ���5���f�`CK������%/��\>�p|��yF��6�O� ��`<(��H�|��9���j��d��ޛ���<���ì�-'	ʕ9��.��P���l�mk��E��js*��ϼ���Y��|q�|�~����fW0��Ej����Ԝ-�9�����A�עā�[/U<�4�"��xE���ׅ���1$Rםm�9��qB.?2����G��Ť�L���#U���|N|I��!ٌ���Z�ބ:��Y���}��E]c"[l'W��? ����(oծʐ��Η2{�T1ʹ*QI �"�qn���X/`�Ʉ`
Baڝ��k��=�K/����m�����	z�1������pu���z�Z�����2*e���ؾz�.]��`�:;[�������_��S�{��nh��h��C0�҆���9�m��=+'�(���"O}�XY�$�@Sd�@mQ��t�9��Efq��ii R� \ �t���x���r��9i�M}8�{F%3�$��hH] ����(�-��,�4�Ee��۠<���	��P�O���|�E��G��'"�HR`���D(�kȅ�L�њ��*��hdɄ���	�E K_�P��~�Î�'���ֲ43�t���3����O�t&��%s1�6��lY�c��8{l/f��G� #0z�Q.Y��]��-3[�[�]��|)/��B6�vZ�O�ǋ�6}�đr.1�����t�2��������4�	���_��otᇴ�U*ETܱ�7����q������L��� c��z���]]s�v�no��;c����wr&B0�a���b�F#��F�7�gh4��M%sG�D����ɋ;�fpis�y�����wv�����ެ�)�g[�������(���,�F�ENA{��� ��|^��@ش�m�xۉ�m������m�{��
?���~'�S停2���(�w"��L��<��B透߫҄u��X�HM�4�h�`)]�9����>1�#�tr��d
j��Û���(7Q+��Zgen�(7A.���Z�����`�-h�����짥�L������@é�[a�Z��Q\��j/<w�'�ȡ�B�\�U\�t�kW�����F��9��ß��������L��ɨ�����ɾ�l��|�l�l3�����)f�9����m�Ԝ�I�g��DU���4K8![q��%>7Vr������Xr�2�0�'5e鄹 C$��K����@#J��|��}*+
;C�2��4��Yv�dd�� �������T�	�!���t�Aˡ�� �U��f�6�4IΟ����;�����6q@��ܘ��U,+6��W�7�t7�N�V��G�ơr(3�x�l�4� �U�H�lɿꁄ�J�ig�$R��Ren��0��aP��/T(~�vN8\D5{Ƙdo�9�.��}AGڱ���k�&�����π��7��(�[^��>m���b�l�L�Q+�����[�
3�^�0pa���
�x��˱ Q��I�$�H�yz�Lf��c����dqzV�xc4c6�٠�{��9����-�Y�T���%�i�E�K�+u�u�^����An�q���(sT#�9Ҵ�u��t��P^?m���i7������� ,;.H�0%<�x@B;�Y�*��s�Z�규�3��d���s�v@@F��-�����F�f�a�ɶ)���v��9��*������ہ\���PFUؓ��k�T	��.2�uO�Y��6��|z�A</�Z�Ѩ�x�94W�������Op��5ll���_Gn��8ʖѨ��s��V9�A���|	�[[ߺ���������#�y���Ə~���o����|0��l2���##�g+��H�=����>��@�if���M)�6����ڡ<3�a<��s�kt�Y�0$~�RX��ZʺɃ��`\���AD�y.3a��D�_:aw�<?8����u��2����t*���iLc�G\*�XfF�kζR��[_��o|��Bfqv$�nq�f�-؈QVf�-ed=�|�-����hӐ#\���Ω���;����KRFNz݉��3��~Pb�C/)D��"p����y�1p��f7y|����В6�>})��os���abkIB�Ζe,��[�+�^wg�~�;�m�=t�s������ h9b�waM�}�6="��r��,�g�>��6��/G�BO7�ӗN;��$.� ���a�3��p�n��t�$)���8<>��1����ࠌ�.	-����b�͍26�#�ԁ���2��t���ƖI��P@����KT(#�V���?���x�?@Z�p�?�#G���M$����$�����rm�0��$	1fa����s���r�ꑙ@;U��=�C���C��*υ�h�� nr�"!�R�����*o�)(i�t��:~��v�ԃ"���wS:V�V35�[�D�g��4>�Aa#�A3�7��0C�N�Է%M/� G(UJ�q��?)�W+^x~�<{E���گ0�q��M|�/�������BC�c�F[k�Rk֐Ͱ}���+t��3��ݸ�TP��>��9�����򋟿����x�^�����h�X:[� -�K���ܷ2r<!�џ���X�P��L�S2AG�֠��4�d��`����]���-CV=��l3o�|Sy6l_9'�(}��I��Ir^V���"�S(t|z�2g4\�ٺ�VԦ�eمΖ���ը�o~�
���2J�]2c�2+���Ψ��A~ND2ƍF�6O��"�0(�Уl4��z�K�'�Wu�<�^<3�
Ip�v�0��g��9wq2���_
$�;r�>��m�>r�Q��Wa����-���8[/Y�����.��@b��(�5�O'����C�����}�ˍ��2�;����,��]���l�ߒ�M�]��a��3۴�����Fҟ�9�dN�J�iY�乥+$�,����Ύ͟Н��ݛ-�z�3�T�"�Bs�s�����w�p�v'�&z�:�]�=d�cl_��ʥ"���M"����|�C\��~�a &�Է#7o�VE\.a8~��{�ٯ�Չ�/a�Xcx��C��ؿ��R��Zd�e��,2F��0O���if��%%`�]�U����%#�'�36Q�'2E�{�<��+���#.�r�}@���<�h���XbSԓ5��C	��'IG���`C]�Km8����QF�*M�"#u ��G���y�u���{m\�R9�(����#���w{��#���gq�u��޻�}����ؾz_������b�I�r�l�j뵼�(��.PE>����ooo?����~��|$�-��~���޸��wv�xҞ�t8���IA�nF��aOz�������b��b��+ڳE`��a�#p�22T��ר	)�-�::�p\ӓ4c�i�14�m�&�	urE�n�u2���f�RDeF;07 {L$�ll����UD�GG'h��`b�xP��٨�9����oJ�����.9�|�|e_�r��.
�!2����s9��f@lE�<%X���<�QD�m�86B��� E�28[�鹺��}[=!�IW3�	J[�o����w#~ް[6�vFˬ{�7�����SHz�?dji�l�K�.�L���� f�� #�0:w���~��'.�������b�e�m��������@ꢳ�LR �p���&7�k��|�O�&��t���fI�X���cr^�:g{�~,g̭�,��3�i���L=���5�2C�G'�j��ǭ;-ܺ�E����x��BX����Vj�*Ds���%K%T�Eeb�EI�j��m�!WdO����.������m#o �F҄+`�,��K}�pY��c���xf��Ԅu���e��6�\��-�|ۛ��l�K�=k�e��!xňQ���N�S��=fbZ���l����!Bѐl��� ��F.�D�grJ��O�����et�̀��F��%�KY;I(��0j9��p8�P�VEy1�Je�o�\�T�O_�;���!�+i��cϾ��߻�ݝ6��M�eI�գ��(�.�@��"���������wG�a���8�Gg���՟�z��]��d�����'�^�dH9��D	Ȋ�w����&-�-(�et��<��-�l�8�'\���ٔ�x({���2^=hѠl��&$���ї���Q#��Sx���	�>g�B%Gq �ƒ�)�\F������v.>��,������"E�t�R�<��� ���U����.�E�������-� g;Y"�
,M�gˌW���6�(����9[//�a�̖�t�0q�癘���9��#�=�JWΗ��eX3&���!-K�FϚc0��㿷Җ���4�	�=;G��4�^X[�6�Z�qY*]|,�S6��,��H� "Q�I����r}�Ƣ|c�-���밶�����j��.�-�����4i������7 X���y�2k�3�7���#9mF$V�⩜�z�ҳ��9V�Vea	Pfs,��^��V��3��pz֐��p���d���kuܸV��JV����J�y1	*� �S�^w�z�����ȕ(U�8�񳟿�7�:@�_@��*���r���J`1���U��@Z���~�	3P�t��=������0����������.��NM5;�l3о0��/aI�}A�����9U&���>��WV�4*Y(��$�+TiL��E`�y���A�Y�ֲ���,�E������5�H��L�G�DJ�1�þ�"�D�|(�`�>k�(��z_��3غ\��！ÓC\޺�z��8����]���������X�[��X��Z}�问��ի��~��wv�/��o��/���[��8E�.f���D�LL	�}�Yd���eyyB�����qr�$���u�y 5�!��z�d�*�Ij	��_&��3KE�#���������͠���e�9�ћ�� m����q<�屸�y-,�+����~�HW��H��@�eG�����W���/�Q��PȘ��\�3B���E	���@V�a���J�[ !��FhV�jC���Μǳlc��0���KuDv(''�?IgPiN_ݟ��:0�g[2s�v����Y0�^δ�fK6�Л�5� ^_r#i��"��RLN���3}$����/+�vKg�鶅��yG��6<�T����%M��a3��� ���8.:�0�k���q�n�MP�~�z���?7Ԯ1gk�Rd?3g;��q�>��^����#�J���8j�����89�a23u��b�����2������V��"���T��6�R��g��v�(�bl]]E�D�Xz�{���)�}��YY ��"�T��5ϲ��y�� )躲�3U:[@��A�V�sS\�Z�N�#����ێc�:X�����^Da�A�)���)-c?ɞQ.�3�>�l���ٌ���44�Xn^��o济FC��h'&㡰8Q>�"�h P1�Y[YE��Q�bo���]J�"�|� �U�(` <�@cEdHZ3����Ѭ��܍\�n�`��d!���^����x���U|��7P)-09;Vu�X��R^A._���?�r�ſ:�������d�D#��O~��W�>���hM�a.g;p$g���Kf�c�Hd�],�d'#��c"��I�E�=�L)��~�����x�٨��7)݄yB-0f&���|��m���ec-FR�љ��˙?+�Y�EbmE�@"ҍlVY,7�C���l�	��+��dن�^����\d��E�,��gqn�z~�W����|1Vf[��X8��9E�g3+H����(����,P@�L�,3F��/s�Ƙ�$�H��3�����l���^�/+/���C��s*��#8Ls�FG����nC��<�W ĞZ��g���6�"V&�� E����؊����2�w�]
8���K�~��/��T�h�c��\e!����X�I�U��<ӧ�U�v�˿O$ӟ��Yw,��X$R~�}��,B��Ͻ��l�JթL�tF��� �~K	4�r*�9�힜-�~N�3��N��a'��g+@~�|n�˗"\!�9��Z�*�x#t�cL�D�P���QY��*&��#�SњJ��9���~���"�������\���=��:c���X@[�����\,I!h���|���R M�"��?�*5Qf�н����,>m�s{�� �P��؞Qf��8Q�����3�5�,<���ֵn�F&s��E��L�$L��NTu$y�LεH�rQ^�S�6.d������1NOOq|�F>��ӟ�l0�h���"o���Ҏ�J	�Ҭ4ѬE�Z�ak����:����1�p���ƣ����Ϭ�k��fl����*�u:�?��z�_�����G�H�����ۯ�ݯ���Ǚ��tp2ʡ�^����a笟(��|�Ǽ��|�Gv:���D�ŏ'��Y+#unV��Yb١?4B��=ztx|N%��T��2�4g\�`i�J�	��7��WY� �0GEm��"|���ȓ|��e��xn}^�|��,�N[A)���X�b}}�RY�+���_`%�㋟Y�|.�r��Zq�|f�l;C(}d9;�H=�/�Ȓ!z��yк�G�0��g~���s ��IH�E�Ff�)�3��k��{���t�Կ�H��6���,N�P���F��F��Y�,Xz��w������Dk�er���
�>M@�$�_:�#�%    IDAT-�m$ʃ/������f��?���K;fH�x��<���0EbZ:[�Q�`�6	rl�v��F�<i \��Yf�C��{��&k���-̡�Msr:
̂�5�C$ӡ�5꤃�t��<~2Ã�%���N�gb��D�N������<�i�b����0�i{�����ڼ��9����qq*ɷ(�(Q�N［�[�w1����Ŝ�#c٭;J�?��G[a�}���9b��M�P���$���r��ٻ=��+�2���f�KE�zI!���z�b%(�-�:�>��( Ƀ�{���hW²�V�.C��s1[��x0�~|p�	F���{�(����N~V�RA�!������Om�� �Zg-k����qMZ�;g8<i��idr�q6��899�$*��S'�#��L���R���Z8��pxJ@m�ª
�+5���.��JI�f4�"�#�E�ַ��ֵ���9l����wo?:��{C<9�L�2�y��I�MjEL0t���^��D5�ɐ�@3�t;�Z��7�y�?U�W���R�!��f�h��<I%h��sj��q~���9��=&"�D���s�3Vփ#�˲>���/��"9^_�QCc���W��`��O����:m-l�"sd���r��!o4��^� <@ÿpuc�W�VD9~��lG�t�bI�`B��Y+	88�@Q�q<*�Ѣ0G�����i�Ό�`��)*V���Y�����A��	����,�Pvd�\��tЇ�?�rQN&�1���:�$e�����?_^b
�d���}L�j��.��>��0�TbZ���U@�zvɵ�,Յ�Ճ/���U`���_`%��oMI���@@�do�"4A.oԫ����,��I�kR�fp�h<=�U���qy��`ɞ:;����z�r�Ԃ����h�9�L.O	
Lp��5�����U�`R6ٸ������~���Fk+5͚�c�C��]�Y��R����M����I�@+�Yeʣӛ�۝�ӝ�����6&��U�2Ѳ-E�2�
�XrȞ+�H����kcwcR��A���霽��t�����h؜}TD�H��"b�9yZ~b��Yb5b�������֕]'��H 1�pi'yTb ��g�d��� ���ep(n�Z���n�''���:~\ȁ@�Q%L���ޛS����l�A�s(@,�{��M����ߗ�@w@�*f�\�N445�̄m���L#��-�C��AI��
,�S;M�ZD����+u�7k�gt'h��q��_�|y�o/��������O��}r�{G$�`�SĄ�	�6��FBǕ+E��G=9��b�b!LgZh���g'�O;99�h�Ӣ�n4V�Dc����4**��H|le��c���..:�S�`���:Q����bd
�������,�A�W��x��#�m}����U�m��0���5���K*Rsf�$I/s1����U�,*�9�����7X]�&wP�����3�<�I�i
*�P �'��,GR���эj���Y͒YiI�@q�`4�vQs�!3���@�Y���:*:8j/���9p�����4:H����f�h��xT���H���Y ���]�e�I�Gg̉��iJ��<�hɥ�r�v�B�;U��y��.}���,񜳺 Ԡ�e�ɱ��N+�'�HĦ/̌# ܨ��Q�8� �D') �����>|K���<����Y�^�S�y�߁����ζ��xb B�q�q	��.�	N[�:��v6q�_�`R@�?F������ؾVB�Y�Zsq�*��C��D�P�o�V�P��#F$m��LZE�&�
���ƋN;Y�'V����+�h�e��OM�@�u����P�MԲ�X��Z��^��Z��YM�)w�hw�#̘��H:\'\q�*O�4�����-n���yB��#Li��Hb�v�z��+T�e��in�81ahwZ��s�b�W���$�i2!�9�k-��ڬ`}����u�	�~���4Bo8ŀA�*hk�5�B�O�RQ �L��&��p`�{Ł�d
ڗJT
Y�w��ԑ�fT��hn����u���	�����S����ݽ�{�~��b�����1�5��h��U�a4�cF��p �؜�^J=C����u��n��j�T��{��X]�j���u#	��m��za�6:Wfb�l�E8gƆ�`���?M���H"R�Yـ|%@Ƚ u'��z�&��E]�� �Cމ�;{���5��ʝ\6R
�J�2�q��b�+����7�H�����z�B>��������-d�q R��ҏzx)%��,��;K�<��*]	ҟ��B�P�I&�lu�lÈ�J�賜�Mz���aV�N�ʭACU�_�eK�s�!X2�؏Bɗ������R�Wo��CzN��ni��r`�Kd�����z/سX��^�M;ދ�m�eC�r��z �Ǭv²�`YR�"w�z�F������T=�J�yQrw��D� 8L�)F+/�'�۲G$P*�ǅ��jG}9�|��B\��i��ǭS���y8���e&��8k��������_���v�z�f����4�a���PD�����J�ʰFa�*6$�)
�Kf:N$D�BI�g�������!Q(�^��*+Z�j#q`*g��NAb� St�B���ull�aee%rk���Ɋ��c�@��8o��&�0Z�u�y}�Nj�,�N�k�~�Ә|��M�;�l�]�9�Ұ%�����%'t�RV��"����	z�� �}��J��r1�Ri��f�ZQs�G��w�:�/S���r��J��u��rcF-�v�ԐsUBV3����Ō��R���qn�b4�j��8��/���eܼ��ݼ���G���n����O~}w���U�����p�Yڢ�k��^Y�Ypn�%OS�
N�۝S<|t��3T�%�j54�+6�AR�	��m&��π��#� ljh�r�\�������
�>I��|v���q9��h�Ԏ2��,���1%s��l��e�JU�S� ǋL��t9W�s������(_�$U�VC|�U<�,���{x�e�@t�)��r��<�=�@�eM�G�:�2��݅�$�2�"�r�<���r*sz�L�������F����?Ke��ϗ#H�n��K�_YS%���3��T�P�k����y��K�� ���ey�ʫ�X`d�ke�ý���s��$x>K�t]�{�x�t�Hڏ);�qS�~	|ʽ�	Z�9��T:�c�3Y�T�b�����K�	��P�f����1\��� [��#�u2�؜���#�'{������	Yn&�w!��5�}6���)��>n�k���*�K�e*����LF�\���O�b��t��Ҫ��Q�o4����K�	ph�g�}�A�Fa�rFK86PM<G�7�Y��D�5ә2���%{�En�U���Ge�z�Z�bI߳\��ރ����`H��yR̆����3VǤ���Ãm_{�|����5���{�n��]	+�$�@�K�14#�p���.����!N[�zr��~���ؓ΢X G5I����C��a:'+`]%}:Z��N�G�'h��8mw0Z(i�{@N��+Yi\p�Z���U�<P�NQ+P�Ш6py�n^{�?�q���;��~�$ ����g��ݟ�~��.bf��/��Ii9�3�<��N��?C�z6�������s6��&�Y�X�W�qJDR�1*����և�Ո'A�i�}8��l<dC��an�X�u*�f�C��6	���*V��LG�d<V��,�ZtaR����������k� ������aφ��e0Ҋ	eQ-��̍n�a�q�Z��hAZKF�e�*ق� �9{�c�#:[��l�@A������ۖ}ܥl�VS�%y�^�M9��>���)İe��\��\je�;��O��lA�,#0Og����"��S����9�U��r���!:�)3�v���BƜd����Y����d��]��<H,}<�ә�]/���=��%���$�:���*H�:g�*1�L��C��,[^��?W/����q?7�����J �SXVnԚ�q�L.T/1�������!N����q����1�m 59]��|���<>�B	�:�M2bnk�7Ѩ4A��q�"�}�XW����o��V�36i}��o����3�&f3�)���JC��k#h�}\����W�"g�0⊰�hx��gNB�>�Ԁl��E何��r��?(�#R�(0�]d�u�k��i������4S�c���Vy�\�(��v�aϰs��F��:��XLȩ0D96�b:��;��h_�(U�`�>x�Y�<>ii4��lQ:�c�uzj�Y�A��@��]�\!S/�Y�)UeP���b������������������0�{�?|�;���������K��p	�(��d�b�� C�	�6���(AJ��d�f3=0eߖ�R:7C�Z�ɯ��e��ۚA�	�A��eZ�A����̈s�8G2A�KC�0F��76�X̸Y��2N����_���a10s���F�ҵMn�@�a����ٌ0+q���׮Lq����'�Wϐé��)�5�Ȗ0"Yȴ+�[n�(WWn�y8ϼ�٤�[���!C��V ��eF��2�Ġ����˷N^!��P��R�e��/���������Dl��z6e�7��B�Uk��.��Ѹ��9����i��5�d?����{��p(��x��0p��+��T�����޲V�� s��^�_�K�I4q�~�c�˅�l�����*�Y@�
+�{-{�~�� ���X�ú��Lg���"�ё�)0&^!*Tqt�B��G�l�no��w�xtP�k����Y\^�q�F��@�4l�kh6�dG���E����x�|o���g-nbN;��A���;Ax��'Lgt���G�%f�%oo�8w�Yol\B�VQ&K*D�����[��@���X��;R�Vh?,�� ��/G�A��{�+*��2����ϟ���O(����lo:0R�)e�<6���q�� ���fŎɎ�Zr�����g�[�u��/<�����)&�,&���Iv�0���v�LB.���%���0�N��w���S��b���X�aց{���ɘ�
*E�@�Ȝ���n^��_<s���������=If��I�c�ׯ����}��Ȗ�҅���|)�U)`:�j@��9��z�!�mHDGK�S:5��#�8�����cڗEyuY����f�7����VV2��Z�&E@��k� V�li}��sr�t�ζ��B��(p�Ҏq��2_�\}��亖�lb�!�=�,6W#ܸ㥏qiu��2�]d	~�9�|�&�"�I��.��A����	��q�f��/�������θ��2�Þ�tH�'O3(i�%%��YF���`��H��3c��n@I� ?/3Z�gk�Fi���\�gg��.
��Yy|�R+I������'NZ��N�<^���{�|&zr�[�i�g@=;���8bڪ4L�u�TJ���m�e���,3����Eg˹v��|��M����K��g��#�]�t�A�͔�(#��������e�����NO3�u��'GU�r@TR�����Ե&nޠ-�#eT�-j�W�ה��s��'?_�#2��"e�b�&J7�eKA�Ơ#ʮ�(�v&��t���B�l�Zu�ƪ�ttd ���²j��3,"wx��C�����ZPz�%��Y0���ԿB@?%Ebp��w5��[���["?ɲ��9���A���{]t��f�{���2Ý��8�sv�^��~G���:�pL	?����P�>C�-�樔�ܺ�(.�|�G?8<��I�YFζKy?�I��r��X��j��8�C�P@�^�J����]��>������Ƒ~��~$�vg�������΃�>�7�c�<V%������(�94�0�{z��)i�3LQwӧ% J\�2�*P�Q��S�T�
�=��H�KեQ��W9�d#�H��}A�%Pē��r?��,Ȱk�#���q�8p��<"qs��M� ��(<�&cM!.�n�Z��Ic���f���nl�a�y�(�Qv��8#�:[��F&���B@�|z��a�ed�|�w+�?`����$�*#���������q؈��im٪w�r`�)lY�;7��q��H���b<�YQ_�I=+��;�@e�HB��ن��n�8�;V$< X�D����3t0S*#�2�Mz�s.��j9�`�L�PT��8��gk�v�L�z~���=���>�z�X�jX$���L���i*m�����,4����5�Ld&��4ְҔ�

������f���;�:�=*a�b��a��^,����sU�
Cą�FCrY�r��V��E`220[B�G�N,Z�G6"܆ �)O��HZ�|l�xO(vOA�ry���u#�GOb�6��@L
�pV� _g$�0YP���7����e���Y�kɜ����z�^O|n쳪lD�e�DGK�Ri9��.A[�<�V���9k�J 2�
$)�
s����= o´�ɸ�~�x�����6��[O�5G�Y�RA�_�b]S�vgݞ��z�!��	r̆9��"l���c㜮�ʪ.V%4��f?�}�{�ŏ��Ɓ�6��H��ǧ/��ǿ���N��N�=�[p�I�x2TI�D�����	ƃ�~NRn7�\h�~W�>w�e�M����$�� ��m���K��v�@#b��@|���ͅ`5i�l���Ǽ�DI�
y���]�x�jF�E ���v��8G����Δs��)gG�e�Z���d֓Ǯ7W��C�00����k�u|��>��}e�Ji��JQ^��3�WvB�%i�bC*;��oTuX6�sIҴ������#,Vt�}��9�Y��LE�k�4��x�v�5wr��8��D�����7 ��t�[�2' �z�6o�Ќ)7��o�ˡrp��x���1~%�r$�^��Z���9���tI	�� �zj��7�;[3| �cAy��|
�5>e�w.�@�����5���`'��t���b �\Ҡ�&����%Wr(x� Y6f�ZC�C�}�{�l��s����a N�>�^��}��[��8�ԯ��2���Ox�����k(���7
(�9�C�ӽ^YYQ��2Kn^���l� L�gزt�h2K%B��w�}c8&�$��e�9w�-�R�����s䣚����Q�eւ��l���֟����hc�/�?��,�vr�g<�y�d�ݫ^����$�3ߓ^���Ih ���A
�<S{L�t���^�����Dt����
��o�C�I��u)R:��� G֌�`��N6}�z]����.��3�e�k]���Y [V6�����YW�Ҍ҆S�c��F2-& ��ҕ�RG&"1����R(��J��K++Xm���/|�s��o�H?�{?g{��3����ko�?��=�L"�G�E0N���дD��g=sS�zG����3{%��dB�b���a ���e�+W9�^Pc>�����J,�2%!��K��(�Ӗe-F�z���+2F�)Z��Q�ZȊ;]Ε���tiVFd�ǅ���*�)� 	�L�V(��+�C���*�"b6�c��m� o_ZǍ+<}m���6N�ŁDJ��(�i����,��<G�T0��^.��N�v������専���Z7H�Q�E*.��Q�I�rH> �*
��t�,�̟�]b���I�I�i&�U��'a�3�Л���H�C�%�`+�:]�!����gRZ��
�K,'����rps��-�'���~���iD%���ʟ��L[KQQ�+-����$)#����ce ���g%�0O��<_��ƊԔu6�@��&�o�Y�y{���총/u�q�� �F��ρ���˱J�!NB�������Q�'��z�'1ƙU̙M�gsM�g�ެ�3����fFΖ��"z	�"S�`�v&N
v��U����8�=f@��5�1E����e�<G��,�|��B�����re]���m�|IY9�'+Grt��|@���z��������vA�=m�ns%��'b��7K�Sjz,�� �;���F���_��i�38GqV���	�Y��N�±(�i�0mTψ*�=�[�    IDATJ��"'6���n�'���'�4�D�ʬ8��VT�G��6�Ci6�Y\��c�jq��6�X<�&�Z�N�P)R����f�+���s����a�o��پ���?z���{����(`2���2՟٤'J~�j<�b��>&1��\<50E�%��6��x�ٛ�������j�`)��h�C����'�&&�ǇM�:#n���gy�R��O,��C&��6-�T|�������H��A�Md|s������q�T�:�P
�&-Wjr�\@f�á@a�B�˫븲Q���������^�����"�Ƙ����*'!(h�>�]���(dfGc:S�n9:�d�	�[Z�%�Oi�_�3��Fu�@����s`Y��gb0��vCN��2�bjrd\�ee}�� ��A{;�����y3��(O��C�<5�$�u@ԇg�c��ݟ�����Bm�i�Dٹ�r��Ξ1�'�q�����B���������2�q��j����:��� �X�<{Q�`�H��R�y҅s���
���!-�Xて�e�$U���+������'���iV�T�6�-��3ԓ&BfQ��Qwn?��v�Dh��@q�|	�8"H���U���n���*j���
%�=3[�C($o�3�J���y^>*��Z�|贉����R��2(�TYG�q��&r��ا�\	��x���-p�;1^�k0ل���4�fp����-)H4l���K��21%��8��,Gd��}Zw�b�QW6W�@^r�֯�ߨ�<'/}B	�)-�����#�z�#%El!�*���gݎ�
�=@����DG�����ϊ�9�u>�r���g:ߓVm�!J���vS�"/��V+X�ױ���?������o�H?�{?g{����_�������{x먏ք�k���!���q�W˸Ԉ�,-���a4h��n�X�i�.��~oI
��/�c�V��>�	��d��Ɏ����(����)ʠ��,���K�;F�F�=U����|}G���[L������zJ�%4�����}F�y�9,ohR��ط��f�iL(I)�z�Z�`���Q,�1�R�%L�D��j�Kk�yu��Y�Y�csu��f��k+edsj0p�39X����*�x�0�\�ע^�}x����19����D�F���̞Bf�k3J@�Iʻ6���z�rp�Dl^�f3�@Wt�ޭ��F�(t�!($��>��e��MPV0|է�Ηp�8�w��V�a�Q`�Z�P^:��T��o)��O8f`�Ѭ�䲵{F%� &[*M%�ʔD��dU��x��)U��Ϯ���3=U�f\�T�v�!3J��e���s&����Q8�K�*K4z W�'�xZg]��Y����{{x��;88�_G�WD���Lc�>&�
�,����/}�&�{f�JNڸt<\K_� 2����3:�)�I:T3��s�wF,9PJ=^� �I���r�2��+(�ԧeOzJ�ҜU��]�b&��e`�+w��:��3Do��XZsb�;_�_:3U&�'�
'���A�<g}�mc�A�JjX�,��8˜?n�9:[�Fi��崅z3���̤�`0��TAɋ�-�+�l���͑x���<��G<هg���2�̿�Ћ�]N�%d�k����;��Y�<%J�ܔjZ<��)A��%��j����_�����@��|$�����������o�����)�Ԉ�9�gT|����f�� �ޱD��� ��7�u�!i��e�ʛ�Fʳ�>���zd,��֭[x��`�\�6�G�@r����P�65�(jP���Ys��N�h����:^x���q�����Ν;8=i˹s3#b��3�ld�#+	�5���u��K��9>rǅ&�f
�{R\26�r��}j����.��#���]�5��ZE��h�J��,��T%7��!�!|/�k���0	�~��'�':��)A����_xy�ь�9a�Dd�"K�ء.�*�|�=B�(p�v'�!�I�i���qQ�5>��@��L� �M���;�E�e��f��e}GԦ�=�4gz�k�糼+��w���"�3�'s���
�%��]XV�4���2�D.gP�*,�ӥ�Kg�j�2��lq� ��N�������,����6n^N&B�~7��ߌ&3�Zm��j�pz<�ݻO����Y��H0_��,��h~�٨��"��W6��?x����KY	���6QuM�G��>� �vYFv�E�%��NXa��A�A�/�A�e,(|Pj�^��biq��-�D�]��Ü<����t�8" ҀY�.���}>/�F��|��s����dRB�K���{��/;�&�B�Ytꔶ��)Iuk�����e�C�at��Kd�����ၥ���Tl�k����� " +�p��i��(k��{x��F�>*e:�1�+5�E۳+��h$>cz�	���p��$FA��\��@gШ��lo^���{����8��ޏ�پ���������ͻx�`��a�Ĳ4C�¨��F��?�2^~q��t���P/U�nw���vvw��Uz`^ڬs@<F���^�SO]C�\[T��o����}(��llhd���u�	3'�7�����9�Yr����@s�:;�I��9z��{��Z/���^��&�?:�ݻ�Տe�G���ֳ(_����5Ǎ79�ϣX�����'�8= �'@�dI��U9�Gؼ�ĕ��Կ�M��0�b�����R$��J��h�:��x�h/�<����27��<��L;��e(��5F)O	����(�qh{�2�g+�]#`gCJfwM�]=�ؐ��rP�;n�+���e�t�d)�̨��u(^�����ud�k��h���-)�' (/�eM�_3<�lϕVS�67�ު�lC_��6��>�H�R��A��ɽ�{Lr2�V^̡��534=��%J�����*����s������z6��ʮ�f���4�B���
��K��@>>�H���5��QO�_:�|��liqm�q�����Y�K�������<+���+��E�R�l4Цx.&Vbϋ*�9����`:��I����%��+h46P��i�n8�j/j�P��fH4G�9^+�?c������� ��+`<ȩ�r(�9��}%�x��.ՐX���}��Lw�����Vה}$�P���tz�ޝe�R�g͜��C�IV0���-��D���%������$�R�����g1$�Q��ް'�X��m�`���l�u�hVEfė��x�A��S�O��c�KZl�Ř�~�m�|�8�r�2r�e��sϿ��k���?��m��8����ū?z��y��	�۝�51pDo�E.?�t��Z��?}��Oc�z��Ѯf�j�:����������.��{�iq���ի(�8k���XB�e���89>�/���-�1frظr�o���Ǐ���#eׯo�(Q,�?c����ZD�z��{ʐ��.�Yk�Ν�8k�*�V�x��簽}U���X���;s�\�M4�eo��IC6�k׮���>��O������^{�<|�G�?d�D*�S����V�)z�M_:p4��9���}�=~��x&:��W�������&��q�� ��}U�xnV�M��m��\`#
� 9�ŧ�f��v(#S��zxևS92�2�9�DG���șݨ�V������M����a-:��}{3��¶ ��s�Ҡ5�ɞ�p02U$��/����1c0#�e�� *,��=F��#:y��^&N����GS��
X˳E���eI6��m$�ˑ;���-1L��73rt&"
�q��_��x�˖�R2ή�_V:���r@�:B��]^�$���D��0]`4!���#�#i�x�g]DQb�(=�\��|e�Q�EK�j�!�,��/<�o��i�(FϾ��zC�_�-�Yd�-�3��t��5B�1��\�V���f�Q�_B�ZGT�	]M��t�eb,RR�TyD��T�k��r�cF$��>7����i��)�
�_ΡrfWU�@N""��v��"����*wt���.��A����c�Ȇ�=�0%"�,gۏ/:������QN3�0$%��̎��sf�8cE���(��-��U�JE��7-ǭ�Nq|x�v� Q<E��Ө��C8ڤN�o���_����)u:�P:�E�ĳs1�Q%m���Z�q��2D~��_��}���_��G���޾s��G��L�h��P*Q������'_}��ۘt��c���޿}�w���l����*�z�TJe	sq�]�s��I�~�<x�H�C��p����W��
b��/~�Ew�ꖌ3L�\o<���.Wǧ'x��7ԛ}�������צl6���K�#&����{{���=Po�Fq&���Ej�1��d{11�R9������/p��U�<9�~�S���=,P���}��oVpu{S8�ɣ>K�]�<z���=D�66����� b2��9Dv���(��<#�P��t�&b ��{�5��e�9d�nP,C1�oe�*UF���A0��7Gʾ�=M�L�J:/�w�<�dbۦ�Bp���m؝	4��e���F�qC��p
`�&3������{H����/��'��,��<T�qΛc��zԲK݇@�`M�d����J��m�$�cZe ��4/�0X�7�E4��G]E�+ lx�NE���E�MP�>����G���u���.G�Z�rV���}y���n�U��3�����������"��q-Q�՛��*������-��KI�9�*1>����?�VW��L��dmM�-� WI=�� �7�����7ZA\���c�X��m�Z�i�j�m]e"ą2&�Fc����H�{�|���f����[о~?=�U)���͚s%�b���De%餲���~�L�w{�.6�5�Q����p�+��]
%2�� ��`b�|�����)�:�u���u���т��Z*T��372�e�5�u6!Wvg���!�2����u�4V� �d�cQG���>)>ɪV�Dik�F��+R�Zk4����3������p��}��������go�>Ļ;}��s�R � ^����O�����E�+��<��ɓ'x����d��2�f���5*f�(�9>>���*�,FG'��u�ޭ۸}����I��?�c9ٿy���C��W^yE��Q���<+g��K�Ң���9į�+���7�|]�Z�F���˸z}���:.����}CZ�Y���{}$��&W372K�,3�z���O��׾�;��{��~���I�H�z	�B�Qʇ���ԍ+"�2n��'x���p�X��O�̨u�N�ݣ}���D��z��[JS�>�/�a�K!PL�s^�b�"g�Ҳ��2w��?MC!A���ލ���(�X4va֗NP1+ka��c��@���l׌��i![t�$��1t�U�h���_��c���P\��F�!J����GC��d�r��Qǜj 
���dɹL�w�̞x�%�l'gá�=�����!^���esx=�ʄ��4�d�-P�1)3f4��@�B�pQ� �#E?�a���p�KG��'S�"�4���ҢH޷K�.s���T`�ʘSg?��G�)l�����������"�"�z�Zo��/?���y��^àҨT�=g�G��q����5�Ŧ�Ȇ$�7d��Z$�����UԪ�!*�Z5BA�ˆ<M���_3��*��̚�����+
����Iu��ܶ���%�*ڰ`Ъj̈́�?��Y�N[�����rݔ���03st�,�B�F�H�`� eEJ{H����,�z�سm��qy^�c�,l�H��a�l��5BD�
���&�G�;���w���(�^V�

nX3\�"F��@����=V'J%��Y����W�������}���ٛ�q�p����l$��i)?�F���O� _y��KD(+3쏺�H<�����J��V��QYҞq�Q��S��w��;�h��X����g?����_��^G��o�ڍ�x�hG�������.���/�c�����W���o���ܾw[�Q!����x��gqrr,g{��9[�OG4`@vn�NZ9��L�92f��r�����O��?���	�ſ�k����;`��E���|�޸�f���u<}c�(�ɨ3���prL*n�2
$수9�73ǰϬ�����fC�:�R:"��t<��\�Z��#%���:�t���	����-hi\w�B���(\<"݋��J���$		LE.�.g�N9?c8	�v|�CT˕��d`%/�-6
?��q�t�2��W(ǥs�l?]'K`*��5��U� ,o��8g쥼ev�m(պAU����|��Y�P�1����IK� ��X�M�@������+�|�=�T7���xLw6r��OC�[�{h>�\�,y���rm˺��;����e~N}J��3x3l{�=�g K�yN��d�1���&����pi���^��Z����ٔrF6C������TF�{!g-.�����
Z��kX_	���2�d��k��R����Y��G�\�y�´dQ����V�b	L2lCҖ1P���W����=��5GmN7���$KG��l��zm��Mmi�`Ӄ:�Jt_,hЋZ����ن��}c�t���yx�����Þ�#@�b�eƯA�B+���g)|����r9[�a2p"9_Zˋ)�����5�=�,g������{� �����}��o3=�
��E\L-CY�([����qYI%�8�+UV*^RIU�$Ne���I�r)�ٲESA��f�`���g���w�o�����n&�`�
���U�A�t���������<�sҹ�H��X���~ﵗ?�SF�}b��W���o����@���ݷ�.���������J�e_���ګN[	�ci��zC,
���t�Q�e�X�R��׬Ď�P���IN�a��{c���޵�/�U0B9���9���[
�T.��G�s�>�n�N���g��o��o��~�fgg�_������ا�{o�cw�ݱS�l��!���c��7o�������I0�����Ӣ��)y��I����_�d*g��7�����%ku��Ul��K��mj�l+�Sv�Ȓ2	��:�ww�l�L[6SL��4�鷺e����]�6wlñ��7*8�dPe*kA��S:A	�Gc�Q���`�^����y��9�S�� #7V�1#ָ��X�pq�@K��%�0f�Z܂r]��{�+"ye�6d^��'��Z�Zb�'�/�V�3��aL���ܽ&����m2a..gB��`�|dU�T�2Up���=_*r�O�o$�D(���:4W9������xS��p��i�pBNك�I
4��Qq��E�C�G��\���~��`�C���iDb?���>����1��Nt���A��xl�|Q�6�7Hz���࿑'1��EFl~�l���6�����?e�O,���}���	�}�瓴���'vt�ת\ޔ�x`fϊ�M�7IX��b���h��B��#p�c?��A���(��������;Be����q��1v.�C�3�&��|Z�r�"��F�����b'[��W��j6uO�j}]�8�h���8�VELB*�O�����5���=ĕLog�h�wX^A��=)�����;
��ڎm�<�Q��*�TN�� �:r���-�Oz��BA����nAv���M����d2�3g�~������_�`���k��7߾�_�w��xܵV�oZF��T�'F��_x�^8w�ғ�3�4�^��� ڶ�Hة욑��9��m�gMd��ݡ������.�pic<�\�`����+��ĉ�v��	�s��{p�N�>m/<�������>uV���_��UJe{������w���t��_z�;s�z#���v�[Όs�-Bf�@���'ψ(Ł�I(����w���j�N�����������hR�Q2g�Q��U�+�
�l�^�RW�@Tջ��\Z�X�A7�7�>$�r���kq�    IDAT�l:|��ǵ�.Ds�AĄ!�U����u�͡�~0���h� ��Q��D8,Ja��a/��`��L�(⡭�9q?j*1��bZ�_����A��j���s�~I"�l�6lAK*��tLo�� ���]���q��J ��)"O������6�X�A�w��i�#����6�D;�׎}�X�������2�F�����;N0�2wB�C����.ҵ��m�U쉇�O���zP�����T����Q����e���u��FJ9jLD˚�5�{��A��g���O�b����sG�㯽`�چu{u�= &R�O��MH$��|6'#�Q��
R���k�SSv��6;D���a��m�RC����e��'��)c%�	I�!פ��;2ŵ+�@�]�]�]���?)+�K�}#7�̔�`�wyaQI)��GܯT����M�
s�C!~�H2��g&�d2LC�$m��� �JN!�|ʙ��RV�V�(e�n�ꭦ��?��چ|�I�%�g)g�F4N�V�)�Ř��ޤ���1i�|�2ɒ�se�����{��/|X���U��\���������
��4~��Ⱦ7��-;��������©��VHO[�2ŠJ�K φ`�^C=Hئ�T��ʚs���eZ޵w�}�޽x�u�af��¢���Gu���~]��ڴ�� 6@ɿ�2���W^�{kwU�@z��U[ZX��'O��|����L�L���?+F3_�nݺ%���ZC�toa`��S�U&^-b:�Z.��?���d?�S���/��?���o[2S�I�dM,�����|֖���ȡE�*��`C�Qk��]��b�t9����?@'�RֲɁu�;d���UR�R.�]��� �/�vسy��4���]�?5FC���0�:�wI~Ae����g|cƯ�U���p8R�8L��/ė�{c;,�$�Ø�����w��f��K0i�uգ���A���M��:�̧�y%��R9L
�Ѓ�6T�(Z��EH�:�Ej|��k�!��TӅTV}��:�׉�|�j��*��(�g�}�21���\�#�����^|�2x�}��FD��x��Q����҈$�d!#����+1^�]��ٜ�e��
�Q����;;]��9cn��L�~�K?��ۭm���~S�Lth��=$)e���>�0��[vq
7��5�c��?m���	�Tr��!���l#����= �:Ɍt�q�`H@�`_�?X9���>{�ׁr{A,&7I�.�B&U�0��9*i�eT��5�ܰ\(�;��=�k{Lu��Tqo��:�������g�����m\�{~.Ȧ���;g�ÿ�3w0�[�TT1�9�ڽ5�p�C��qN��9!�屘�gyb��633��}g���Q ��23L��>}��gN�������[�߹��_��a��ִ����Q�z����ZJ����Kl�]˧��9�Ж�b�Ϟ,9��-l��6��#Ű��ٗ���\�f��\����+U;|��fM޼y�6w6�̙3:	�de����g�	:^����flan^�K̴
�4.<mǏ\{��}��-��݄����� �Pu-�2y6F*a곟�����d���}����߰La�R٪5��G&} ��c�Kv��6�����#?z\��|��{!�QJ/��׷�uU	��g���.k��z�g�&��K�3s��yTS�3�8?���I�[�|��1��Ze���a�R����G�.�'yMj��v�� =OVLɀ�x0ƀϟ<3�=V���Cf�G�Y���H<bU���VE�7o:m����������I�=�ZpR��,U�!cU@���Q�H{e����r<�� ����v��AE8������OL]��C�1N�r�]����������H��U�M�}�q$p�X�)O�AO��G` �&؊I��X��X���-��7��Ԡ߶����8�d�o\��`�𕟵�_Q�c΍�1�+/خl'"�龫�8{>Ĝ�`�p�i�̌;y�fgf,���������x���`�P�#���:�8��@]��ε)i
�]�r�b��'T��>�ش�bA�5<�YC�p�����R�a��;$�J�۸"�]|8�1�<�DGÒ�Jx���דN76	�Y|F�V+�拗.٣�G��n^��!�(E	�	����e�.e��y�HyX),����o���+��h��|�o����o�w�?��[���˷7��N�v�)k�K�u��)�g��pפ$�X���ĝ���ʤOSo�(�aD�������i�����׃��o�#��EevL[[�x�lr*��t��j��&k� /�u�G�^x�Ο?�E��[���;�`?��&c�1(S<2z �&�<����c���}�����Y:?#�?J[��	�_�N_�����<!��m�lskW�U\�苑)�;�֪=��-��l�b�B^��*˰IaT���j�`eA�wݩ�T���<�88 ����l$�p(��%B�ܛ��$�����X��I+�b�D�(�sƾ��Zá�6��W�*&��� 5�p�%��@��+�x�E(�u"�[��y�7��v��9u��I�����ߓ/�C�C���5����'^O�<b�+��ˋ�}�>&*
p�u�]��9h��Y�Ѭ���AO:[��?��K���`��R{�K h	R�bŊf���+���?�1��G��1�;I- ��@d!� c�AOi�f*��8mwn\�^�f/=������Y=$UC�߶tfk[%d�+��G0�qs?pz�|�ɉ7y*m��o�n{l���C�<��B�I^	˧�=!K�Ӛ��ɓWv��-?5���.��X�D6�|��,{@�wi��J���x��9� [�l9w��k�����	"����*�=��=�p?�OHb��`���H�u�-��i��U
T������c8k��\�L=|�n�������0���c X)y�-��
}�c>#ݯ�%�JM��ꊝ<U������|��W!�P��~=�`���n���o�޿�e���V$��^���Fu;�b����=w氲�䐩>�J���'�8\�j�l�^!�jҳ\���lu���˪lY\�:��>L�~�c���+�g`=U�L$�P�abᐴg���믿*(�$`����,"2�t�.zAf�r��p�d͘q{�����v��i[���6jmK�V�0i�((��S-�ԉCvheF�	���v:��hǺ��l�
��؜b���jm���n�l�R���%�����{$���\���;�u����2Vo6DF��QWkޣ��Q�m��'%�P6l��!|ps$,��X!� �:y�����I�R���^3@��s4ҍSB�����X�/��ZA�ʡ'V�1Hg��]�$Y�y�{m�lB/-���0@[���{x�S掕�-�{�<@w��%Vl׉l1���� ~�H,�	�'?=bn�}B^���}�^���˩�WE��8`��V�+�0L=�43�1
09��k(���X���:�'����5{p���ZF	I�,�vΘ�	2�dE�r`й��U+y{��f�VM�����h��̧�.��][GDO>��丞[�d�$�-�CZ7���}o}�666?�dG���CV�m4�B&�'w��ېhr�0k#�㉶��B(B[$Vi������`囱��{8)�-_,X&�Q�FҚ��9O��yMf]�T��oi����8ΌliaFxġ/1эg]$��^����Ao�\���C�H�?T��Z~J��`bY�]���¡-���m����ݽ+i��҂%�}磊����1�q]�c�v��pW@)R���O/�{h�ЗΞ={�C���şH����_�o���`{�1�� i��I77������C	�3_��=}bɒ�'Jbr�9�T
ZItqP�@S M��l��ҥK�(�"��jX�5T�޸uG�,X�ׁ�΂�Й4�� �����Ci.���cP@�{��Yk4�ʎ�_~�*4V&ȑ��v` N�/3p�'�Um�-,��Ҋ5�#{���P��Zk��RF����,������nwF��g��"���U�>X��}k�nJ��<?gGW�X�\RFO��g��\��ox���<��� �S�����a�x0�]�f�S$7�g�7a<`�^��i�u�g'f㘿Lش�c�%h3�l�51Ľ�����޻������d�R��N�?��}v���D�L08X�F�hd�D�����z��o><ȖV0@�!`��M�<�"��+,��c�0�������ݶ�*�ؓ��?��x�.|}��뒡�����d���sFIm��L�[�[LaT�g��[ujZ�&�z�$\�Z͆MU�V̦��ز�w�A?{ꤱ?_|�EkvZVkl��J����������*Ri�����d�/�Yyj�r��5�{�pS����?rԎ�Qk�Z�(ؒ�RY�4F":�σ��<ERԁ^�Z	*c�&�W��P�b�ޓ��82�I��\�Q��nO6��o��nmmk?�\D���ft~��h��znT�Zo���`�����O|]�P�g��#��Ϣ�ù��뽕�3V��}`}�h�µ�G�)C�|^�?��Ġ�v�Ţ�&��.�\ϼ�����"g���[��˿x�#�g?�@�{<�`�'�]������`{�!#�2�Ǵ�6W2;�<��|�5{��!�7��#��)�R��[�e݃W<��U�j��v���T	[[5k�[v��=�}k��=z:��������W"2F`k��B��i�GJ&�,ꕏ�$w)�kknI��C�T�gtP3	hw��E�bG?��U� ��_\���kuG���["S�Bu�{��ǝ�&��ꂭ��Z!;��d��	��ng`�|E�ݝݖmmo�u湇c��|h���dLF�K9|Ȫe��Fq��t�������U���zh;�X'VT��a��j��ڐ�p���M�3;��1P�j����H�=�ZA%�o01����� ������\{>k� "��bY{$��$�q,B�^	f��=Ә0Ġ�F�������t�v#�$1��$�أ��6�� _�*�|����Ī �H���/&� �D �F�� | 6�5���P(��}��5�J���=�g�uD��w���+&>�F��K{���xkӮ_�n��F�Ӑ	v���[� B�>>	p�Ӗx)�����Ma�){ȗ_|Ѿ�s?gK+˶��@���Oo~��q��\�PG��: �`y&������̊Y�5k�%*�Jv��I;��ls��4�s O�^��پ��-Η��g��D�H�����h	j��۰�)O�H´?¨@�X1ܤ?���8^��6[�sOv��VK�H���g���U�C���+��g�ؘ ��,���@��T��*�%���NG&2��Ǡ��5�Jʆ.7"(߽�>~dk���fϕ���u�nZ�T�b���O�)�$	,���$����W������[?�@�ă핵m��e�T�:��n0��Lad�F�g����1���6�:�4W �a3�)�8�\E'�j�v���r�r(ld�[5Ut���2�Z����0�3`�L��땖&�/Y��݇�������Z>i�6�ٳ�5��#��ې��vaa��SӪ���I ��m�a���dK�ׁ�����[uz^~�T��Q�2�i�����I%�?�h�V笘ǝ�������`�{����:��Ŭ��k�n)�r�!J�8�:w�-��:�>µ(��J^�b�Q�%h�3�"Ǡ���2���5�:�vxq/��=*�?��9|"��(8A��űj��F֨���G|DbT!&���a���Ǥ�/�f�B�˚��~pί_o�����`Z?k$������2�."�����Ҍ�2�?����ȃ'~|q}��c���(�R2���:���C��rܫ`c+�I���7�q�!`sߣ�T��8�%&���M��!.�i�=�ݿoW�^U�(g��y� �L֊�ґ�g���L�	��~�!�O:��i���W_�O}��6�0/�؝�{�?��=m�b���g����\A�%������p��v�i��Kv��I;��j%zʖR�H�����`m���J�5��Q����EdwSuh�	ߣCc��@l��
�B{Fc�ܪK&���i7o|�j~f�j�<uޞ{��.�#߻��؆ *4��I܃��xvƶP0�eN���=�����(���蠚 :��������P��6lo�X�qB䴂�qξ���"�ægM����4;;��zd�/�?��o�(��o~����[�gW���Vm`�d�:���P�dӎ�������"��7ǚLA�f~~N�%I'�)���677���M[�[i[�]�ĝ���|/M�`g���*M_��؇p-�[A�{���CU=�l����	XL�aa>���6���ꪐ/i!=~�H�i��N!6U������/j�m��W�mt�E�
NV �umv�lǎ΋ U)cٵ>0��iKf�S��i7o��C8���rA:����O1�I�Lر�#�8���Q�9��^.'���j�|������}1���e�٠��ß�I�}��(�����2��b�� ����� �B&pރ{��éPt�(r'���Ý�=K��P�r��Jƥ=��������4����	b����j�����U�b���!�F�j�g,��'�̀��}`Ӄl`��מ�0�>��c ց�u;��~��dB�UX��GE!u�&��0~^I�(�w`89��cA�{w�>���U=���w�*�)����ߙl�R��&cŪ�gOE�v�V���F�����=9u��̗�d��9��ݶw���=�|lI\��0��u�G���vK�xqyI��ν��ܲ�����ö��d�BY.eи@ށ����mA�!�泬;O��&����z���w�&{��I�HmZfT��_�U�c=�f����C�ur]|��Zӕ2֯G�O}�363;�g�~w�O����Vȩ�<�0G9���W~=��p�
�R�Nd4��Z��5[u{���� w�ɸG�A2a�bY���$e�q�-.IA��T:r��bH6�E�,��(��cG���s�>�����o���z��߼��k7���N�4�A��a͎�������3'�-1X�޷��׭�m(�..��<��UO&,���v6��-�ښ5w��MŒf��~���C�cOY����dÁ"$�{z��i�=q}�YA�>�(��I�ހ�_z�e;r���,Zz�o~���훶��X�(g4���Oٹ�>b�A�n�^A
o�d�"��ф)C��*ڑCsvxe�J%|ha{�d��AL"��z�+[�-%r���n�ʶf�T�*��aI�Kv.��@�!��n��ڲ)8%��`�aż�t�*�Iz���C{9�o����W�*He�Q��@Tt1p=����cSFBGtX� �`�n���V�~��Vs�%�K�
��!���UH<�NU�I�6S� ��@�Ht�{��b�P+�x#{�nSN�+h����"��IK�V�,�AS)��d�Pc�͆��I�b�ʚ��Z�hýQR����aEUN�!IU��@�BB	T<W�b%ʽ�{�]w�Jx<������(��~\���Rղ�iKg}��={��iaQ� ;��/`� -S�jfd6c�y�^z���޽tѶk[2��t�%[�*[1_P���[U�eF]NTm�����5�>��V��Ҳ��̪53=5�y��l�L=<8�5]���wD��ВA�lH�;��Ar� �8<�����s�&֧����N�a[�]���fn߻{�vj[�V'�~��?m���'�<0�ѹ�����C����XD�#^G������+�TR�<��8R	�G�}��ln���[T>(���T�b���Ҋ�K%F�����^����wt��_:}��?y����7�{k/�6�Y�#{ ��`ˎ/��W��Oڋ�ؤߵv�k�o����{�h-.ء#��D�?�<����m[�{���]I�Q�[�2m�"N!EY_�"��YN���?��8���_
�&�2;ql�`�%\�����0� )8\uSB    IDAT����ګ�c'O���`d��~�������[�l��UM�2�z��g>k�>���?ڴ?|�-[[߶v?e�T��c<bGr���D�:rh�P� #��O�ZϘ��Y"k����Ff?�lgc�M��R�������Z@���hu|,�ϪV8��)V�� �Q ����&�� �8���8����X`Ǫ/y���4�����}��l�s҃���)��CD�������]�OL8r�"����Ņe�n�*�80��a���������L<�8c����WE��&0�#���.�AAQt���l!���`���zS�1{�y80��v�%��ߣ���YB�3��=f  �!Γ&��c?>[�X���w�u���M
a�,� ���$�~�o�o:L��ͺ��k�:c��9�"�@�l�������%Ƃx{�E�^���i�{v�����S�`�5���H�g��e^á�m5�z��"j��6��G���Rz����L�J�g�D�Z���i ��A�9�G��0���Y&���χZPO��Y�V�m��3�HIh�Ɋ_-a"��͝���߾�f�/_���{����.�s�?����_��v��R����p�8Z�� {�fXGZK`��"_��k/!K��7��w}m������-��	%+�v�s[=nF ��6]�Z)�S,��t����8 ����o]9��=z��'h�X���ۗ��7߹�רl��I�
��ć#�[�Vg{��?���z�%��4Ѭ>���8�t,�0	�WQ��ҧ¬��xd�5s��65p,6e@h��Aİ\T��@Y��6���>I����1\�V�{_k4��	��fC"y*[��矺`���1;{�imt q*����߲K����p��3b~�_��U�u{�~�Ϯ�z`�A������0G}T�l�d���SǗ,���qF���5}KeK6;�l;��	��vw롭ݼd�1R��2)���ʨ��Sٲa8D4-�\
B���$V1�M����i�L7�+[`d�7T$�x��7$_�GCRd��<����{�����4~F#��%LU��6��[=z��=!�k>4�G��C�ɼ����&M��{V���&���:�ث�}8Z'�(��W����E��f�U&ú�􍹥"ר�t�o��I5�[��שC�A,���ѳ��+�|����w$�ʖ׊R�X��~]L~�O$#�V9<6A���#)����{��t_�-a�ٓ	���[6?k�͎�=����w6�Z�٫/�`gN�;7o�;o�����y�ż��	+M���_�t!g�������P�����L��V3g	/��5{-�&�V�45�6m��!��^�+�V�E�s�z�j�u�$C|n��oT}{���=�~
���D�5��
7�)hDb�g�/�������4����ݽ��nܸ��.�	��B"�K���쓟����hw�l������mtO��<�mz��y�h��7�-7(A��L��֦�I|�y'���G�g�f�\iܞ%CBֳr>g3ق�,���҂~�`��ȧ3*�V�����+G����B�I�'l��Ǘ�ַ߹��W���n=e;��u�~���,�G�R��O|�=v�
)Xa�@�l&�N��J�ff�Ef��X��x���8}��e�S�i-�8p��+ڮz1��i����(s�	*���6A*%�Usc����\��g���&|9Y<�wԆ��mu���>{�.\x�ʥ�=~��lr��к=�}%T>�s��+��^���rE���7��]�r�v[#A��I�2iF���Z����Ge��N㊄��o���ݽ�غ��;q�2��M�X1��ڣ��v�ݷE�"�n�����5�/����A�Z��T�����(�gkF*��sP%��
�Ĕ�C/Nԉ�D�mt=R��bc���
�3�e择>��Ͻ�j�{@�%i#�ab����Z�w$�Y1�(<z���^��옍K���i�l�R�D$X�}���Tv�Ģ E�-����LIEGH&�*�#�@����ܧ�Dp���{�Y���F�=&���q��~�W�ܚ?�0p�tI8�h�D8��]*�ו�i���U�eLP�A�R|O��s�͉뙚�վb��o��u;v��mA��ϰ�����s�.L������2�R�Z�^���Y����=��k7���w��1��h�,�Rflϼ�^=j�}z]�޸V�`�I�[�'*>1�y���RC��t]�!dB|�a�'���D�ʹ��Ug�*r�c  �MHl�'��U�3�^��B�4WY��=��m��O#"AJjB�%H�9�i�Ñ�[m���M�v�=Z`�Ʈݹs˚����g�?e��˿,�����E����NV����D��38܀��������l�ްF�m[;:+�`$&ZŊ�8'x=��D�t�JՊ��=I��s;�0kǎ��wƒ��s%[Y\�;O?u�ןt����D�?���տ������յ{4��V�i3x��Dv�j6;5��^<m�N,��BE��n�=�kk����gQL�C#`��,���$�e�m��!�`��@ءgCF�fCP9`8J�L�PtU�r&	'>=�DR�=�w��l�C}����|ѹ~��737g�Ν��Y-�Ǐ��>�=��yk6�v��5�u�ɳO?c/�����]���}�w�f��ܲZch�f�Sk�բ92c��,[*ճ4�і�F�gw�lص��ҡV���3p���:m�w�Z-�fX�i�*����U1w�w�Te5tBA\SR&d�x��4怇)I����`bg�ҟ!��T��� �M>~h-���y$6���S](�vf\��k�	s_z�$B¤���'����Rff�R�]B���j����o8��q�JW�r�d!t0�@���B�c�D��â�<�=�Ȍa����¡en04��T e�a
j����4��CZ���&�#%�j�	�z�'I�꥙����맇M�_��5����SXY�re��A�p���C��FyL��=>�ɄM��4�/��҃w�zf��p��We�B���iK����}�#0�[M��yl����S����8y�Rɉ=�O�����X3�v�#���Ҳ��-k��_8�a^�����T̻ot�'?e
�r��&Vk5d)� �����$��j<�Lىx����>�e�dd7�<���3�� �zW*^C�oI�DTr	�3���Be鉕��h��F$�lc{�.�Ů\��$�9���;;T�O �){饗�s��\`�;�=�z�d�!�d���4�LNB/˹y���f������?z���о��q��� 5j�S:�r�z]�-��u%�TP/�E"e���./�ҡ%S��\�r����c'?�px������|���~�{��������.�Ë� ױ|�o'���TibS9[��Ȅ��U��[��w���!`�-7�h2���t�V��nl=V%�æ'
�bH�H7���긥��Zg��Pj�*�A>��]Ȕ�ٙ�ݸ����>�{�\Ϊ�'6d8�����wt D�;Hi�d_���ӟ����߻������ZTǏ���'O�%������iwlYw��1Kg
����"�ڑcsv���%R}�Āq��h����{v���V�,X:W�T>m-��[O���]��d����Vg��ʂUI��4bxl���ٽ�vC�\�Q6�L_�P�c" 6�m�ru���}��i�F��ܹ]�����PI����r��J��Z�fkG�:8�\��|'�A�{怞�Vl��#�8� ��^�`_�~�Y�P"D��*�0sU��s���
�C%�"���Qgi �9	��Ӟ�t#��ܺ�4��qd��`�H���EW���
s�4�[޲�
�EK�c'��h�:ҥ�k!�U��Zvku�F�D�7_���&eəZ.i�C��c�ӂ� <�7&8�T��jD�>A"�y!g�@������ݡ5��1��ִ��o+X�j�5J��-�.(q٢���EZײ�wo	R���^��nkw��=UoH�j��@�	�\AA�>!𦯳��O.'���Ug+���5�ʛ�v$n���ƮuC1}Q>��Y'�Y�2L�G�@��Z�R�]��>)�]�
����T*' ��g�m�p���¬�!�!"��J�HbIxR׮ߴw/_�Q�33�h5��5�Y@׬W��x�j=1�[G<��%��n#q�݉j�v�"�a��G���`
k�w��0$�Y�9���0�>�R+���d�$8~�H�]���Y�*H�`����Μ;�����'Z���7/����{��6k=+���8%�`��	��;V�þÿt�qY0��K7e�7��ݱ����S��8p�F�Ł�̏T=�0��[�+��y�hs �0��Ò��IKP�=9qr�l�ZU���ۭo�&J�
V��ּW�H*,�(��*�(�Q��c���}�����i�y���eT`�T�¾w��,�_�E��t�l�~���Q��jq�ؼ�9}Ēi*�l[]�����w��Y�F�/��1�q��%'�mL�j5o�/���MW�J*8ȹg�ۅqvL��C���#�ݑi#�g&Yy���$ӳ��(�U���X�aT�8������y_A���T "�1F+��Bx�t�jZD�r`W����T�d\�*���rĮE�&Y����@F��O���f =� ��aL_	`U�``��G9
�y��G�"YqS�^�G�1p���)_�
?��_>}��5-�D��`˛�ru_���@��'��礲������׎�(���ܔ�A�	"�Vel��V*p�+�M���*eV$kTT{|f=��[
�=r����}$��@�|Ҕ�,��f���l���ʣ��ڮ��]�		�3_��]^�׵v�#�ڤ�D��S�ʅ]+�M����S@���X��qR)Z(A`�Q ���A���U���vxeَ=������h��6��Xg������w����vi�O�±J�M(��vwj>X%eJ.!YNU|��̔�s��c�Es��o_�Y�C����O�*��h�&��.���6w-�Y�X�7�
%�f�//�hߔ�=;��\�=�=���?�1�1�bY�!r:K뜤�}�ܮ�f&h��T�&:�-�skəM;�����܊_=b�٪�o�pl�����~��'����������ƥ����]�+�a����T�q��?0��UW������c*#J��%.@��l�4�~��sH7��ç/�C�PK3�Q&�L�\��J��� �Z�%8Y}�m��!��`�2�$mk5��~,�Ⱥc��\�`y�%eT�NѻYZ�5����d򑻴`���Y�) ��l#R�
L�g��P���V�y->D���ۥ�7���]�f��,i	|��1�4L����i�6�6����t��g+J �Kp�tlT�~(�GMߦ�f�y �$!4xU�j7�Y#��X()Xy���n��y�|���yC���(�6{��w�q��+k<Q ���~�k]С�}����!����,���f�S>ie4K�*� KFr�@� ��YZ����ͦ�VkWlT�Ȋ��̃����%s�զ~��ZQ�,D�81)��X߽~�D�f�\V�K�]y��{}$@�i�u�lԛ���-���\�*@��H(�>v��#/!��!��~ٍVܢ20��+d��=�dq����g�S�V�i~`�l������E����^#��{�іmlcb����8�w�..���C+
�jZu��:ڟ���t��#]������3��*4��-9i��9"����o��򶲰(8Y���6{㾞]��R5�����C{���ֈ�T�3���15R>�ԏ�s���b��|~Ng�����)gS���4,�����|J��V6з�P��4�;iv��1!@��m����Q|T�u6�'��f@�:�@i`	���i����NrB���=7�Y���/]ur�ۚ�'�F�c�Vۓ[, �X��L�b��[.��Um6��ós�~��>"�H���E���sO$�����?�{��/3���ꪲ ��m�Å��.��	�=A�����˃BH�c�@�^�a(�<M�#O=Ad'U�b�b���(i ���d}_L�n`�F�&��x���龰b�3F�9����A���'H�7TY�3��lβ9X����Kf ���Q	{fg�ņv���3n�z`ׯ�Y��.F�}�AJB�\����O~�;�~h���Y�}%'�V��M��:\���W��!Ά����5el8���Hw�L��[��x��(�!�l9bZGK��'YN�R�
L[�#��r�hY 0�����K7���m��b>c�4&�N����?�`�����Yt��q�RzMI��h���jA,r�����3�5�*V��^�c���D��s2a���'{H~`�;A�	<%U�.�+���;���J
p�����I�L�6��5@!bE�\=^�Ψ�rI���D��]��u.��S�KRR�h3��m:�+� ��Xۻ�u%��B�JժJ����c�جi����~��J���qf�m��!�V
�iխ�j��b���/J�:���l)ؓ�Ir�ɮJk�f�k�����-_gM�u7">��e+fsBG--���`�Iڵ�C����*u��=�5�{ɛZ,컄�������PPӗ��҉��ly6�G%���ĳ�=�4͇Y�2U�� Y�~nq� ���@������#���֍[>ްє�Td��lH�|R=l]_���Z��H�HعN��T�"�m6^�D�{�n��l���%�lg"��s�����V�Tu�Ȼ��fmif��?��_�)�m0���"���>�`����{��{�_�*�#'OIGD�ա��X�F�~OU��������S�*;�e���	Ik7��@!�p8��$Ӣ�e�`8Y�z���WÒ��+c�Rs@+��$-���V�
9x���߷�� ������="|,x(��;��Y\e�2��Td���{�=�<S,��[*͡����E[LYB��3r%���쳵�k�oY�� 攪[�3�;կ����{8�ٸ߱\��9�)�f����u%)4�i*H4}���$�BA�Ӭ7�L� Fb���>A�Hd�
�{U` Bp]l�� ET!l�4�7y�	�f�����&�*7���\�n~n��ż������X#��`L%b#����Peq�Il`��FT_^E�+w��$,�O��RЫ�m*3��Jۡxt2O�`5�<�=eM��<�"��lZ#$�]��Ir=8�!��Y����5LĭC�q	��?��̳W�ZZh��!�0m��<���Q��,�s���Q��cu����Ӝ��
��$.�"I�	mk[�8'.\����w���6�$����s9	_ �s�BLܛ{nvʎ=l���6�-ޱ���i���U�S��m�F�n���T����}vtǲy1�����7��e��z�]A�AsE��0+5�
�\F�RZ5�^O08lv���L�Bdu��#\��ӆ�2�F��uT�!	�\#�;��$�d�G�'_�@���oH��z�"�u8g����ͤ��^���Ç�j�|�a��Ku 9�ԆqK�h�������'�@�� �{�uP�BtJ��裘U��4N�oO��@��;�6_�v׶�NSz��;{���;~��W~�ӧ�D4����Ώ>�`�O������W�r�����Z�RQuǆ�d�3�M��J�!ːͳ@�mXWP(�ǖN���C�C�DB~?LXy����ʉ	�XYeЅ�LTfb*�sv�	ik71��lG�d�a�o)���R�H�t	JT]4�y��Q��=��(���9����C�TW8_��^�h��ﱰ ��װC��,�,y$`���ft�M��sX
X�q�>"�o�d1�������sSu���!�ß��U)���wj�8������,!�<�e]GԣrO%��&���Q���S�|��jA���`�;������6T3�!z���� ��i+�T���>Hy@DK�n��`���8����ױ6Ӡ�F6��#���3���u��*wuW    IDATu0\��=$s߸^n�Y���b��둴�b'��Lp;䎆	3LYO��>�iBK���{�^9���YL� ��F�	���g���5�+z�����2n�f|�AJ�����n?H��깅�t���c�<)�C5'�KAZD2�07m����\�z����s��qm�F��A̓)0�L��C�{���;����R�`�;�~h91�]c�$t�>�{��5�r�GtM������T��.�Z���$���Ft�tGr��'籭�T/gT<�^�O{E�s�:Iāq��5���LF&Z�B�d#�Š�����GղT���i;�HOX��B� ����=����K8r"N2�z��e�Xh=s>�C��7	,�8^g�ю%���P��N���'���c�|�?����U�H���o}�y��K�V�k�-�Y�:-W65Y1�b`U�Y�r��@���L��l4�
v�]������ �%&w�Ђ|[5[X�*��F<���u)e��a/��ovA��ɔ�6���aM�Tѐ�4�5۩)��q�	��~e��?F�9��pc�I��=�#Y���>�>���ύƱ�k���X�4%itma��_�1Ax聖��� ;��]gjSM�Y`�BD�9��	�V0�zd�7�M��C �F<3'�j�� ]RM�I "���;�g�?߈8�d'�ZZ�@z�`bA� J@��u���,�H����E��3ބ\���{�di7a���51��$�naN�=����La�j�����1����=~�Q0�94T�f�L0��ꀹ�a�$@M�a��%�D��7G��F�k�i�7���_���k ?D��?)���! qm|I.��`y��������P�!f�M[p��{�t���PG�`s�H�HtGc��%�-��J'$\h���f�6?�&�5�[\�RB��rI��5�H�%TQ �0V�U���=����4�
�9T_���5�-�L���ag�2�=иB����"8
�{7�u^Fd�d!��sQ�҂a�� r'����*Ap���c܂$*��U9��IO֥g�xj[�	&9�ߐ�	FǛϋ�E
I0m4���A!C�`m�`����*�s�������s'-����T�b�Z�㜒�@���$I��[B7ZͶ5�:4�N͇��"Ž�۹����H�S�%;~���=v؞;{�_�ُ?�Å�緞H������__�t�߾��e냢Ya��1� ��u��+n9�F�f+S���5�[��<�����Y��k�|^�X�L�����Q?a�ʈ�J��^Q�Aud�r����*[ld�㨦�ᦝܤ9�T��}�, �hXqp�	��b,��s�U���&5U��L�%�A`�1���]��'��z�P�Y��^���ii?E�̀= lyA�X 	b,X�t����	�͟h�	sW�`����TMI痶!�k�D�%'+y��+�`�nȧ���k\�z�(;w�6����C�󾢻���d�ϣ��)ߴ����͝5�$:ޢд�$9�> $lV�O�G*��\�1�ɡ9���g���ML<y��4ס�{�)V�)�q }b���5���n8�lWJ�`����^j��qq�����	��$4�������Y�� yE�J^#zUs0�9x&]M�+�Ú����{Ŝ0�d��%��~�7����	F�B���V���l��׌z�H���40rb��'�]X���h���Rɫ|���כ-�bYA�c���5�a�߫8�\��s�N4x��@�H�\��,rd)�6����N���s��4��>������H�8�!�����j2��273eG����YU�Zk����sP_��Yg�g'B��(��^��.��I6��z�ꭦ��|��8��I����܃�3�8o #*���zJ�`p��L����yqn���^�CC���hsC���t��iwmg��$	��Bkh��a��pbX"��\i�f�gm~z�NY�������������U�L���o����?���[][kd�c9�����4�P	S42��;��;v��oY6	�a�	����-�ϩ����}e�T�ȉ -�ϊX!�}6K*�@G�&[*Ho�c��v�:��;��ZQ�H���+`�;�H:�0�B=F�GE�BYA��C���pW0����Y��ł�L�myaގ?j�!q�"آ�#JN�\^��$.g�3�633��G�@���/���烉�!s�#D/���	1�6����`qz�sve�*����/	��_X�qs )	I;�4O�!b�7
n�������\IC��~(B�ٗ8���'��p1b˫�ޏ5��7)�d�h�5ل>�_���c����akKstճD��K`b�?��,P���������`�Q�
zX�-<%�D�Ʌ
yQx��88�~��o�n��&������5(磑�f�������>a�x�6ce���D$X_�����U��(�W�� 2����g�����W�zuy�S�T�$`��IrG�N�]��1uSc���mzf�Mdre��=2k�u���{��'XtB{$/w'��I��<U�	�J$�BR�� ��꒿��d�zCd0�I!�j��ѫ.��3�M�ͧ`O+Tg咘�Y뵝!X�A����S;u�Z^�����$ξ����/��"�8�@{0�d"J�-O���܇�v��#kt�J�I��5M22vɒxI�#؝r���'6U��9+�P����<s�H	�B���~wY���#�ᚢw<IS�# �b�{�x�<H�-_����9��������������W������	���ko��w���[͡m�s���	"z`z���M���v�-���ڃ��5�0͹	�t��*x{k�j����$nI�����v��Qg6��Є}��X��~)���nW�ݰ��]����'WD8�<?��ٹg�uz�L�Sz �rذ���t���(/i+K�zxI0u����faaN�_mgWRo����Gv������%�T��p�0���!m�F?�?�*/��C��)�������9�$�@!�8S5hʤ�+	�.돃"d�,��3'�ᰠC΂ft�$Ȯ�95�)7�/��'���s� (! ��`�&���\�|��znX�1S5h��w�J���E�v��B$=���u�xdS
Xrn
p��!�����J8$��$�$Q�@AR��=��L��>\H6�W�4�����~g\�dg2�P�K��ĥG��?'R�V
`�>������B0�*cX���e*�4Տ���C��^Q����+H,��$��<Q➺�����ԚaЂ ���C&��&�Xȫ�1���`�8��	,��r1J����0T�gf�kW���,���{�No�Cd�2�|w�6��֥_���T�.--������]�oHǒ����$�<��}lu��D�n��9+�:���߷�ݚ*�g�yƎ���e����#�Dx4܏��C�s�{G���$+d ��$S¶qcgG�}Y��rY�--*��������y�𦵾���9P���sb-bY���#�(d�j!�@�@Ue���#�dZ|9�q1�ڊ��N3+T1���ű�3�¹����/��cN���^���?����N}�ۃ�5�)�������`�͖
�7���9�do�O&��^k({B7�6W�rwg[�\��Tjb�}ڞ��ia!��=�Mn=��1<�����߲��Ic�h�����
 �`|��Rk`ԅ�W�F���W	�
Dr�S�8}Q>���v��s��	����O�6d�߱;��ڥ�?�������#�b���5,�I�@�T0�NE��H��RE�!&�7�E�;�U�lg�v��E����نb R�O��	 �sE�O�pIXؘ�zE@%�ɸ�G?���أU������c��� j���Lh�轂<��O��`�S��<��VO1�v��lspNak��=�lԳF�}�-�n��&��ԛt�#IA�C(�u��;V�~���z^����|�c��ڧ�B;`��=��9�Q�3P	$>fN�"��/�{zi���E�&X��_1ؒ��|N�T�Ť��f)�&���D���>��F�!I����-�-��(1B� ��}��
w�I�|A���D0v-U�R��@G� �,c	%���٬�`�' n�X���:���>QU���h�V,2F�-76��vMϓ��|�-�,Z6��������j�J��A��K�^(HZC"[¢C��D�3��?�>Ӑg���=u�醃�v�/�]ĒjE8B�O.��!Zr-ZkHGc�Fv�Κ���[�ش�4�އ���6[��\6̌f$����b^s����r���	�l<�Y���#G��Ғ|����l�і�Θ���åI�?��H�(x��Q��Ѧ+٢��VlfvQFCǖ�셧V~�W��ڏ�pa����'l�������m~��]`U�_�4@A��M"4ă���5�����vݶv�6��3�L�C�G��,�����8jǏ�r�(oR$������QY'v�W���m���� mQ/�Em~��F���	9i��y��c�J2AX�����˦���v���̣u-�]!ps��	��B_�پ�_�a��(����T~��1I0(�3�Q��Vc��XL²�g�@�̯%!�C6f�	������}�������Ȇ�f�r��T`|Q�C����sPq���0�/@a|��*B�l�W.�Q�zZ�6B�z����4�[T�AU$jn�����R,���H	�$Le^W{?��6f	Tr�	������0;H1\��2�5�����x�u�-՗ ������!��A�80��FT �YNg�IzK�j�V�$�rb�oGk�4A���݃���E�i4�dA(�4����w�6=LؐX�?���Jє�[#x�������U��>�NEݯt��0� ,�8|^�P*!��6����\�������v��$�ʬ���@+q���C˲�$���@���ݺu�z��$����/.��P�7���k"���ST�A��U���&%52� )Zc�T���C�<q☽���ҧ�̕KE���p�"ic&u���q-Rz8��P��{x4�f�c7nݱKW�ڃǛBX�$��7���\^A�����l�A&���%��U�l���g��`�Ν��7�cl0L��@"C��_�>�i���0�Kg@�y/�ꕧ�����KU{���?�7~���p����O$���w�}��i��֌��p�Pb���k��h��� �N�R��i�ީ�Í�5:i��eɢ~װ�N����*3'm�h�(@<�TK2ψ�V�Z���l�Z�?�f��j� ��#+5N��]�*���� ��bE��j��Lz�{H%$��\Z�٥�[Y��驲�Q���H�������"R<XߴZ��,�K�,�v9��e��shiHM Z	����)K�_*ft�g2y+�+�<��d*"��
a�)�Fdq��h��,v�v�h�M� �TK��2{����#	P¡�$�Sp&>.L$��!8;MOϑ������^�Ϭ�����3���3l�~I<�ܻV7ë��KX�������.ɜ����?��:�Q���I�#%
��E�E���������U�;2�-�W1WT��^1��t!���@�a��X�t%�W�$��Χ��]���6=����	��+�h��}AU�i�3O��EUHz�NTŽG"!A�B&��ґ ���{�8~� Ċ^k�w.��v�偈v�VEMB���2l$����ԟ|���~���D��y�1�����'OU����I9�`mm�+	�dcyy�
����/�U$�ɘ���L����$:�S���d�T���A�p>#9F#��6,��QD!d#;3�dPR;[���~MD�ǍE���ow��Ʀ�[h���,Tc�
w�i����ԵN��l�y-٤Hz�L�IO�����Nً/=k�ϟ�������v�a��l謯�6��s�h��%�����)�NSn��Ȗ�\=��`u�d/�_��_��Ǿ�Å��~��v2�$��;ߪ���j�۶!�@r�Rt�,h��Np���5�۪2�Mi𒉜L�7k��9���t�k���r�D��\�l(!c`Uz�/�b��P`������Fd�RiiQ���ᒘ8��CF�A��7^Mި�iɡ=h��5�6�pڝ]�*��z�gΜ��}F�w��m���mk7{
�$��跢��uI�O��=�R�nBF���d��8%O��kS����rْ%�D!�x0Ҍ��g�]�g��1�c�#?�"�(��<�[���!)8��S�Y�����+A��0��	�h�%6��$y�s_���u�cJ3~>�I�8��~�Nj[�z��UX�4�7Jǜ����W�g��ajc�A�>�-� �
4����bM��^��=�T���O�G��4�:ẕZz��Q���A�U�F��`�m&f�T�m�5�g�f�Ø5$�XX�B���!"|�,ቋI�@yy�+�f�(I�1����ӢZ�g$o�$��@��`3I( PAU�S�&fl>ڰ.�+X}����׀��L􌜐z��;�{̜����T	#!'�����عs�l~aVH�|ͳ	��!*^~�m<ڔ��L>�k�t��>�p �*��#���?Z&"~��!)	3���;��<���AD��\����N�d�ў��9�XX�2���M_bKNV����9�Ԑ�v��@�	�ם1�_m��e��+��
rhV���+�Cr������W>��]�����&FCk5zBeh�3I!w�.�ڝ;w����g}�9�m���-�:'�L�J�Pٖ
vd�l/�_��_��k?����U�D����w����z�f�gM�P��u�I��/e����ö�ݹn�����Ma�^�fk`�[={�5�T����AOF}�a�ry4���h���>W�v���flL��5��>���u��a���<�d�ꅪ��!�t�q���||T��a�c��*F�4;7m=�I��pͤ��_�W_}U��+׬Yo�?;�"dCQ�ɩ��{}�\s��%����u!���#�67[�~�a�\B�6-2�|��H����3A�bB���H�}��4�T��~,TiHC%*�6$z�a~��F�C��`��/�~2�D�*�RZɉW����%x��@ �PDr��0�6���R���=���ocYz�X4�JFcin@@" m��*��It��d�R�'h3%��W�'pF?�%�Y��Z�G �����,��-~_�?��� �:������IВ�2��fRR5I����A�T�d��<%<��v���hb��Me��LjT!9U�C�'68ȃ�vŲN����t�L[?��Fr����CBBKIˈA���NOZ�8gWD��feM�m�Ǭ�����+��[N��,��gqa�Ξ=���T��k�WEVحk��֭;v��a;y�Ξ���KW���X>L��5|�E"I���I��p#��4.�p�*�r"��4��T�Ru�
e7��Q,i�_��f]p>�\��ȡ|�;�=S	$�����є�&/0��P����[<�5��}��r�#_��HN@�^x�y���`"3h�i&q�Ӱ\��iIԀ�9���`�u)7�/pݸ��V(�ٹe�	�.��ŧ�W���/�pa����'l�����^���S�����bW�,�_F�Qv;�~�}p�=�hf^*��U�X�m��H�Nc(��v;��m�kY6=�~wۚ�-�5����Y�2c�����X�����ϰ�(��݉u{D_���]J36����L[6�諂~b�R����T0�( ��%cN'�k�|�����}+S�j�_���y&�UU�fz9g �L�E���$R�,?�g{�����]�-{u�������^y�k�E*�IQB�D&rL��ι���� �>=	 @�8�9䠧��v�����_�ˬ�7<;5^���%�|�jaorF;���    IDAT22&	!<Q��Q���\��!�ML�,�epB)�xݚ���y'D��TBR�NP��\�ZIb�7���B$I�.O���d��VD
�X�o���&%��rUy���.��7S:hΛ�M�j�Ȫ�e����k�;V��+���n�]4E��
�����[۝v�RSjD��NASuH���N�.Eb Eh�)��H�N��E�y=�Y�>�͗��;Ĥ�aE6]�9W��lVV�}����1±��Sk����'����TmX�C�g�F��ű�a�*#
�ڴ�sZ�ڰ�A��@8h _,�m��x���T't��Q�x��'�>(�iKs��8�U�2i�]�v�؅jU�q�w5Í"	B�w�c������艀�,X���o�
Ԛ;�J�\�t������Ǐ����޾n]��𰼶dg�\o�R�w��*�C��		��(����J�"%�4Oa7M"�[�ƔegKlF��
�!�3&f�u;��xvu�HLb��hNS�G��-�tB�2ZC?�J��F�?%�vS6�U�ē����ح�Q+���q��L���jl�\���t�W��!���:�x)p6�o���id�1�,"�l�Gƅ7��Rp���_H��=�K�A*I
�k�(n_��O����gߟ��ޞ���غ���_�V�:SI&Ku���̛���,��<v��Ί�Vc��$Q(�Ȗ[���O ",�l6�P��F7�)��ʥ4:NAG �D�����2��� 7�z��c}�|�(l̓j͒NQN��r��چx��F<M�9kUx]-	/&M���R��SnX4C�e)�%/�Ύ����#v:�w��$�� B��P�rW¿����Y�z��2����iIry!'~jy3��0Lt�(.!�Vk,F#xe� �+�*�@���C���g���`��������2��<�3mv��YP9��E��F�S,?��߁��*؞�	���-;,e���/vdU����_v6z�������S(���U|�9s���N׼b���9��m����-@�&%�"§��"��Y�ӑ�=�	�����]��v�>mH�]t��'�ms���*�s^gKs��2�3	�P	Aj��fz�b/���?r
�ֳ�������h�Xe
��C��4ֶ}T׉����v�P�:޶D_t�5۾�|~�&FYp��H�x�ܺu+FF͡�g�z�@PB,]y,W�,^�~��5]����%�g4�>ܨ×�r��|\��Hf�3��I�b*���s��$�,�3�xӀf����}��ټV�)�C(��E~t&E{�8���C
�����"t�*!ʮ6�Ų%�խ҆dmi/�0�%b�&��	j��9���J�yޯ��z���\Cu�W�B�
D�h���� q�$�7_4��p&�*�E�j��9sj��+�Kju�:f7�[�1�Δ�nu-��6��/f1%׆0:���n��q���,D�	������fa�˟�����;[�]���r�O#�ۇ*m����u��@��"@6dn
f����r�����S= �pd���)��s#�"3��X,��X����!X͒�H3�%��p��+��	\&Ox��Z�YX=H${���Q��rӊ���s��3� !���&RI?f��.����`�9>9����'��h���w��PMZ���}6#0	%H�=3�r�$���0=e���IevV+��OK�cg�v@w��+�Q�PpN��B$������8�:Ch�J����Q~�I��zl� ���^=r�u$)�6d�a����E��М���"G�$7�È�͛�cb��Z�h��i��"І��'h�b���[{3��� YG��t���Β��wu��t����&��.TO����I�<��h�E�!�0��:ŉ��-�%�ŨKm��:�O:�޳�׽�:s��k ILZc�{�����
9�8F�j̡:L�����aG@5;��۝��Fz�p�"����/��w�~�9$�C�z9��.�-�G�(��Mi�	7R�ՆƥxK�$��a�Q�vlێ���������R�	���<,��n�c)e�I�'��O!#�����󈑾K���W,��xJ���ߏ�Aɢ^�tRIΑ���Z�ov�[�n�hk�e�d�ȅ�5Ǒ�0�[�b9�����^c��F��;��qF^z0�,���Ur A�bG�4���xVb�%�}�Q�I���ʫ��X*@�U��*��L����SȦ�&����rNK(�ݹ �</#����ij���W�E������(ZnQ�$
��_�ٸA*D�*��� K�`7�C�U*��W�.��C	u������:�y�����i�7�c�����u�ls�:�� Z�"L�+9�2<?����d��2ٴt{}�惟��3CK[hX������aT�������
c�[�TRK(�ĜE��09�P/dQ)L�\�B�Tn9�H{z�J��gkrӊ�������T��	���e���v�t':�]��$4B�`���΀��,�^�"�F�:ْ�+�!����f!�	$�.z%�3�d��,#�VN��d/��ɮ���Bv`d O�>]�l,ZЇ�������N�$�E���R�J$p�2���V涄�tț��^�ga;&�yX�！��V��(��t�YZ#����|G#ޔ�-��M��ϛ��Fº�%si��"�:5�Z,x
~���R;��d�ZR�R��f)�T{~*Y���4%��c](R����������TM
��HMT�ª�NʔC�F���pDi�t�2S0���*=(	]mF�*���Ն����7�-1?�6QK���>�/;%��b*3�\���א�'�����N�gY%��X��ߔ�dG����?������![x��W86�9E�5+py�	�d	=|gO�QkO�/��N�d?
�:�
�̙i��f�m�:�4�b�B�9�@����/�-["����m۶ahhH�}3��t��RI�ۦ��p��oQ��%]�X`	����y �]�I��7sbU��f.�h؈ǃ�����튃\�d�
��W ;h[�n���̌�1��,����gE��2!���i�#I�4+ȗ��f�csS��3CCH�Q$�:���2+ɖ��R.	<�k���b�A��H&�5*�=���&v$�}%��D��c^��pf$'�uFG��J��=����ρ�6��G8O�=Q�]��ҏ~잧������M���6N�:�����������Ye%����'7iH���5�l˕2�IqG�5w����TɅrM��i����@��G1?ۤ��dv�����͖��Zj��(WXli��٪}=s��P*6Q�0��d9����"��\�Hz�n�<,_>a�߉�S� nl�|���������$��y�n��9�*��i�]ؖ��dPF�qt���Oz;�8����As}���n�i��F4څhl��\���@����������4��b�T�jJv�@��FW� �"�e�T�"5$���J|�3bf�4��a��Np��车|��������Q֒
�Q��ܸT�!�E�(��*v
��L'�@�[�h�5�!Y9�;�Xۖ�RP�;lkH�qش�&�g��4ܰ�:.E�����NҏD�9d%98ݦaf�C7;�e�؂��49�2�K'a�B 0$�f���)����+sb�wAd�����d0�ʠ���șC+ȜUT�s�����q&�͓EQLQ,5��fUL�^��Ȧ�χ�f*}>���H����O^I�!�йy�ͽ3�e���cH��|�".�:%��%O��p��w&�&3��,�e�t�(���gW\���C�ң#����P�6��,Z��/�d�W^yE��\^����u��c�x�嗹�I�i�L��>�v�JCm �����.�F�O*��x�n�3z:�kM��~��y!�MNҰC��,2?�l�;�]�7�+������=L���V�\��l��dH~"�A�bU�rA-8�#��^�f	� �6'�V~VbCK{J�#V�nW@�R)��L�8q�·`�����ҙI�9�}��}��Q�GR�xxP�2Q9�㚒\�C49C��f�İvQ�K���t��rl]6�/-m�^�l4VT�ե�z��6[A9���ZF��F���Dz\`�����O���AOT�+�BFP���@�<z]je��*YCn*�o0�J]��WG��C��EKS�<IB�5:�x儧H.��ݔx��X��wܶ�3:�у��Tz
����å˓x�ͽ8{fH�Gh�VF��w�0��ʊ±���2@�lź*����S��Bw�{����@�N���\N��@j8���9]X�|���3���D�b>/�?�+u�$:H��H1a�FHP�M9/V�7��/z>a��Wi����:Sz�Y57on��ѥh��Ɛ��k��Ѻ�N�F$���E	���UX��I:�>�:^�2�",%sf53lä��r��.�=�{��T��]~$,���wI�Dc���g��U,�:�(�͙�:��W�@���4;�em���}:ߗ���|�6[u�cӓ�y��dg#EՑEq�gX �d!�K�EKĒH/�I�3m'%9D�Jeg� ґ��6�fк�{JC�Iƾ"��*8�����yHy��%�y��kH��K�[¿B��҃�=OV�gJ�$�I�  ����Ξ��j	y�P�܅K�r�ĩ��,q��F/#A9��ZRsfv���m:"A%�y
�gϞ��˗c���^�u9ܴ��NŰl�b�v�H�ꫯ�����Y�>�ɊX��p���>£܇��G�t��w��Ƭ�ZfU���������$qM�ݸHP'�Z���0�����V����M1E�n![����4N�A>OT)$kN��l���B��a?�P�LI�UD:���O�X�qT�m�������P�Ѵ��U����#"����į<HRI#Q B.J3,(��3�^D"1D~��a����̳���&H��}0�O����b�8�Z.m����F���c�SΜ���5.NbׁS���EA�_p��"`��DT���7(�p<	�f�H��Ġ����@�X�ɋ���dmN�ӢE#|LS�F��X�v֯Y(��� �(�����Yȫ�l���g�8�d�Q@��KH�)n1��sd"�0�E��|$��N3J����Lx�p+��wnw�;
��*2\�;�8�²��t�L4�YL�;9N 	\��x�@ p��\�z�g=^�y_��֠�V3j6�^�4=?ږe�L�mkn��b�����tM7mâ���lY4wӶ\F˶m]�M7��鵚���ntӶm�jZF�l�����8��^�9�N�?g���i��kv���А��^[b��t��u]7Z-��4�0KȌV���n��0,�����n��[��ٶ�[6E6�vٶ��4M�5��̏5ڋ:8����V�0��U��J��l����KT�e�����-n�-!�H���lw�r0p�y_�"G��ֱ�J^3�����S9$(���!z�`za]+�Xu�����t����>&匿GNSl<T	�UYh�i�/�E,����p`�gb��$Ni�[N@y��k8Y�'����M�!=6"rv��P-âe+p��Il۱�B�bU6�wwۨ�Y�^�!�����-���c+C�����ѣb��/ɹ�m)3�fH�ߑ���2%W|�WC<J�J�|^�?_u�K����#an_��֮@w�jM��j�$c"n�"g�^9�(3����I]�|Ot�.F�y	��AY�'��$DC˰P�4p�Ro�����;�uE8j�B���b�JRl{Z�nW�.T(Q���4�#L�YH�mc!o���z�9�%��1ǖ�A'ዟ���M��x�zT>�d��k�����d#�űb^�7?�ܽO��zs3���F��78<<���ÿ8:2���/k<Ο�=3``(��{���s���T���l�B�`�	�@rd���!�*�]b,B8����ca�6�L�Ã�ON��!�FCC��4����V�fq:~��YK[�_�k�7�|��o~c3�='����M�X��]a���}�(�7M!Zp�BV&	<������	f�z��a�#]c2H ��
;[�le�yi
�հr�,�׋\vS�a��$���J�\H������}�ҥo^���A},�Sx�:q�t�4=�F��L�XT�b�h���6C�,�����V�e����h�j���].��l6��mۆ�e隦Y��j�<1���-��ې����<��i���T_-]7�e�-b��[���u�z�˟���-��]-Z-90���VK�m��l5�iz5`Z�Q����tA���2شݦ����i�v7ZZ+��:Ep^�2��H���;w-O�e��u����-�i���Ms5MS�2pϴ��W�4M��W���,�ú4��|�a���a�ݞ-�SRLf�K��tL-J,�*�v��\�/]B��.�<!���ڀ+o��S��7�"=U�$	�,���DMؼU��	x2�ptĢuB�S)&�4��寰��{P�j�T�!��:�ȇ�����.Z�|�7y&$|2�Qx���kd���޻o���n$c~X���%,R�b�BSy:��E.�P
B����˳��8�����D8,S��b��#�f��&JU�c�>;���2,�Jkh4��\�8g�H�*�y��UZ]a��G3�
���b�Vi �д.m>EA�>�-95��{�s�z.)�#	G�c�@�F$g�Ļ�b���X9��O=��_���{ݜ����Ǐ;�'�l��Ŷ+5��a���"Rl
N�e^����2�qH2���̈4x�|"3&�5Ǚ��*�W�5Q)W��1�)���e�~ЏDW'�.��eKf���I�r�){;v(�7hx���ؿ�m1���̔t��&3���+�fn,���[�XB͒[�	��S��$�j%��iT*�4L^�*���S�*
ڪW�ɸ`n?ғ#���������9��WΚ�}�������Xbl�O�8�D"F�P��.]*$���d��ш�u=�-�˱J��u�\#�B.W���f�i����zm�[2�$�e������@��4e#d�J��_(���lv���D<�̈́�F%X��\<pr��x�2���v����?���g/��E�]k���T��ћY�@�X�퐥�K*6�IQ�T��'�@YJ{F�B���&/�G�=�g��[8��_��H�d�*�Ͳ ��������ᎵX8o� t(Q	a��&39d�u!�ۣg<=����� k���4e4��:]���Zy�B� ����8p��5zV���@�\���H�Z��"�4Ju���A#*W��<�$�q�m�Zd^+�dI��Ywۦ����5�Ȇ,z�/%H�0�"	J'՘�!(|l8�D(@���ܾ�Z0s�?q�C�;��پ{��۳�䩳��X��:�ܶ�H+�/a4ü9� �z;���F�!y�J_���-%����ʣ��EY�0y3p����Q<x�)�wx�Luc�m˱r�lx=&<o6M "#bP�E�H�������#a�u��#�5�BR4���z)�.7�����<'���Ɣ��$!nz��߹Jل�r�D6_B:���4/L��̝�/^��d�;=�߼��;�|�.���2�W�ǏM'b�r+U(���Թs��%:��G�����o���shڴ<����ZM�g�^�#A��!	S:2-���Yrw�t򢍩�)(9C/hZ��	�#sfՎtJ�W��Q���$$A��8�3a�t��i<����a��>���xt�]������z.Wl��Z����5�7m�V�Qt�|c����2&�۴�-_�QNTK�5�rey�R]W��"�_�������Tk�04Vƾ�g�I7�ĥ����2�#W�Ex�������w��W�Ԏ�g���������,_�+2�q�ԘB�g7���Yv�O@T�/r4cP�7�hLbE�0��Ê�3�=��;ￚk�f=�*�\�C���86:��ͺkV�Xî�G�G�z�RI�mڰ��2v�#ur�#��Խ�g'�CJ��ܐ��:Ul�$5��;Q�R�    IDAT2<����Bn��}!�`��a��~��<�%ֆ�mG��,i��o��Ǐ��@o_
wޱ
�v!���6����3� ��H7(
o���ޕ�t�7�ئ��"�)�����i5�`�"��9�������ksf���%K�\�Y���^��{������Ǟ���;�&�{�~;z-�>�a4l�m̴�ۊ�L�2�h��s��d�fSF�Tv,-�Z�4�o���bbC�&ۤ;ZP
<M��dF�� ���lF�ْ1	x���M\�p�߸\z���
^����MS�,�%;�K{{{+ײ����|6���l�^[�dWi������<��?��ᢐ��rG-8��pA�W�˜O01K�h��ғ�����E�z{%�^�L�"BG�.��?,P7�]:�1[X%#)�1���Nx�P�x"��j���%��H0`n_/�ϛ����w�������[��rAN?������]'.\B<���5�����B����5�3E"���V�"̓]����Kje�K�\%6����h�wB!׀�@s�n�mX��K�m�G�!�a�����pN:]�k�o��S���zRx����M����� B�=oBFeї�L_����@�6$ϘuŴ��g�Jż̛��8/t�0(U��x�Y�����-]���+}�/���^���/^�m����p8����K�|>+�Ha���h\����B�=A�*5���^欱��|1�JEg�C䋉c����B~�1�t�P$" h@��u���铓���!T<^03�x($�Q�>x�߿x��w��V���u���ȹ�~qhl�7�;h��0&ŶPTNy�Si隈���E�[ɵ6�� �L8�{�)�"C��ϙ�P��X��ŒΖ
���W��Q�\�"6V���T���|I��,�m-�?��?7~ތ�d��D�`Fω�ߴ�.�u?�-YlGFF��?ܽ��O�D�3��V/��Ӟz�	P�J1��Ѕ��D�)Z��!8'���dC?b1���nU!Ǚt^�m6C�S7|�8�ް��t��n!ȹ��w7�1A���^{c+N��$�3e<p'f�H �7��2��Ŗ]9�u�8���� e��]6Vu�n1��g����Rqe�Y�t��RE�G�,�?������{�W��L��pv��ާ'''���<4��xiPؾ���>NHŀ�N]�EZ<d+njr�fI��Po5��!DFp�%J��B![P�⨥�U�D,)��D��''M"S������lSS˂D��G"�8��}�G{l�߿�K�mǶ�9?|�O9�=7���}'-,�y�H�Б
����F��]�|��xA��V�UjV�X��IԞڇ�5N��t��'�;wbG�.�V�LGw�>��lN�K�iH|^>.��
i���TW�@�Zӂ۶��DF�}����sݮ��o�b+����~o�ί��0��TkV/���F��lYd9�$|,
�+k�\[	�➊!c�婌Ŗ]����i"Ue" �j۪ػ�02�*�U��7>��:�ؒH�$J�^^hlÃɉ����95 ���	�w�z,Y0.�D����������<!�IjJ�U�VY	�Ŭ2�P��dr�BM^Y�n�ip�x��O޾x񼷮�B�~��
�
+p��q��Щ	���ti �c�"�sS�b�P�*i�L��}E���t���D�]�K@��ӭ+�&>6�ɉyG��渹\Nrlɶ?b�d�ЙH"��Vm ��R]��N��~��%�::�)��������?��=�ܹ��^�W�x�K�F~i|���m���V4���.4U!rr6ʝ��NK�9�K���Hz|̹%�I��Q���&9a+�pD�\�E���S}�l���p���S,
y�$>��%%fDb��t�~2�� i!�����4M��} �n�b;|)w�w�������Б����K��0|�(Cv�����b
�IE���'�bQ*�[[��DGF0&.��F]�[�z־k�Le�(V���Bx�Cbޜ�*�n]�>��.~@&��RlϞ�_ ��$�k����m#N)�P{�[K)��J���3�T$��hP+�v�L�r��R�"��zC��mC�O$	�l�,=��Ǟ����:�~	�+p�+�c۫�ʚ��d�Y���˴�B�.�V9P�\;�H��N�Q�n^����O< �1T���rA�$v���$_�ja�v��8��b���y;&�Ɍ&ш����D��aFw�4�>���wܱ�{W������>����#�/gCo���ѷ�	�_�X(�r�G����9%��|�.ѦLBb��	axF��	mD3cYHZ3z��C�'������	�g�g�ݎO�4�י{��li���ϫ�� �(,z�V��n�3gN�=.���[��NL���~w��GOF��	�^�7O[E�D
�__��A��%�Vή�f�KN��T�sAv����bK�;���
�nۋ�t]�u"�q<�if�&��F�>�,-����c|��o��g��I��v��+�J������W^���xjS|
.Xݨ�R	o.�DC �
C�Yh���EԪMq�ἪX�fPa�������;�W��N��h��[S����rS�Tjbg*���U&;O:'�����@ɼ��gL���)�S��jn��|�T)p�Q�*�d)�p��( ���/�	��a�W�<Լ�&����W������-���~��k��Xޯ}���?|�ѭ��ay�ӎ��@y���̸���}�Hu$EJE��ɩ�h�ň�A��OR��>k�߲��AmW�r�ĸ��P�����>�U��B���}�ӕ�)\�D";I���=ntœ0kuX�f��O}"z3��j�-[lm�����o�}�����f�j��1�N�ζw�C�b�)�u�;��2����ӛ�tf㕹^�Z���B�P��-�11ZA������6`��>)�~�`	Q�L�m	����q��(6oރ�Y�UB�Ѓ��M�C{8,�a�.Wke�GXly���Z):�=���U9M��R���XB�r�l�J]�;؍3��T*c��y�^|�S+���~��
܊+04tq��M�G��,p�XS��Z�x��dQ$��e��B4��mj2-�d"����ф8J�����eť�$E �'8�-�1�J��n��e�� ���u�dq��Y���D�P44$cq�k��g�]�lٲ7�s�ގ����}�s�����5���!w�l尟/L��[�{=�n��#�	�m��R�C\���b>�&&��,�,����bPb�.�j.���Ï�����Kt�{���t�b��PH�m�T,�ΰ�f��矋ߌu���q+[㥗�yl��cK��.�X�D��̈6�tM''����N:C'�5UX�99�$*�pI���!0�}J4��l۷�Cz�a\�*�~&��L���6����	���Il޼c�94�e��^|�������uǧ8��`+�I�pir�-���R������W���g�+��ސ6!�b��/���6UA�P�sv<��{����W�V]�m[�v���3�8�-��V�d���x3O�E�HŠ��#Huv�O��ˌ��nm�>￀/(�~�ٜ��0��	z��ł�,���Q�'q��D�'���#���}�1Cq2�&�^�C���zj��U��n�������}�y�A�.��\*J�fSf�S�,�VU<�a�n#p���7��F�Z�@��}n�	��
C f��9����e����&�'�W�U.�`�bW�r��:��~��-�X�h>f�'bQ�-�'��Ii�ef�}����X����l��|�o���d+�/mt	���G.w�;E�'�#���*��
Ơ`��uxAH1��5Y�:���9�|'3y��f3�MFć6ރ%�g��|�k��R��2l�.g�u�~Nȉ��;��>tRQ)����Xl	�脹��F"������@<^m�'_0z�s^j��Ų\�<���R^@�U1�0g���=���U�j/���M�����������>�{�v����J�ru&L�!=�+�H�э�-��#�(��)�\��a�1��[M3V��5hK��e��SR�Y$:~sXM��m3��{,��K��B�:�	̙=!�O��\}ᅏ.\����#�>�ږ�_s�~)�4��Ix��AT�Si�����\	�U��ք�Ƀ;VA	u�x� Ie�4�iӽ�W�E�&�,�c��8p1	c�"��h�%�M��S�����C�ڰ?�h8$��Ŗ�p���<����rͼߏ�e�-���կ�<���d��^�.�&!Ɯ�V%m-}4U"o.�����IGب���iY"�23�5Tf�,UD���鏅Rń�J�]�`B:�
�M�*�fˍ��v�:���c ��/�G6m@"FRTMY��-���ar�*�bo��=~��kKڳ^Ȓ��P3![�E넾���;o��7�~��M��E5���+�ϽǏm��CG���y�	4jn�5��[�����ʈk�e	����Y�G�{b���Œ[z{�c��\{||<Y�����ٍ���O�'Vf�?�m�R�&	O*X�hY�Q�N�m�(�"�P�4�~��1�'33��#){�G�����?��f�c�|���;��y�A�.D�Qt�]�yY���b�L��S��#?Sθ�����ܣ�ш[�{ ^�Se#�|l���������`��ǵZ�f�f�Z���\H����0��l W(H��s�e�
��sy��2�lԧ��������ݿ�V.��?}���>qz~0���+���VI/�8xg�R�^����v{vx��=0�3���5]��ͦ�V5o+���V+��:��b[��ԔZ�$�6=���=��X(�0"�����j��"�Ug�Bn3y�ncd��=���q)�3fD��Cw�#��LK8�x�H��$|n��f�D���[���>�nV A*��|>���1!lp�D*>!-����+�?��?��O|��tN���x?V�����ȑ���la���n�*M)�,���[�[��<���]�p�˳f������{]/��Ҫ�O}��s���3����$�;n��4/J}�#-8��,$�q��:��	yמy���-�a��F���c��[w���{�T� �#恟�(&3�(��҂O�H��*���B^��ю�"�0�Ʉ�sĵ�R�U$�1!)�\����#�Ͻ#��d_�*�lv�չ�܋cc���zJ�
��H�� X)�!�G_��׏�x\����tg{#.
>�����Ǐ?5'
b��5W�-���b��*�Ű�������ڙL&/j�F1���P($s�̦b���byٽD0x�T%�$�Hc��c(t�l=q?��,�����B64��h=f��Z�c��#��b��܅���:%;u�}a$��t�̹P�!#!%|�GSL�Dg:�����SF�X Y����LȌ�J�q͟�蛏?��*v�F]��3��^�#o���o�<�����k6ju�hl���D��
1
�8�Q��e+��ڳ��׺�_�O���7d�̅I!��k�ot��.�,4,R���$��e��02��T"I�n�駟��x��k}M���G����wv����t�+��'�k�9E6�e��[��C[�G��)�!��#�,�f���IS�4DCat�:s���D8��K�,�����[948�����G�G�Qm��d�&&#Z� �@�hT2�k�r����|/��~��-���r����r��������[+�˔�p����*���.]��X����.����yS�����'h���f�d34<�=���R�o�Wă��Y�y���w��b���N�U����v�9���,���� 6>|z�hTT�I"Ì�>$�1a��*6dCh��B���uB!�a*,K�P��� ��<����L��:�MMA}����y_����<}��0����UW`��W���c����R�2M�I��Z�ôta��"�0�,^��>��/�����?��_8r�į�3Yaʊ ����GQPg�r	��b�n��cQ�.�X�;Յ�=5�~��7���`��n�{��,�SY�HF�͢��Jy!<IC�)ubS!�t��XQ���Vlg#AA��u$�3g��Y�f�ܺիw\�Z�:u�����;y���$ш��*gۺK\�Ȑ���b��$�J�8���ϥ��w܌�ݲ�vd�бm����]�a��c��0x!�x�nx�.��R�E-���u1��/��J�˕��	��R���}�[Rl	EiA����)9��J��XB��6�ǪI��wb���M)��>z/��X��5�tw���CI$E�"���9���Dx����	E𾠐�ƇQ.�b;62$?�����k`�%���?�µ����W�V[�];��{�O�ٯ�l�"sr�z���Ծ+�+����ӫ׬�x��g��믿|s�ַΜ=��h!ζ[���ǚ�(�P������b;96�d<��3gѢ���s�͜?���X���w~~�[�~u�����L!�P�D~���[#�H �U�K��uk|��C��16��$�.Y�����+V���C��}G�����̖���-SE
�F�%�AOyf�K�<�l׵�����l�e���{Ν�x�C�ښU+��Jw[�U�����|O$������}fl|��n�����ĩ�g�{�A�J.�k�����5�?�����z�(��6�����ؾ�-��r‒Lz����ˉ��B�`��4����+���ڶ=#�ڔѴ����"���@��EzbD�~�����se,]��ˏ<�����zL���
�*+�־W~sp��o��J�*�9�2�5%��'.F�m�/]�?��_^�{����Ë_�[��X��G!QL
k��,dJ}¡�J�1t�Ǚł(;[�6:bqv���|��+���]���޹��:y���ܲ�&�g�BGL�iU��0�C�^V*	]80��+W���
� ��Hѣ�ݦ���*˗.{r���߽����s��[wl�:82c�e�^��|^7�� R�!H1O��ˎ?������z?~�.���];�]�t���p���j������\2��[�����������f�����ⱱQ�8y;w�uef����m�VbFoѐGR̋e�$ۑa΄��F&A*;�;�Dҋ�=�H}���)���l%RkKTܔ@6��9��Db����.E�(�xǐ������Sl�,(�-aْ��C�����?6���
���<����֪
��I��U=ސt��` ����w�u��'���m޼9��+�\�py N���2RS*lZ�z�(=J�bQEp$��,�+�2*���:�	��ܸ���ׯ߰�z_������[�ǁ��_�޶��H[���Gg�@Ӭ�4g,=�R�"����S�ļl]��� �A�_t�$y6ku�BA,_��?=��S�|�^ůny��:���Fu��R��"���HI�%jP�eǞ���=W�o�cn�b;ܿs��K�._�y�n��0::c�9�LM�����p��<EK�Rw:��
g�FCC�x��)l߶Ŝ�L��Č����I������Rf�Y+o8ہ˓ضm��\Z�=a<��#3ҡ����4 e�N�EWA��|���Vy��تt��22�q��b|bDd@f]͜$�l٪�޴��Y���^��8��_:�%�;U�9n!�WIYl��n�Vԓ�<��?�3�o���������{G<���X�m�_�򋅞m[n�ζT,�Z*
Y�Ŗ���}���>��7o���Aϳ{�/8u�S�����t3f�D*ΈQ����ؖ�U؆W�1���+���V�h)���`X6R�ܳ���-��>��}c�w���Sj�Ieh���.)�,j����'^|a��^���F��ܱ���A�h�|�	t��"�iu�:���C���b*_,��=�U���A�9s[��E.��D�G�{��A���*s�v��ْ�X�/�a�=(���4̛ߍg>�aă~a�@@qx<����Fl'a���~T���`*�_Td��    IDAT�Z�eӸ|�&&G%2�R�\)�K�.��Gy�'�gM�vzn�8���ap��o��@�l�D��7IbT���Y�^����#7�=���~�ؑ�o/�HK�Ѹ21b�ʑNЯR��=��j����7Hܪ�Й�Rl���G�ܰ���~��=x�t�����K�%���0>5�R�&��a)��8�2ٶd�S#�?L1���M��}��>����s�߈��?_��7Μ;�
I�l�Ồ���d?-��^�ԧ���X𡡡�[��:584��Q|�'��J�hbr���D��<��k���+r��[�`�S��1���������]ȤM�eJpE�x��MX�pZ�:<�]�Z��VC�C��ضu/J�2��b�<����%t����)WAnɒmۓ��5l��6�0Zz��j�h:�6�h/Y\�xc�^��J��E,_��O~�#?{#��9�W����}�K�C�~�r�b��L��R�)v�#,:HYX�p����'��7����~����GV�x�𣳫K�.�X٩r�IT�r<�ݖ�Ff���~��R.��c�/[����z}?�yv����C'N=�e��N4���'0rˮK��d.-ŖV�F�%���͚�K���#��^?b� �O㑍-Y�p�U+B~��|}���صk���b�c5-q�JDb�Ffg[*��_���3�q�\�4�d��]'�GƐ�㑍��MÐ����k�G���k�����O���?���ȥrã������X��*��6<p7͟�Հ� <nZ�5�d�E��q��8�nٍJ�
L�q�2��O�+{�L&��u�2��_r�]���~��w���%�
N6͚��i.�,kU��xĶ�t1�ϋB.���"������	i
%,]��?>���~�z�d�g�W�VX��������S��.�X�cj�!�V��$͜���/���'_��&���/|�螽{W���DБ��c��`Ifn��̿��%����["��Jv�>��G�ϙ󃵨7��عk�+GϜy|��C��@�x#7�2<��s�(�	���-C��İ�ٔP~�=1��f>�3���3�X�z�S=���o�kݶ�Ͽ����q8�b�2I��Eg�b˙m�X�x�����7b��//ں{�)��T�n؀޾��.i,^,�?�L���{ȗ���B������d��W���^�귤�fKM�����u+�d^?<�-�'���Ƽ�T���Z8w~۶�A�\�f�q�}k�O=�x0(�Q,�s��������\.�AM�~h�m��f����wX��tCO�}��91�P�*����˗���l������1��8��7�hp�̿"�˗Fn4ɰaڂ6��vvv������{n�{��/~��[�+�� q3�����)ώ�]!�l��g8[�d�X��=��S,�����]:p�^��lwn~���s�v�;��-e���V�ox1���'���2Ŀ���B�ES�AEö�A�+t̝3k�ҥK_\�b���}/����+;v��B(_g�,�a����Tȧ��Ӧ׻��yv�۶o;108���.�}���߃@�����������H$:_}/�/��<;11�z�Y�0��B4���z���-$g������l�
"�$˒��l-4��.���Ѭ1�����_|a_/N���_�ř.]ߛHt����f۶����o��͟��ŋ��/&���2�`ي՟����v-�=����W�؁o�֥����ޝ~��<��^ѫ���I�\��&������+�_��f����^}���O�=�dsB�d!et�,�c�U[�)1tD�8:����T+��3����$rSY�c��+V\7S�j>�-[^�y�셻w��6ҹ�z��JxQ.d�+����u��͢�%�V���.�^I)�8��D�D�` ��N���~�0�-�z��|�#٫yM��1���o�v���GC���0���2D��G��r���/<��4�)��[��|��Ъ�{���+��Ć;�#���%U�Y�crb�`4��L,�x-�����&_��
��Ѳ�"�Q��k+�Pm�g��^�s�t����g�m���m�д���z��(��}����`%>��S����`�9`��D:}��4�s��Z^�m��f��#c##:6:*d-���f�b[(c��՟۰��-�=����W�������ȹ?-�K�T8��HG�-���0<���c�mk~�ɏ<���}�/��گ�����ӄ�����hm�A��Բn圸Ѩ��a8T�6ͯJ�21w�L��P���Gn_�b�[��ڮ��7o~e��K���<p�&f̜��T ����'�|�(b���2�e�T#�^v�]�1��g����X"]4�/�]��+W�z��c���ߺ}����pۇ ��t{şyFW�8Y���I�R����n�����vt�����^BwO
�߁X4�2!)�E�Vo�q$��`�s�joʞ��'럚LO���TN��[���L���19��7��&�Q��^ܶv9��I���ѽb�&����YB�a���a�8~�"M/rX�~���#��������������?4>>���+�_���r5������Y�L�FGG?6����DF�e�S�4��ª�k��������}���M�����o������a64�ccY�-.�Mz�6ivQB"�D$�s��{�X�n�5;͵��رc]_�[{F�&fCQ��Up+u�Ȋ��܋&�S��R���|n��ԥ�Ι94��������M��vۛ7�sص��WN\x|��#8����>��
�Y���R^�l�ZC.�uۖ���L."S9��D�\B*GOW
�xt���'f_�{�������T��
��s���Зꖀ�l&W~����������n��޲�v``xÎ��v�F��}�:��>xt�P^:�4����\^��t�];4�S�o_�m�bfA6_�D�X��JŊ���.�lݬ��#��t���=�r̫�"�Ս�n_�y�pi�,�իe5�V�z�NO��/����Z�a�<��F̙5�-�m����v��������~�۝���������a�57���j�G''&~��J��l[��b�A��pc���?�d��?����sM��q.����c��^�!��`tt�� b�Ζ	=D}�y�]0��?�싿�^ދm���~�o�t���?����&Q��Q,W@ so����˽����D�Oeq�ZRl�Y)��Ѓ�h�ڵ����u�?�}��_;qi�ѭ��ƅ�*z�fa^oV� �2�/da�&l�%Ŗ�#紤mҙ��	�egGB���|�b	�pH���S���oÂ��������ٻ�ѱ��{S�KF4�4����{�l#�͖����b{���{��#��ܻo���(f�����"����,��^��>蚎�����8ʕZ���n��=���n�k��Ъ���Z�V+���j�K�ULiѨ��U]WNLf�xc����6!\��!љº;Wa�����k�|[c��fJx��9?v�B�R�D��#������Jv�r�V�<x�g��B����02�X��Tw��=��m��P(Ge�RI�zca��z�R��t�R��lV��FS�))ٶ-ej�b�j��Y�`�5̓o�g5��+p�W�������إ�3�:8?�(H� �Q���:Lآo��/ؘ�x�o<���x���[����;�����QW���ᒮ�.R�|�RY�2w�ߺ�5��y�^�#Q�b��l���I�y���nZg�y�+o�ش��I���9���JV�n61���is_sC��������
H�����U�T'��l�0gf?����˳O��u�OMN��ڹ�+�N�������&>�O��̲��wfO��e1����=]�0���y<����{��Nb��YX�v5.�D0�F��S J�"����H�`�@�9I��� �6ZR'P���!�XL
i�,�bILfJx�;;1>I���xw޵Kv���MC�Yl��o䁋�:9�f�)<Y��{��}���"�L^�e�b�#C1^�Ԫ1E���ex
>`o����`YfW�l�i��yj�TA��b����hHG��C��������r՚O̟��o��O?��
|�W������ѱ�?g�M�rLLaZ���5#���j�(�bƴ��f*�����~aݲ{/��7x����/���塡w��O�VC2�)�Q�d'�j	 ��0�q�����4~��V\��&ZM��w2�e���c�޻lٲ�N��a������q����N``����1�;�e\��da��BKږ���I�;̶-e0c��m�|NH�^�!��K�-��M��h$�\����`�ș����{?GĀc�2a6[�ǎ�c�����B6Wߴ��x<���u���g.lڱ}���t�kV.��c������;]]Nc�ܛN�+OD�0���A��uKE�*݆��A�ސPv)ht�F����{[�cp8�ZSG��[���E�pUxu�c��<�R2TE�f����9'��`��8�A����ғ�f'��L&�UƦL��N�,�<ER7[��d���$՛Rh	���9#B�	��� �{�W��x�M ���1�׹������?���r%L�P7q���(]��z	>�[
 ��Z�^�G�͙�ծ�ԞD��HzN:�ht��^�F�f����V���J�O��k��%dܴl�O�x��a|lB�E2����p&+���+�~�G�\&��3���V[�M�i�m;^�Ι�#w8�KcuF�CotST���-��`�4.Y�f�y��^]io9C��,�܇Kż\�K�,�����5so2�,|��{hh(yq��#�G�>s���G�ryA�*��D��6	����i��Q��b._���R��}���{��[�؞>};���)T��Յ��������1_��W[�|�Z6�]z'�Eׂ�d��7 ��,aֱx�غ� m�&BO�'�L�������PŊ�xG7�w=�.��U��:�K�-'�r��r���<:�f݄�U��EI<��Q*�01>�Z�,�Z6�v���7�?/^��'7'�*��mπ�Պ�NXh���xUl�U$�GZ�ė,_������/�=]e�?4�7y�~忎O�U�r�t	�̆!Ŗ{��fp~[����w� ��z�`0�	�Be������4�!˴�9o�l��L�%Ș����Wk5��8�䁞�,�����:��⣮��D�Xtg��J�⾳�፫-Zt�f,ߖm�~�����݇N��}��pf�z>�Q�%4A�%UM�d���&E���&�Vlk1��P2=��^�l�c�?��HmŢ[�8G4�B�J5Ѩ7掏�dpxtU�X��'�"��lZ
��ڻ�����>����Ǟ�۱�؉�qqB�n^���E�*���P����GE�V�JP�V�TQ�� ^mR0	�4�	�!΃�1��g������[k�;7�a<�վ�5��{�=����[�o}=��d%0mm^�w�`�Tk���~ۭ�l�`����g���w�|v���Ԍ}{w�2]�U�*qI���\,G�"�G����^N8�B��ST�(
�*G���5�>��r\�FG��>C'N5h�m�2<Aw�u]w�n�F)i�K�=xz�	i~�M���=y��0�P%4���C7_MSm!�%4=}�ʢGC�5��0<L�Cüp�	C��C�FÀx�k� l��i
x�#���g9�숮��߸����������8���?wf������L�sK	��%5�9%	J<!�}�.Y���T��@+	Ҹ�gh��T��P�q�96��Ҍ8�K�%W���:�q{�@E����� d��hƘ��x���pI|m�F1b����\}�e��*}�y��gOM~���Og2ڵ�bڷ{3�E�*��
�Q�(lq���o8����t3|���2��qn���arbG�8��Z���-k{nn��ACWhdt����n��8/HW#�қ�� L1�6��ew�~��k�M{��=�����/,���6�:9F�22��
�Dy����\��R_In(' ү"9(�|��j(Fz	3aѢVi����L���4x{�FW]{�x�>ں��`���#d�B�tv�E?~��>5G�V�	�Rھ�F�#U�ƒv�z�� ���رh�GX�fxh-���� Aɂ����^�.�B*L�Q1~���4�jvi�]y��y�5X��Ǐ��ߜ]���v����V��� ���N��@�!ơϣ�J8�M��M�ƱË���FT����7�:�Z���#���2wZҪ�H�^��~��b�À�_d����������������+�����>tbvᮇ�������/��6k/�h�FrV$����n��@�B�z�.�n�שˌ�Y9D�l�0d�#B� �{8b#�uY��pZ`�0���l^�-:�7��-�u�� r֦��{�׽��-�v���� ��sss��?����={S��4�$Mn�P��!�3"��M�V�%><�f���(�5��<=c|�S+ ����b<��cʩF����3m�9ۡnY��ݻ���Ў�q
�V�"���BөSg��ggi~v�L���H@�.����L�A��g�SN?W��kr��1#����`!"(L@e���0"&~���@aS7�i~n�tX���yׇo� ��߂���Z�'���gN��)X�YJ�3��=��nU� �x�G,�������c ���$〣�-;��ý��'�=^�N� ���o�uУ�~/�� �5IHI./5{o|���߿����x���|��������Ћ�{���t�ދ�h#�U��
�QG��p0d6�L0�R\��̔s����@�@��
�D0~�EʒJSp�"cCAje�e����7�rx ��3<�jk1ö�s����#���[n�urjjjս�km�lO���3ǿ~���p������W)�`�����-��͂�>���4�r����G�e�P�`k��$ZD�>�B��P�V�hv�MgZ��GFij�m�:FcuQ ��)uL!jR�U�7�^^��!E;��h����`�1��5�`���
� }e\�Ml�e+Ԇ��#��p �� �M�Ann��.6�_��ۮ�����B����H8��/}i�1�� �Ǽ��@�
i�
����c��qM8䬊$<	 	������J�oE�,4���N=����O;0E�&{Q��}���EtI
���)�haa�8|�}7\s��'^�>��C��_<�Б���LF�쾄�?����9�hG,Ʉ9:5
�R�[ɣ�V"N�;�e[، �,?�{Kx>�����!�XC3�2��A�\CB��`3ͭG�,$vVP�P%�2�V*Upmʻ�w�O#��ʙ���6��|n~�`�"}���)�DV� /I�p��F�n� ZD����h�B�ܰ�L;|�PI��s7��5J(��E��ҹnNii�h�@
pbvf���S��qޔ�f��QIM�h(.i��x0����|F� .X�������.�� v!��N6?K��o����ל.o��43�@��_����z�G��#�/���x�_|��5n�r��
���%X�=qƵ̀1��P���N�1Hc��(�G�5ҊA�(���BH��<�V��s����H&
�g��E���UW���Iiz����[�~���_�v��|��GO�����#Gi���}�죛��K:kPL��̨����� z嚭M�fh_���
�S+�4��\c�GH�r�`�nq9������`���9���A)��Z��n~~Ѽ��;'w�ܹ�Q��Ξ>��fs�3�n�Wt��(v
�~�2R`�� w��	+�AԒ���`-ᕕ�9h9jD
����o�!AmI���Y���U���甤�YS,h�5܃�c�m��*L� �i�UECUM�=kHw0+)W;����Aċ\jA s�,k,�����
'�$ ��2������[''��"�ʍ�P�}x�R,,����=A�لhLһH��8�E٣ ���Ƕ\9"�Hi  �IDATsNkYH� �b2MP��A*�Eul]����^N2g�lM��QȈU(�j���L/<�"���x�o�ֻ_��~>�;r���O͟�����ť����K��EUզ���G���  ��e]{�!d�X��'ס�����sbA�<�B&}:��, �l����+n���ëę��8S*�P�(�B���b~���l�i�U�c�_|n���,y��bW%%9�# N���V�9p8��&l[���-�lצ2�Ԡ�*$r�&DA��S�T�=��.4HK5��Â�4#mb��T�� _�{#��툾r=�H��ʴKqH���.@T�{F��CP�B�ͦRd�J�Vf��P.=�.7�zkȨAmEj�5��-[?�o���ʏ���[`C[��������/Z�GZ��B��2%a���f0N��>�=�jHR|�Ij���`�)g�?�3�����e���������.�� ���!�(�R�47�@�>�"Ml���ݰ�����}`qzqi��G����wҍWJNa����B8f
�� �B�"$���S�W��KP���M�BC}�EFJz:b'2f%�}"I�K�"5�@�l�@W9�87�����C������)]o��?�W���}z�ūgN����,jpE�P|�&V,�0� �C�ʵ|���L�����67F�F `� �KM�P��
 V���P'�Rty��e�B��xhJ1�V��K�XH�jD!@�g%�ڎ�L�Lכ���Ny��-�x�跕:O@IW���-��x�D$#���o�kx�?�ܵ힭×̮����-��,p��}��<���T	����[� �1RPJ�d�CZ�Q#FH���FFwwK�`2`�H�P�Kp�"(��������=�/p�y�s�s�|���5��UP�PKm�0)��. �l�f�
��n,�f 0��afǳ��Vo,TA����[�����9�|���V����9��9��?U���xL`��7{�@��+��l�*Eq��z�zu��Vr5��Hi��O��?�>W��(u��=�Lw�b���O'���^��K�|��HK�Y,����Nl�a2̟�_�t%t�~��U���p�ʦ)2��� :��)��B���_G�=�`�J�2�q$.��O�o��E�O�\�x���ѻF���x@ґ!�	��`�p�#^΄~�HB$TT����
�R�5�rDy�e�N��qL��(U ��ܧ�
uɣ7��\
uqh��D����3JUt�����O�[�p�H1���4ፗw6��1�߆,�B`�L�o!�gJ��n_����}.������hS�3��Y;wA�i��JW���>A�$~���:�-<�~Pƪh�0⾢Ədsq�0k�Qھu�P�Fx�1��vԌH���$�+xw�=��)>U�,�Q-d`��ZMW�X�!�}�`I$뽑C��n5Ek��D�!��FF�&#�sW����J(��,�����t&۹�։���'4�Ɲd�^��}������`���i�{��Y+a����H ���L�[ca[�H����������b���X��<�n�'y��V��R��T .����1��@�N�u���>i�;�z����X{���L'��Yb��=0���.�#�V���|v:��X#���p ,f��@����`k-�S���q2^�8��r/��~�Ct�S�᱾A������L�SRS��REv�\���ٜ�E�yY��ؤ��������=��n�q�y�.(T![�G���m���0���椢^����ORm٫�3����fg[�Vb�����C�	c�T2b>.A|��E���Ӟ,�۷�m������v�
�1؎�9����]ka;z�G�#Q+:ʲ�Ee�F��!�o}�??[yǆ����]�&�u4��Q�n-��o� ���Ӟ��A7A��T�D�2ڋ8��c��~v���|�l����JS���aɷæ�rѣ�s:�^�T���S�/�~rD�����W{*ve3.���b	#n�?��޼A�Ї���=�⢣���3�,&�l��`�^mb,��d{A��-����W�|P/��;Z5���E���|.�
x���������$�&gw`�}ڿ��~&7��c�H��OK��rS��,�L��rI�����7�5�vFY����rcc�]�K0�Q��:�<����ڡ�:���x@�����`�W�K��.'��"]��qΗ�;{��BV����Z(~���<�7�r�oۥ��AA�)^�wD���+��\��(�$ǩ�ye~p�n���ě���|0d�t�U���-��%l��u��hȈ^�.N+�S'��
�-�j��W;����w��{��ϦO-��~/��}Bҿ ɰ���2����j�ǒ��%��t���w]��A�ɯ��.�� ,$�aH�A��g�&��L2���L� �	�v�{/g��u~�D�!�kZt��BͰ�����T���������B.�,0={������O���3��s�v��.�ƨKl	e��B9�&_)!�oA	 �O5"�^��OD ���&H����?R��q�iz۩�u��zh��,����{8Z��Ia�lN�������;�8G��\��O���>���8���X�F:�2��y!D^5��]�� ��r�sR%�uK_.<�֬|�(T�_���e��(v�1B�
�w��A��ڷ'�,�_��}\��b��(r7�m�KP�?���g��瀤VÌë�q${���ׅ��{	�II�^V�r/	x���@{�K ���'���~�V4I[~���1QT��wd����C�c�r�����-rD�9&�'��@~׌���(�L�(Aj`I�ǖR@���o(�=���3�?��2����BP'S���q�J6��}b�u<�C�"@𡐳<KK�M�Q%���~��h�6',�-��d8�3�lTBcDSw-��o4��C���3q@�C�	��/��-}&��I8K}�N��ԿP#����݊��N�����[��j(��[��3��xiU+Cx$��05�p�t�v�=.Tg/{�~����g�7�xЍ�4I6��S4�z�#�{��.���eliJN�빙m�)��u��#5{w�9�������3�kcs���{��� 7J"�l�غ��������� VM.Dt��)+��5�T�9�]��+)�v�1��;�v��F}D �SmA%׵�f*v28��2k���X����"W�h��ݭ���
g�@���ܟBH<�t@_�b59n3�jHB'�i�.p��1l���9�w��o�$�{�?� �P�*��g�]-��?��.P�s�e��eC}���Z�#���ݺ�����'��^qbgm���}t��Ѥ��9��3�.�"u�$�Տ?������vP�y��>۱jq1���*�|��|2����f��e1��N�E�a���}~���۠���(.�)�6�M[�e�%�tN��gu[��GҌ�t(�#T1�mҖ��"�����y��^B{�Q�7/������*����y�����5n"3!���B�h��n
.�#Y���=m�'
 f)-F#���8���&<�d'�aP>�������@@��=�����������MP�ۇ��N��>�swΥWJ����m]3��x�Íp�~�v*Y��߷=Ô)I c�)I�=�>RwZcs��D }$}X�!{O�zo	�j�#�v[�M��2URJ��-Z��6������+�iQ������6"&w��bHt�6�+J��%d;.�	QԒ�`0�~#�1��i��<V�V%(KP�gA�����Y����N�&Q\��o�{��c�B�1]) m#�Iy�oǢ�	��d�X?��Ȯ��/b2��`�d�IFq���k���A<Z�t��F�X���������a?|{HCr��g��*t\�lw���Z{@:����H�6��ubm�3+��F����z��a(��0��9�m��ظ�4i������<Jai�����E�GÞ�s�So�8���:%��Ώ��2N��#�7lRy����.&1�<ZD���'�zR9	&�M�s��{�i�F|�U���j��
W���%�Bx1g��ce�I�{�m��*Z�Dh8�5��{J�0B��W�y�����@F�.H@s�1�l���IG�/!�%�a���������O5X���^֝Y@�F�Ʒ���n�	��f�]H���4�L	.�b����^GA^������2]���|�b��;�I���QD�[�����7��/ഒ��� �γ��A����X\JJ�-��%��=�+f�G�L�uqM4G�<Z�w;���.��� t,���]7�]q��kN�T�J�kD5��F/CM�C>��fL���4r[9#C�ilt]�؎^���1�{�ˣ�O�W	�m� d���g�>=�`�YT6����V�
�L��2�M�#"�u�[B*!k�\ % 6��o(l�x�ޗ�'_�d����vM�[~6�1����WJ�%8��*v�A���弹F�72�;��x��lQfs09�; e+-/V���DL7��r���H��}�����9���3�	|6����#��8s���g���?w'#���s��O�V�ɐ���ٽVZo��]�n��R��E6����>B:�E�Y�w?�,RZ�Us�����Uc����D�j� Y���bˢ9gЄ���,�D.<y�EC��7g�WY4��}3�fEL��Ӌl��G�%�#�+�:.W�裂�K4?!GgGy��s�O�S����ԟ�f�Bu)�1
X�Ss��i��3b�Z���:��B1�P���N)*������՜�y�}#�K��f��\��)�A�p�r4��:=�R\��/y�˙������n��ľ�24�x��}3&�����usn�{�u��ع;�eĪ6����+I��~@V����_�+C�K�SH�Z���
߭���vs��-?N�kr�v*�_�RqX�g$��F�d��!��w_<�7r�bfc���>i^����l�>0i#�b�s�C��'匫�����\Hs%))	�bd�:��2#�z���j@�w/��������M"��:�`rȾ_�#`Ue���`O�����kˣ���6ۜ�u�Շ��ŀ��[Ǔo?������Svl�rc����9(Y��'���7'/&��Հ� ��9�\#��셼h5w��4+�52N�u����1?�������v/N@T��]Gi�BR�Ք�����͒�+C2��X�=DmLݐ�$@V_M2�i�5�y=	�Q�E�@k�$���~묹��K�E$�a^�V�1T�	��,Bδ�M1˴a(��,���s�\k\�3ҧ��
��ed}0����R������������xm��0"s��֣='��A����9ܯ��:��'�(�$n_�`ya���̷O��]�~Ӈ���֎L�?_�_�|Es�9(z?�-8��ݐt���J.>
ܲ�oHT+��Yw9ˑ:��<�|����<*e��Qk�G8��8Ғي	�ӷ��cBG��<E������5������r���hH�D0�y���^��n��NM�hwM��M���r�Ƽ}�٨Q[��U�,��L'_r-c%8���ݤH���-�8E�>(zz�U�_n���H��t���X��B����K��D��G�X
#�!��x�66������BMӝ�{��~�]ѝ��[����_΢?�D�y�fӢ�_QH�����sǣ�����C���E�� ��_Mh�z�F��#��/���R���C}��v#�g�Oh��A�U��PK   �u�X�j�� 7q /   images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngT|	8����R�$tN��J��%������&���-J�"KB�}(�JY��6c�!��G�I��g����*�5��y��~��}?zz[_���&&&6�׍��X?01�9||'�F_|:�����a�t����_�7-���>R��ku41�<�y�������=����%GW����������U&&!&��&���Kָ�ލ�)�N�>,ie�8z�ｰ�Q�>k���]��cr�c���e�kw1Cο�n�r�<��oL���G?[p��?t���7F��J ���}��)�u�������T���%�RtHQI�Ly��G"ovf�}��-��4(pTr�}�һYH�j$�A]�`��eE;�	��݅'�b%�ĦF�lt/�DP�����d�����sՍ�s���-�����/y �ȻX��e�g�П>�J��=H�m,T�k��kT]�t�K�H�`����k��R3�2�Y��O_�{��X��&�T���]U��+�^v�����sq0��96]�D�,潕�d ����6h�8��Z����-1�r���vsѱ��b0彄c�@��)��|�,Q����:��0�����o�t-O?�1�rͮĤ^h����#���M���@�g�p�F�(�J����pd��k=r��{ �zq��-MN[�]E�>Ò��!{��y,��3<��i8^j	G)�P���ʉ!!��[W�JՖ��N�����b���4|���N���.kK��t'w���$-���##��0ֽo��A�k��K�^/�u�w',T��}�E�	�i	��O� {���+m���.�����bmic��w��1��c+ۋay��؜=��H����:�޽[Y�^ȥ ����m�m�%{B��|F��=\��뚞vW[���.��h����?}n���ג+�KE��[l@ af� ��2_���X2�	�n����O�~����Ql���)v'A;1��7�}�Q&��&��#�d�^J�%�wxϩ�"Co���^3��ٮc�$�4b�K���#���e��ʴ�'z����f����7��f.o)��4�;�%]�'H��ĳXRˮ4�������3�q�H"��H�b�þ���BG����;���
��b(�}��De�0$��H��G��j �� ��C�*��X1��D�eE�@���]�,�m��*�$�QB�g�X�g@@���b�q����j�x�˂��ـM��BXep �r�t�ʉI���s�n6H��Xi�"I0��|,#�&��t4�/&wͲ��$�����Ǉ��T�iB�f)s����9�"��'����wB@#1�[�H�=�Ge���y���m��_7�:������ �����A�`a�O�eMS~����&��&^�N쀩ϻ�oʴ�D������$�(�Ѻ�CbC��<�t����G28�H䱹C�xK����� ��	���tw5��D�b<�ˏ����"_a�B� ��B��#�D����ŭ�~�~B�`�@|)�Y��r�L&gIϕw�57	��Z��(F��<W�g?�L���fz���؀g�]P�S��í"Fw�JLF%*R}ߤv�'��L@ri�%|\ǖ�pb�d$�i k�w1�T�Y*�,u*^��v����6C<	b0!ּ�"`K���7��C����Mlh$q��|�@�%6-"�k�OF�&�~�Mԙ]_�0Ҟ�Ԝձ�5���ќ���8vT��d��a%�8�r��3�N�Q\�Z�1:��N�䆸�B*�qx��P����t�@5?��_�0��*9�{R8�q�A����u��E�c�bJ��z�J��D�N�S.t����B�@�/�� �gh�[ [�H�����;R���So''�GqK[���51ӦT�/�����W�*4�k5���_a{H��^�(u��:!
-���Ƴ[
�,��Ä	�~X�aQu�~��p{<��S����*���詎?�A�-}ۯ4}	�S��bJq��pCLJLL�+)財E������[LA��VJ���D�Yb��������ހF{����A{d���������@������_��mQ�C�ԃ2$L��
�FZ��F���~M��q#�ā����׎�7�}�ۨ�ѕ�Q77�����mV�+�ҵqҡ����z��J�Oco�i\�ߐ��{�U�>�l��|��o��!t����������B8v "����>��jF��F]k�\�ʐf�c��1_����ٱ���K��I|���NG��1�JLn��/'�*�ˡ��5�-ڀ0r2={�,��)C����/$��v��^��������ׯ�n��x�����خ���kKۓ�N�Q͙�B��a�˟�CN>�z�Dlh\�C���nJ(Q��������6*:JNV�<g����5�Ԯ�x&�\� J�j�jltۿ��RS[�@"\k���+�Z�]i���GG��i�VG����s�V,a��F%�U˒0Bsl�!���U!;��Ш$����J����e��z�e'$�ܠP�U�Zo��jb��j�|��������9��N<#s������Yt�����B���҃Z�&�!,�(�<uj�c�8���b�ɦ���'���<:::87WXS#�@ԕ���/�?���N�����~jnǽX;f��}���	���Z�*	iދk�}��/w�r�T�����q�q%&JU/�M^��x��u�b\����QфYÄ����n���S鹈Y�Lmm-�P&+mث���x�-h�n/7%�!d(Og�q(v=��E��<AAL�ړ7�L/	v~`rw
~��ؽ
7ӵHaS-z���#�b�C�cw�%
�U�c���!����&�y EnH�GE�=�*�AA�^�sjR ��u\�0p��,E�b�v�-C���������������~�U��B���?ںfDd3��yz�*��k�QY��oPgnk�2o�	�)^k�f���:;�=�����?����	1�����];OI��5x\���������yډ��(�1ٶߔ:����,� �t�Q=|��ufu��a��]�L��/����jj9?~x�%�A��o�q�DL��=��Z�x_W�8'Q�2f	���`I��P����?��8����d#7�A�?nA �x�E���!el�%�4`/�����:�!���uZ���������ٶ�Д������D��z��g�4�l����q�Wf��?��bd�~�?؞�`��!;>В�l�1EX��`㤱��.pr>b�.�3ҵ�w�1���L^�e�h�t/�>����xezi8����KHioo��U�|09̤�T%>p�l�xk��S�#�ѣe�cɴ�6j�5+�����6k1��l!����D[�#+����=��O������C�Ш��}Lk��dMˆ�#�X���q��FN����9�Q��I���k-i�q$���1�s�q��%���2��\�6*�Z��.�%$@=�r޽����x��1_�@#�����..z�P! ��"�q,kD ��
���{��_�q_g�1�����S�@B����ܛ�Ǐ;�ʪ�Wt޸���!
ҧut(��9Kc8e7��3���Z)�f��;v��iK�{�4=�'zY����Kr��6��ntaI��c�y��?��Ib��acK�=z8��x/}^^^K+h��]S/S��7$��iIr�zE��5z����Ծ�h{���ݲZ�gDR��Ӹ1�?U33�3	����J����9���5���[��K$�Or����:�������Ȼ��H�U/�G�h'g�[ ��i�3�!,W�B�ϔ8�"�h4�=�y�c����o�)�F��fb r,��>��F�M�>�V�C�Ղ�"һ��؁��.�����8��9��h�hGק����9ɛ�2␋@�@��|\wղ�9ğH	1��l@e���Je��.~���{��)�2O;��x��n��9uXY����k��ɽ.���#��5�IW�+x!��,IP��߭׬�|�TC��~�-�а=�J/萭��7^�?^VF��F^Ώ�Y@9d@�S80�j[����̇�3H��mi*�Á�氄����/��k�t6�:¦+���k@q3����[R��:�����<=udd@�%I��ef�|DM�ۚ¹�R��TDSSȣ8���'��IR[��E�6�m����0M?����%�^�XX�#Lл<�ƔRP����O;8P��7��������m��t���w�l�^(��X�U�?)V.��@�U�c=ӊޛ��Г�I�e���m���:ꅎ�O����p�ף��*/�mi�tm�w���nsљ��OY�������x����F%��N�tw;� ��B��X8���>��K���j̵��M*Ss����+��%�.B*�3��	NM��E�C������|a������n�����m ߙ
��N���u�X�!ݒE��B���]����cZ1�=.1��jnW$�d�����[Ub��du/��(�"(Ky
�n�d8���ŏ?^���9���R-��fk:�q�Az1`3��6��L�Z��XrLa����r٫W����[� ��D��}}}n��Ds����k����R�4��vn��M>�<@}�6�4�"�~�'�z����/��OK��fwl[;G�X�H �"%5���@��K'q�*�z��K_��"�����3�+����N���*��Ռ�I����m���_��to���e;���M��
ViVV �.!110:��Hd��垆#��GC��X���X���^�/���O`2����Φ����*������D4�=��bDDc�-��ì��m����XjK�]i�}@\��=��O���S*�T-#Qu��(6��K����/ȩ_������Q�xߜ!KLbJ
bw���UW�
�����["��6[���x�!|�0gcs��@�/g���.)}��+^Xp��xbg3�9+�?��b[&&fy�r����9m�{刧�m�X�=���f�N������0����P=qw`�&�7S�GAyoO���9�FءBr#�	ai9*�PYY)86�>Y����N�q�]`���3�g)�c������x�n���R��PD��v��A���܁�>�UI	�� ̀,�Hl-{4|�(�c���lA�b���x�M�k�P������)H,,,�So���9�i�}����ـ
�C�g���a����E����vK�G���Ǿ�@�g�!��HW�R:�x7��� �R��sxb::������k�A�8�Z 
;,�ĂM		���_�/��5���i0�����UF6;�/���qAF����J�`H,TH7\�ۃ��d	�C���sU�T�Wj�R�(5�3d��g`p��c1�?Y�|}���E�@aF*j���NCخa;|r �DR���|.������"7�l]%����V3�l�]�M��\k�9��y�1��#���i)��j�%�\�Ç�pU�P��U0_׫�RW`U���#��{��M�FKWShC��f�H�x�_(Q#u�H�;��_~U�K���\" ���	eZ�\��c���0��ᶺ�3Z�����$:������8	T{�Jo��B��
��^����獋���Rrm�4M4S�h$A����
H�����/O4ѹ.:�����?�2�p��;'	+��@�~zU��5��~�r���#�.b'�A�j�>�>y�-����&^x�S*m�ɫ1�p(ۯ�2�l�3�q�o�Be�y�Q���2��ͩv���rpB�v�Y���[l'P��B�C>�{�St��.�-��!g�c�.	���!����73�OW�UlT���_��ڷ�G�ro���*�t�6V��p㳁�V�����-������_B^�MӬ��#�C#u"B�N-z�!�����w�[�0a�9t�r��l�RD��Pi����?|��g{\��WR$&7לJɣ�ベ~�D���\j��I�Ek�	�����FW����O�*⛮�nHnb��8���^��\J}��A�Cz�=q���	k�6��-x�#k[���MV~�F2��t�p��*>V�Ua4�ܮ���0-0���ߛ���ⳁf��0�p��6�mBl��q75c����M�V�o�X�v��hd@y^�U�;��)ymg��4g"m6��\���q4}u��\�V�Y:���l8q��򄲲rW$;��v1|���O"1���J(f;����ߙ�~6��E���ףX4K"��P���Ļ�d�ݫB��^؏��g�0���4a"1M�`{�`�qD5QO���:/����qqq')b]��u���H͉z�.��]�`o�-���ɲ�$�D��v��0�&O\�<K���FPc�G�C�bQY�e#u��Z�)�xq3�a�nue@<�>q$|�V�����]+-��W��a`���;*� ﶉ=��bY62b���geu���3̣�������+�ŋ�b/9WH��h��_���.�>�i�Z�brk�	{��qs%��3zz�;���˿�8} �d_�M4�����%
G� (���� L-��Ѷo���d��O5��b+�����I��֓�H��Q�B!��]�:1�ߟ����~o$�hs�͟uJ1�Yy&&Wr*Ի��Gr�f��D�Ի�:<����_�s�V��p^'�ב=rm3ǂ�cr	��{5o?�F�p�.r�R�@;YW�s[Wy#�T,}�x`��}*��%r�u����o�BWl}��+���%.y�;�ЫFE�;����N���>`7��z�B���K6���^t���y�Y��,i�s���w�r��A��I29dϖ�2'�50��P���< �$/��9F�xT&&�Y*��f�w(oa�' �oKL4z\���"�Y@C�����kmg��݉��:���bT��y�6X7�k���Vɋ�g�|~N{=�P�}f���Gc%q��@[[�+�C�U�k)�p�� �t���$��{7*1$�Q4��������x���+�|Pz\r�m*�>E>�w��X:�d�7i�3`�%�u�~�!k�^�Y7S7�RVL뒩��%�O~X2S �',Y��j1�*[`%��s�n]E}��5�pJ5��)��J��UBg�D�}q�gOA9��jp/���ID�r^<���F�H��l��'�r��+�&�RĿ�'dU�6&'��Y�\L>���NN��k�5�|�C#|��:�d�dP$1��L`~��<�Y��Q�e�NJ::�?y�U�ci>�<�N�u�tQ]c�l��§�3S��"����{��m�c>��ⓔwḑ��|��G�E�+Ĝ�l���(W��$�O��k��?�9:2��Ë�n��Q���!I���}~>'H:���URG[�\~�_�k�������!�	9.��XY= M	�!1y��x!T�L$7�����؛�>�%�k'&uc�����[%�K�~��ȑP�oT�H����1y����z�����'��eJ�4����Ѣ9��`w���7(�,��
��Y�)����k�Z����̍�-9�U����Hd���+�0 �#���`�0x�?k�4��.��I��u��e;}�d$=��u(��YZ@�_�{��kj�Y_9�� �?��o�D^�<J�V�s,v�l����I����Y�"p���u�G���_g�}��FA)�"p�Bi"�W��aX0P_>�����N}W0��kXrwT�)U��D �Ĵ�Ĥ��Gv����О�
��B:<<���kIz,��r����c錪��+��͆ʞ~��o�i4`S��~c�S�.�fj��^:�P<���<��pn[_k��|�U�K��:�(tؤ���b��	���D��p���{Z�p_��+��Q���Q���u�M�D�#��PW �Ĩ�w \V�D���� �c~\B�RA�R�J�YA
��E
�i�^y?d�⶯���A�oҏ�/�C ��.4c��JM�J_��-2�5&�S��T���퇿�ª84�=D_��ec+!�P#���;Os畁FMP�{�ʼ���hVE&���������+���FF��+�M�[�9��`�k6���cY���[�	�>n�c��G��}�ޘ�H![kW0���Oց/rNV�� )�����̐�֠}�*L_���?-���E�~������y�u5�Ǣ��$N��T���m©I�{K[�B��-0���/���{6����@��%�c�6bB�c���Q_�Y�{,���$��+u�gu<@�gǑ�Y�����c �V\c.��Z�7n���}G[�D�}Y	[�������|5�����Z[Ƌ�\E@}�IY�?@�}s��&F�#�r2�H�U��=!����z��򍓗<Eô�N�\�����.��"���Ȕ{�s��L(7�S���ؠ��?�Ϊ70=�u��#T��ЄWTp^���;��b����c�Y��-��	��̠���h�١-{$��KtS�Te���1��$
��:�"�%==l � �F)����J
}�b��_�]��z$�޷LG[��)�� ���{�Ѿ �����o�=N�b�. uۃ��O�k�Cpp'DiQV}���,����Μ	���PH^�G�e5���4N%&N�eY`�M�� ���8*�� ��'{�c�"��7p��$|ڸ&��2�C�C�l�G%��x\~'a& �ݓ c��ߛ�w�B>���x���bv�9��u�����;�^c$x�om�ɍ(?�5�5�@sUUUy�M��gD
���VZB�)���B4 .}���5�4g<�np@���α�@�7^�m������}��κʘD��2���+�u%�E2���A��bA�M���x&��2m�����A16�[P�����+;�]�Hu��u�}BK�t�9Zm5�$���<Q����@W ��_H�)N`���R�Q���	���A�!��f�/<�Ϥ��GEEɪ\�}�z���d�r�W��x]�ɬP^^8%��@��� ��_�| |�t��)�x�z,�^����,���~=�o8��H$Y�ښ�!H��ޕ���,3�~�(��#.>�r}���O�^�5ꗉ���Rfy����.V���p��k.@����γz�֝>Q��ת��jq�F�C�]1�IɅ�.�#�O��+��C�)ej��gR9���ҒS�/-u�;i>-W��[���~��m��
[��BR�ɨ)]�c���j?��N��/���<��Cl��L �����$~W�t�hеV0yc���,�`��i�� �y\4(����q^A<���᮪[WܰߞI�m��Mx�����S�z�Ma���n����<�h>Ax�٩m]�^΅�x!}��)������tB�>[��o���w�)�o+�l8�@^b����Y#��p8�8tŗ;J=S��C����e����Y9�R�>\���י^$'�S�n뀹Sz�nq%s���XW�S��x���(��|?Sc�V�i
����'�'��4����$|����giNO�-�e����f?b����� �=�q�V�����K�q �D�����!�§/��������g���:;|�^�r�p���d�#�2)|\ܪ?�k�p�0}�x�]���i+Pպa;�j�/�n��ST�q�u�iC����ދW��m<�S�8 ��b��ղ����=�I3���u��kYx'zk�#3.�u�E/S����Ew��xxy1�?�w��y9i��d���[e9�lV4����ւ�SMC���U�,�c	�`,!t�d�ᮧػa	�7�r�zU�vv��פ�������t�@��d	�Q��ge
37�d.&��:��GP�����_���������Y���E
���m�k�;�x�r'MS�kn�Qu��A��^�Ҡ��������_�׎��C�[�z43t׺�BeC�9�����yTܗf�ʱD���iy�qBxo-��{��M����+���(�W�M���FkW����Me�>��e.��1C� 3�#Z-�G�Xt2i�F�%C(!W�EX��#j������OK�ǒ?0�7t������H�Chm9bO7�^��
l���9��n&~�����Ŷ�_w=[T9_Rt��D��	�R^^�rQ2�X��c�E"S�d��_����w�r��r��9B�A��D����6�Ča@���"KE�=���F��0]F�,p�y��f���Eݛ����_1��c֏�" -�)ht���9���\X��e��w���Ӝ>������B�*S9p���
��.GL�<�@��=�ֱ�/ҏ2�DbB��n���V�Fd�������?��F�D-|�`q��x��c
���[ȃ2f�i��]ڗ6JNK�]�[|��viuB9pj��)88�21L|L���<U!C}U��Ω���~DI�
9�JZ敻�nk"?i�u�.�k��z�����^ʞ��l*�`�qm/��LK �����7�߄�?{�������������O;��b<����.?@ �^��P' k�ڹ�zF�4j��A4oЏ�t��RZW���!Сx���I�XЬ��,������K����ʆ�7zՋ�V;`{�A� �ݜl?R���H�_f����ـ�2�X�зH֓[��n��6��ϸn ��u��S0�c�WU0��)�n�'E,��]��]W�h��6�;�zh��dT�������,�C��e���lޑS7TBˈ�O�H�g(��j�r�d�?>����r���'���>&�Xi���ݱ@1���o��,*3�ѕl*���G��������p�{�Bd����5��9$	�|!s�u�VU�03�n��|�}�D�ggI�6�_��e���A=>	2���ze�g����ۤ͝����/rS�M��$���V]Y��;ԡviu�:M{^�k�Lc��a��d���1�ßΜ�A'���ڢ�{����$�hB�:�/u���@���� ��O�"}���ݤޒ��|�X��I�ORA敘k�t�^���V�Jo�t�$��Ҭl�L�bA�Jd?���5E�QH���:�����:�Ҝx ��s��øW��ᣔy!���{�U�h��\Z
�O�����OR�����h�,(p���v>S�O�����8z�pU�����hW����B��C9�"�I�w��3\W3��v[�Q���NM��yv���#:LC}�w��v�m��o8�bMB|��+\�e�̲�IS�?
�mZ�� vOf�&��Hj��-=G]���RQݣD�*v�]m�h;�]�IT�;�9�Jt}Lo~����Ӷ|n�z�Hjn��'�<���?�Z���*�wֱ�`����������s��i{�o���Q���9��>�Y$fe�v��������7�_��� *]kL���I_�mh~��k$nk�o��-���@r���o����z�����nb F*�l�S�̘�z����""��	5��5Y��㣣�A������b�]{��9Z|5��=-}&����a������@]����=��M�lt�����{o"������	�+�X�#1Wj�^��KH�P��}���>?!�7�	���f�Ny%Q>F��\@P5{�0?�����ڥ�@�4�d��Y���52�����Zn�;t�7��q�ӯt����x�+��x��kBR�bO�r��p�m��&�j���V���&6��3�,�~��p�OE���@'6�d������˶����έ3zz0�yi99��j�a�\���V�r'2@BR�\&��s?SSS'W׾�9����1����a��
h���)t҅��x{��i�P�؀faW>�^E���[��3��0���;�)�8�o�~7�O��о �|
�����x�l���,g�����P�|�i� �i�u�wR�X�A���!�D������Uν!�G[94_np�@ y�|���0�\5�����Xh���D�܃�uW
]U�߾e�͑�Fp��N���k>O(�y�~-(��ƹ��q���c��i:��#����&�sE~�Ĉz"oP�S��q�Z`m�ͱ�����������"� X.,��Դ`.����j8��Z%.���^�����m�,��\R��X�؝�B������NV���͝O�$U޳�����4��W�83��_ۊ܎�<����ӽ1�#'ǑJ2>Z��<�-����|j��<jG��ER1~C���ڔ�m�Z��>ɂ�[�pQv�1�e�D���Y'W�N��&�_�rq��]Q��u���O?�?�a��/�rlt��
�0��k��z�+Es��
���!JI�A�	���c��qrjj3���n<�@/�==8H_)��&�p�&�V�&��r�������F�
��k�v
�pB��T� �� ӊ��VYxdhp0Yr#������4�����]a�����
LqIIߋ���ѯ��uzKAΜV�j��
�I�����w��9M�
S�$S�,��_1�t.S'������T�֐�^�z������	����������+�[ih��Պ0��j6��2����D��!PM�����g��YS���EXZ�������'�5����gh�,�{�|Ҁ�xW�^��4孤����D_٬�Ԣ{�n
��^zNkZ�ƫf�/RBqY��/�/c�h��z��v�tW�������Q���WRZZ��V�0�ox�����E�֪�a��^�����\Ta�V�G>��Ê��YDݶ�7�U�f����..�箮
���7��j�s��k�z����, w5KNV��4a�l���蓶�'4�1oŻ>T����� ����Q_..Z��?R��{�SsϋSs����TيV�����'�@`��rd��D�\�����S�V�+���2s9U��x��(�����F鹽n/�A��!:FfZ6��s��q�g/*�a��������;(������H�ڔ��F*)5�х&�E{���ZYZ�#�g�_e}���Њ��R�����&{��\F%��z��J9��ck\||}:^@D%F��p��[Ѐ���Hs�����Q��n�ȣ��ô�5���q>���[)�R�#u+/e�q��Dt�>v�Xz���F�}	n���hɴi#,��Ʋy9��C���?�ySW�7�57���1����3�� �<	Xk6���hA0ƇE��DZ��3�0#O� ~Q�8=�_�bt�>�v�ADMM��+Ǟ�[K?�۵���UD� ��9H�k�W}����(���Y�ؠ�����	Y��~z�Y��\�*��"���jԡL#@�;��G�'uΣ�3�S���U������L,,^���a�J��� �����<~|��TS���VF�ݘo�G�ƚ�z���jߣ�	��M`��Z���DJ;��S���+(�U���ߚ9��My#u 1�G���))��UTT���t�X���}��_E��x> �<f�͇of��[���ײ�Fge[| vD$F�'������R��hv�De �u�x�j���j�j�:�boP�.ij��ϴv�B�E�)S�����{L��b?��x�GM+Ԃн�V"�੹{+A�����"�9�Xi�W~�������Z���9e��2@"@�9=��B��$2�}�qYÔǣ�.���yV:�ޟx(�d�.
�nM���(ef�Bh����.,�|�g�ں&��#cK���bqu�V�N��\��gqql 2�@'��[J�u�HN..��<<�I�}��Y���U\�F{�K��[��w�T�܃�s��l]I2O�W$D ������τ�Xmd���ˏX�v�M6t)%WD��]�:���� �ޗ��D�J�5�#w��ź�{�j�S���.�ړ���*�&�u,,F����"y��M|�N�`P���8�a��jPq����-(r�Z���Ļ��TaC##��{�]X�|}�0��;ø��� �<���[*�����<�0%��P���:�S��^�;_��������ȲT�Do����V�ogUz�A[RRn��!�hx4�Q�N�β�Zh]��| �X8��C�moz�{���h����k����������#�éiy'33󟫤�H�4U0��޶���P�|�}Krs�,�M��-��T|�b�U�	��B��.֞��Q�!�l���1���T���eJ�v�>��KL��W?�KH8:9�k��dikk@E��%`<�^�-o��@7T���m����έ~N�C�zQ�X��}�N�Z^����8&&�`��u���p%u��ř�}Ch��2[����o�JJ�'�^���7�#����>y�(��U]���X����1���j+xOD�+@��G!C:�����񹦔���"�NN>�W&$q�W�W'�:;���"��9;��Ղ�=��گ8<�Ijp����N��qJ���H��&$o*4�0Etq1���&A��W�ׂ�N���2�N��漇��_W��U�9Sz�ӧ�~.���ލAl_NE��s!3��R�>��|LaQ!g���HХ}�P7�A���`���1KP�\ �����,�j|־�m_�";����C&�0�����}����T´,"������^7.xF#A@m�@����G2%��
��˯�٨�h���=+�W��x �����%���(y�`UxI�E�[�����h�k�R5XYYY\P̮W��������� l��,�~5�{�_��Ƞ��_�ȠJW����x���]��ߙ�lӥ�k5�,!��Ԥw�j��1-fqU-{;����7�o��,R��ŋ��mT�,�f�Wh�M'V5S������\���MRG��95MGP��*�J�-\��ÁޖII��3�{w�Q�oջ�B)��"-99�6��%PC�b�r�2I�@
��|�@s&�G�/���1O�}!uT��(;��jPD`~��[M��g8�u)��?E�X���yg����y�Pٽ�v����A�T�:b}&���A{mmm�Y�i:�����pXk[G����H���`��� g.���[7�yy������gZ///�e=1�T����|���=�K:���mР�Q0����{�5��.+M��-&�@Rw�݉�)�ʄ���w3�d�DvRO5p���th���Uh�d��xys4��M��\>�f��?<\�]��Y�k�P���i��!�����|�}H��S�x�%��_�~y�M0���Ϯx�zp�8�M�7o�� ��L@?�x`�ϠEx N4�I`|��bȫ :%*E�M=�a��Ӷ
'-�dz����@�H?�����Ĭ�]4@�����V�A{��b|Б�jAw���;io0��x��ҷʩ}��ā��I���=-������;+ |ՙp,B����'Yގ� ���hwu�Q+´P�=�����{rRc�C�j�j+M�X�����T�k]`}>DJ�r
Qo�� 4�?O�'�խ9㶴����n�o@��^s�j{�rek�3�*���eJL�@�=ff153K�f�__��d[��1g���ރ��hW<�,��e��0(��^��_�RR��2��bb���������i��^l�XR�0�ｮv�rY�W
���	����xjb�E�����DJs���vM��S�KG`��h�/�5\Qv�j��UQ�s�W/�&s����$��׵h��ۖ1��j-#ݮ�Cn;n���xA�,?>|�I�~Q��q�$B.Rq�|��~���k({�^i|���)dė����h� ��C}�u�dŚ1��fbfZ�=3��~EC`�����P�3��D{H7Qǲ��u�Г�.��Bh��zj��h�o02�4O�3��pGgg��Ӑ�.Ӡ>�sc
`�.����h��ϾރBͯ<�)���A�*��9�'k�<�rm�:�DҀ�q�ݑ�t�pv(+-��r�$m˝<��m�=�{cN�(�f�/��@��wH`�W)�KI���+p}E�Q���r�j�R=�ԤfL]fpF��ݏ��0�_���ms �4���������1V�z��k~�qm��`�Y[g��R���r�t�E5`���K�9,D��*���n5֌ޤ�`ٝ�u�Α Y�=85�3]\]�%�e�����V谬�tE_�kKkk=�\UF��%@b�44hQ�["��Q�����ktx�#]��D��J%������ft���)'u5��+�|�WRRb��w��k���`W���I�fcph~-�����������MM���"�����&���
9���Pq�E-� vܻ@�}�zj������l�+� 3͝+��;)ꚺ���U ��*��C�
�|�d����B����~CqH�mi0�U^__:S?�+P�c#����s@� X(F��>�_O���$�}T������}/������@ې���lK+��#�5�e���)���^`	+�P��>�ޛ��
�S��\̲��Lo���T��iq��)�� ����X��6���"7�a��,��b�R��?�Z�:|ʹ�e��;)Ė;�ַ͑bc#h�|&�|}}��|��¯�b�\b�/Ў9��EL��צl(�ͣꗁҚ�a��B�7�aU���@ �$�/t�4��K:��m�pv�1���0f.5+�]����w��?�{�PTLl�qD��d��� ~.��:��,m��&?]�P�+t*���ҫ���-qҥ������r(�fߪ�x���_�~��9�Ƒ�h��>>���0>�����i���]Ɯ��ۡ{�������LR
����t��JGlV��#v��*������X@;(c�;вK�2��MǬ�5�Tr�07d����.zP����"eTY	���r$��(ϥ���={�U���>0
��C�/6�QaO?8�[�#�I7j��{U,-ο�V�_{.�lLfu�L�q��ʺ�]D�a�[q]������z�t�������au���e�t��+��jVaTM�"�N;��* �5�@���m���� ����I�WB1Z����|cj�)f�i7DN^�\f������+������冄\5�n�n=���I� ܞ���CQ��R��|�	�$G�s��0q�4��L#��qqq�++�^����ј�*���VS���F������gttל��D`�۽H\����N���H�==�C�%$$�Ӳ�l���N�.E"��|�{���.Ćª�o�;Xc���7&�6li���Ӕz@髀#�vpo(r�>�174�p�2��)j83�tt�4�T&<bH�\UY��`�x��@s�_�ퟙ����q�l� *��ފ�����MQa��Q���8�q5K �P�,��\�s�1����;>�q�/��m\��4�W ihh�'W��w���Ѷdic���������]���oK}��˺
�p�%���H�����+ `�ެr����**� ��/�QӃ��*#�1��5+ P��^c��Xh�Z��V(��߾� 겖^�g�_GT,���|}z�fhS��"�ଘƱGޛ�����t�ɋ�PYi��i]墼��|�b�x�2�<=+Km�4r��D$S��8űwZ]��-�����(�!^C��Յ��r�c�[x�j�C17�]�1䴗��m�/ի� b*���O�u�lG�5v'�9�y�����d�rs�?��t�>�Ӳ��oSX5?b���4���Ǐ�6�~���tn/�5k�;1RNkc"v��fKϝ��ȶ٪7K�,=}d�����W��`����^tIq�m[��>>^���b�X7��m5�R�!�yx�������f!;Z;��SWA*���w��/���ŃSX���͎�>~77��70	��x����B�\��7Z�&B����=��J��aT� TTwU�"��D:�T�U�"�UJ@QpE�ҥ)R#-HJ�H�  RB� B������=�9����3�<ϧ�̝��9���V����i
z� rO�X�~f~���p����w�;���acN�I�������l���ٻ��<��H��cd�����o�ÌM}�����]M��h�۷����X,/\�|c�������>�uwF�7nN/-���I��>@K�ֺ�G��`^�20X�? ���<q����o��"��{/��P֍�:�D�,>����j[X�>}�I0	{`e��|����ۡ�*$IX�ms����ݾ�h�����(erwsb��q���%�m���ħ[�:���6��Hľ�H�������$ܗ���&�]QV��ؑ��V�P*p��w��k�r0�ި�?�w��Ӹ7ο��k�-��4�R�5��:��؃��	Q�����V�N�T��U{ͬ��/���#0^c^f�O��~Ak��uy���a����7e�ȯ����XH7a.J�pG�#g\ϐ��(�����6�����O9:;�J�Wp�5iNO�(ݛ,P"�<Q�����[�%<:.��Y~~����m111	��b^~���y�zx���t�&������X��<Y�7��mT]z�a.*Woz�!����:��`�G)��2O����w9�o��t�J9[�]$v������T�ؕ
����(���`T�|��� ��,z�dR��Vu[\�����n�~���Bi�Ww۴��cR�����DcӀ d��%�O-T"���iP#=h��X�G(Ƚ�p*�4ePZDMi
�ˌi�a$��|���9������X"�%�H��I}3��(�]4>nc�u�gfF�>}  (��O�@)�W���OTA[�eWKJ���
�l��1H��_�!lRâfm�ߤ�پPߑ�6WW�Qw=ټ{~^_]C�� [3�y��֖d��o�"��ȧ��	9<|(E5#��Ln،c�$ew�K�:�,{&t�"��Ǜ6S%��4Zk�fY&�W��x�ӡR��!s��Z��hm$5�$n��A�l]���r��3)p
��|���c��7��u��G,�P5�y�8�Y.�����
�<�b��
@{��| ���+G��}���h� E�
W!k1;`�|�w ;���b���O����_�Ii�Fӗf ����h�������Z��%���[�.��嵬����gT���q^cMː��.$��.�k�v�NN�˂��y��<�j!���y�SJ﫨�
Wr�HL���/�n��M���C�E-yy��Z�4��9�/��'!I�J���r7���\!��V��ޮڊ�YX`K;��@��AN�S�r_/����?�1i�!�9ﷷ/�~T�C??U�F�W}T��VE��Ң�`��Hr���JuH^�{�7�[ec4=K%ư!y���!8{{{��R�;��O�[�c��@.)Oe���{^��fL�I�a��U�&#Eރv3@�h�!0��ɹ��|j���gf"m~[�(�u��S	�9'�h��\d�7T��-�}MH�P]٥�� HBS��d���߂��Fv��?:
�.��rf�K}_.����ގ��xy{;�;Rf�q]�,.�/LT�v@���&�2oqѩ_�{�DE�-|�4楮�jR��h���P�{[w�����I#���Q�*��J��ȍo�7�DiS|���EA�~ve565U�!�1�]V��f����~��2{�Fä,��{<����>B�g��W���v� ��mַE�- ���E�JYȺ �e7����T�.�Tٿ�76.n��#и�mN�!�W럤l��g�y�\Kk��H��|K��wS��2��<�>%.��U����t��p~���J ��յ����70Kg.��ދ4��"0"4��T*�[ӂ��5���0�P��+�R0~s�g˪���8�8��fU�V�p@�.|jM=Y��)N#E*kb"6S�C(ܳ2;w����s��@Y�Cc{����0���HaLt�k�����ꩧ�,HaA� X��_ė���\�IX#��"31��_J��Y�5L.xK�,n7�(��a�\ʮ����0K�������"Wr�Z�����{fU��l��w����D �r��Sp9�����m��V��!^��9�l����OI���4�5��˦���P�����&���d�����_�Z����<G7/TyR����Y�U�ۜ���We��4��(�a������Ll���"�fUQ�E����Ռ#�f�c���w� 1jd��~?(��I�HR��݈��Z��]|P;�kə�.@�I�:��WĀ8ڻ�/��37�N�2#�ڿ����b��$�nD.w,��6�J��;���#s������gf^����{a�
��G]�>�F��X��������}-G2�ʓ叛
~e�� ��#������e!ڴ��I�IL�QBOV뙘�|e/���	�/�jjX�;�qyV���ׯ��)���׼�~���wrh����B3��I�^BCG���19���LP�7'Bڎ��Z0T7W����>C�Z�쵢�N�L�7YG��:��\*9�^ZT�Owe_�4�3`�u������J�d2�Ex�J�T;dw��i.|`�@�����޿ln���d�.uW���t�?R�,,6Nݖ�!�$0��	��d��4f�
���{��-t�*P3V��>��/T��ۛ8�\�pe-��w�F]]�K��K�.9>|hz��u %#�U*���цz�K�
�z��c�ӄ������u,�N1�2����>H3�oG��8��e
MM0h�]�2��������(>�� CL���Ư9n�ŢS�UO��N^ɪ����^����s@��}H�ԗ��KE��{�B�Z詳bs�2���%ҋ�b��3�����\���}��B<��_׍��Ō�g~j��@���&w�hС���(�8�w��w��5L����6ȳtIj�� >>>�����P���paaa^z�v�'�� �)G[?��u"�<��T�H�e`��8�Pݮ?�H��6g��NǢ4c�����2�*Ȟ�۫o���"R�.J�~�%xwh�hHp=H�4N���ʳ����+��W�0v����{��*pL��ϗC�U�2=m�7�嬾��!�K<D�2�韮�
�{�x�H"P�ԥx����(����5�ӡ�ɀ(�@��XX���b��?#6/EC�'����L�&���E02m�����QZ��A&�s��Z�72Ҷ��2%�Kv�tt���SL{=�d%�o��Y��1�{�Ҕ�r�1W�b�k`Z��j� @%-}�H|�ߥx|�u ����������]����������L�A��W��RY�������/�G����,,�.�4�l�6��:��;�7�2���^�]
Hg�?`��m��I��z���bm!n[Ǉ6�"1v��_���#o_�Jn���/��I���՘)�BⰞ+ҩ�>y]���[�
��7>ߘ�n�e7�;b �ꔟ���a��h��I�I���F0ɳI�3�Tt��퟽ v�ֱ@�s����%�����>��v�j��N\�A�$�� G��](?e}��wg�%jcw�3�	'u{���N���@���+��6Y��^��X��ep/��X�Ԫ�E�x�O��V�M��SP14�50ԩ�<">����<{���dE]���}9����-�����`�8ϦDP�I7'���g�0��t#7~́�r��_���P�M	�V 	�ChRQ�7����?�*�I��S�d��쒰
o�U�oF� ջ<Q����uK��(�'�	��4��2Z�ڗV�)�v�Qԅ�������iC���[�f����e`e�-�c���;m�{�[���*	���������)U8DZʰ*�sH�D_9�g�跽~�k~�/�o{���4�/����y��-AYB;qnſ:!њ��q�&�]�c.�h�$�̼�rX�&#mCp�=x��?V5Gmz{/��}~~�Q��������8��X�� 5hc5�������
>7K"&y�6�����n�U��n����Rxe�1�����Ǒc��"���������|�q�x������b��(+ ͫ�a��566u�8���w%Y���7W���q��3�$��>��X{	pߕ����or���,��éd�.�����=0y���&���76�f��-&W'__#]ݨ���R=5TR��d�l���I�����jX1r~�(3%���b��9�,� ���"��Y����n�Z�_�}�N��f��tH��MOgꪶLʮ���*g�a�e�=���}�$P��B@	w�����#�� 	M���<+��/b��CջE�$%F@����CV|{p���ԭ?W� �kt��Z!�`��;x/˿&�R�x�k9������7<g~6:S�O�5h>�vFD�������y/cY�N��0γw[D���_q�:�kCZ���TwS�*�R�d��o[�ޱ(c�j=
��j�2�^<*�hJ�u����1��mm��5�p��H@��6�4[�����a����5���"��G!�Ɲ���6��2�*�
��?��*������o}���iM��%?�x��6�^�V����)�H+�{q�.�v�:�C�����~	�����^���x�UV5+���}:\�:T�9IF�����l�d��|~D��:4�r�ad;�腽`�q��~�(����P])��Ex�=�V��(v�5�~��	�,��f�*_�l�u�L�P�O��@O�� �D�E�t��	�$h?��x�Ω쾤QE�	�������R a\'S&)!g���R.ƒ��ln� b[��i��'��C.���i1�������&��k�W7NPF�
���z�
�TV�Ju9e�w�T��L�#g���ي� �Og��ȭ+�`�'ɏ̀����1�<S�|(~}C�d�~�~bN(��oM_?|�]h���dޱ����tV��x��(�=�_��0(���Ac�j�dJ�7d��]hi�!D��Oٝ'��u~����/g��ů0:�v�*�����"��
E6��;B���v���?*��QwX��)���b+^k����5�w�>�&ppk��_�J�d�*9W�%kP�w�9�?)�A�����b4r&�`�r�����h�!�t.�~[ZUQ
z�N9nv�g�����Y�$"��w�,S����s�$���@��w,��׫��)�2,I+~���(K�*��'���5%N�r	����AN,���.��_9#�j�;�v�bh�xJq�ᆠ����L �z =�c��E�T"H�k@(Xrl��}���O��Y��Ā�4{ '".
t.Mu�#�ʋnkk�1A�ÍJ�s���YC"Q(�ԝA�ӡ<���X���d2f���	Q9�#P�����D��qȳ%GM�����Kx�Q����7WO5�C���$J��mx8+�����w��!y�o�T�n0��6<-r�Z���~y7�� T8$+K�6�+����93�N��T��Z+�:b��F��mϛί�x��5����|����ו��?ip�wg?wx��c+y��ƽ�W��z�t�]��O���
3��Yf����_n��*�b[)�����"�E�U�;�"�D��5�������ɴ}3�0�7�s�����k��]�	�X��Ώq;��7(|J�6F�"��y��dd;��#k�'p�n��M��w��+Y���)ځ���;�4j����#�].���/݄�$U	U��3�,z�vic8�E��_��*��A��&e�Y7) C�x����}�z���sٞ�����bblj�~��"�[��g���o�-��YYY�R�(��`�	��/_�(݉���5
o�cƜ
�v1V{8e����3�y��������ó�����
��%����O��-/��-��$bN��t�� 
�t��s��D]B�Ѝs2h	����U�>yBN��� ��Bq��)�t����"��qBC�hu�iu�Nn�'|�S��F��=>������l���
Z��HJJ�(Q���~��+��[�q���3���V`8ۄY�\�S���&���A��}�h%Z��l���'�>}�7�$�2�n��1�h+2��%N�4*]=?�������:���w�(U#gy0����sH/Ѳ�omC����	�.m�3n�պ{*.(��n"���=��Z�~@�1�peQ㳍��F�U��t��9�,9��SA
t�8ŗ��##i�I���aFg�F��L{�������Uj1�"��ǳK�=4]fs~�֯!v��P�F��6��;W(���v�Ͻ�jЄ�0��s���,%p¨7���>ʱ<ϰȬwaA�O_:��|��F������5�vJ��5e����]5�Ϗ���5���J������v�����m�N	�0����G��GiiU��iߔ�?�/S���Z����ro{�r���me(:����;�Z9���Ռ����蝜��;;�pG�GF�$f�҂v��<h���!������E��[������(«a/ �CB%��f� ����ac���Τ@�C���(Ƨ����� M�W-���_��^P�L��X�����Ӯ4�حO��9BEo���d���������?�X����A�BCò�ڡ�Kk�����}��l0�QD;E������x�L����־}���3/3�i5����m������!�
��+��SN��5.�gy�y��q���X���-�(����G:M�[�h�/�3h�#[�:
t"��Z5?��x2�Y���ꤢ�{���Kp�yu,nWd�B�8-��C�٪x�;�M��#	�.b���5r�%z����;�lyiiԟ$`jyǷ!F�9i��&yr@�t��g�R�N���Omй�b/�Ϡ�R��"�.,z-N���U�O8	�V �a�©^�
�>�ڍ��>(�V��%;�75@5g������!0�U~�61���8��u?�lw��.ޔ��`��h��di�
�63��1X/.6��{�� u���w/}�7�<���k�����S����*iG#���A��T�=y��јV�ڍ�>b_$f�@ّ�����h����C}>��^Y"Yf�wx�B��t���\�<@NwS7<jW���S�7�J�	b�%�k��p�IpÉvНsR:��3M͎)�]J�M?�h��\k��e6G�?C����a]$�k�US����M��4�ڗ�l�M5�h���V��N�T�]kx]�Q���4��*c
�g��|<c �k�����W�J�/���/o�T�u�(��Ү,���kV�St����k��f���Z��R���#ʳ��(v�?5�\�c�X|F��z���������݇��>�on�*<�"�Ku�[����I��7t��=�[lfgf�p����p&�Z�mOƲ��T��6��1�h,8�^>��	�Ң0�i��}MG�I������̨z�$A�`�U�(P}���y�q� uH����  c�IA��M��7w�ړ�1/�v�C'g;���F�7H8 Τ�I��Ih�����VaC���-u�l_��ٝٗ�W����
�|�ƮP�j����1Lx�Һ(|Л;�I�%��k����;���}�k�j��T�ڍ8��br ��4r4}SVm����XY�3���9�P���u��^���c�tU�Ӈ�]��b9�}��V���6��ڰ��07Zҿ��T��_#�p�����>4^.n����u�w�A�"\Uov�.��h���0��>������6���@3���F��b>�(���9����-�k1�Ԫ�R�fT�eI~.�C{}����3�+5C{7g�����@����o5���0c���KM�[	ƨn�M��!�~��5Ԕ�Mh�:�<��{�M�ܐ]��k\�¯�t���ѪhoN�"z?�w�N�����T&�/^�#j�WK��j� �a��-��nf����;Q�g�9z
��n�Ãs�K݋����l2Ko.���A��z�U�)ܿ���f���*�s�Cae��L��q�^�O		���y����:��D�����|~��L+��f���@A�y�����hj�N1ڗ�X;OiX��1!g�؏T-,\�i�|�2x�S��i�6����]�:a������?5���כ�� ��!��Z~(��U���,�X�`�@�.;�w�PrR��8�k�u����o�}�
�d�P�N��X�-���f^��%�7�r���Z�¹�����C'�$C%�n��+T�Y�n� :� a3��WU�H�A4��K@Ԩ֜x�Xd�B�d��C�⟩�������m���ac,9�����m¸���-*h��^A&Ī-��fͣ����J
�,
�5��{�Q�cZ����Z�:�Oz��q����}�
�������|�WF��;TGք��m�q���FI�KS�!G[l�R����ׅ,�tn�s�ʊ�Ļ��6���)mMM���ߍ��K�ؙ�4��眓=��V��md$�ǩt�QK��?�E��2]|)�������5)��q�t�p�C­��ԡ�
��s7Z�+lH.}۩�m䏿������30(4���r���:�. %G�ם��%]�{d ���h��^�`R�TKS�5�#�9p�7�T�ϸ�IJ��!�������?'aD�h^���}*���Q(��N�*W�O�Ҷў፻�Ka�����+4��
 �ne�CG��#����� C<\5�ۏY}D
$�Xsϰ���;���T'ϑ`9,�O�TܕP��8լ:���%�E��eg��}�ϪR��Se�7�;��UIb�kk7��&��ԉ�<��U�b��z;x���N�R�3���=���L4<��K�8ǟ� MA����c��|į���ҋ3%�@ �C"��(�
F��?��6_^Y��b]i�����ƫz���^���
��>�Ԋ#TT���W���\=բD�k1�����o���g'����s�H���N)F�Ȓ���:F
(�Ui�\��]%V59���
 
I��k�+hgG,�h��M���-j�Ū^�ؠ]$|�4��{�C�tzow7H��-������	`R�:Hױ�5Uy�	��	?���B�Z�o�5��K$�_oȱ12���eQ*F���L��`�~n������й��m%c��2�nC�1s9����:@T�����s?o�bB�������{�Z��=D��@�-sFÆ���J�Hm����]�Y>D7��Q�t��d�#]��My�E)��m{�݃���s��I�V�/��Z�0�E۪l�4��?�"zv�4Ԯ�L�ܺ)�a�p �<���F�w�Sn�n����e l�wN�vPP���J��źK���&T�8�gh��C��iW�NL=���h^On��O���-��~�Q���o���j#�DX.+g���o��ɗ0���2|i{���N �!����|h:/~=�C'�`U/�U�]7�7.d��Q_`�Vگ��E��/��|�n|m�9�	�n5�FR�Q���Jm ������-+�q�Xk�J�m�#� ~j����HdHش��b"@�
'��YT=9p�\2U������yhv
��і�YXԕ��_ �z�]}ȧ�W�f8B��f�?�� ��� Mjkk������Y��}y���7�î`* bX�h�Q�$u�n���Cu�!���V�!I|(���V���{����J�$�s�x���8z@|m]]�ΰ(�fC�%t�z��z��/�޼�]�� �\�\�,]�6\��Qw�gp�?j�d��9Eg�>��YMؗ7�.��%ݱX�\��XT�%��(�/`��(wfkk�40G�9B��?�C��2�X~�\���*Ԓ/��}�]��v�a��U.�mmvG�0c�ڙ�Â-��V�<H���6aw��G�ڝǗ��.�w*�%6[{�m��"?��Gfe)��.�R8�$gx?G���|;?%e8��PT�Y[/f$%��8��޿G��Kw�F3��|������E�����PM���O�t�2H�˯]s��#1���J��P}/`PWk$(�v�G浵������j�Hf�# <�fgmo� #=���M�����\u�查���3,TF������zJ'�fV�4	d��Ɔ��?G(t*�7�n�vt*��	D��/��+<�_�{qNyr����b�1��*�Q_�[�@ɝb�c�������P#D�^�d�404O� ĴI��*~�r,��t�*v��#!G'����
�=L��mI+��g-��K�c�� ��H8Vh������Pҕ�RC�LP��fP1�%?Z�kn�~���ՅS͊� #�X�ud�(k�����[�98�,ȅ]�% u¾���� e����v��: �&��JpK$����|W<3�h%ῒ�Lp��48X`�;����	�(���a��Ԥ���hլSmN����.�h�j�Tr!06F u���<��<	͋R�_��LL�:�g@Ӣ.�Hzx�^�v)7fأc����� 7�<����|�`|i� ��̴�Ք�@��������&���;����x\�i-T,��yؙd��=p�(�^2Y��u�U7___��U^��Uk�)pZ�#�fY�ޝ|����NF}tK�a�ן�i���-���d�P U���q��������kE��

��N�pg��o�7|��N��ƕ�L�bE����D"�ɓ=w����𹅅�x��e�6F��-�>\)b|�#�#k�Q�<GhT����t�Fj�b�'�-����w��Z�?P��Bh������;��&z���+�w�Z观**^��#;��/�ɱsm�7ط�hyi�ʛ����18����
d��1�Ċ]�����)�ij�AG�>n�h��!^����s!�i�U��������M&���G6 t����g+޲q�e �R��3�kg*N3�-����9�k��������_CB7 '&^ �6����@-��T9Bٔ�lV�{<��\*����HW�]����`�t���l_��iP�ڰ=��"%U`ꢌCV,o
��՚\/u�} ���I�`"*�$T�vl�B�D����Y��#�k�}���~2����6��1��w��֏�uww������#}��q�=�ov�����m�-Kcg}����J+9e�����r�L�bT���L�����;{��uw�����n����UV~�z�Ư�=�[l��8���X�x��M�M��=��mq���ӿjg� ��@L{�/(��#B����ʽ:E�z܅hc�ĝ>@e&&���~4ٵ��	�lw��F�־B�	���tgE:����p�h۬޵e�rc3e���v�`�j�����2�<:���>���9��d���#!��Jl��&�����t�������`�3������o9��iQ�	j9��1�'�1�����"z�y�4���_Q�����{ĳ�~#�jo}Kh:�3���2677�l�� P�֐H�����qS���?���ݟ�����&��QW�~B�;�{��P7-�mycr!��71OJ�0[�u��N+����֤����`}>��O�V+K ��ȱ:>^I	�jR��t�n��r�s>�ʍoL�e�zI�^�#�䤧���3�_Ct�?}d?�@�,~N��Yh.5�1�����o�� ��wyܻ[tyI���v�0�!��-*��e�(�}���|��б��k(6�B��p�!�5���s\�gz<��h\�lܰ�j}ܗ�t<��5�#?��XcSA�a.v�:ᐲ�������:�&�ݝ+܆���������כ'h�r�B��1����hAD�	�͢��)g"¾�@:;�{x�w�̚��4o������`o���lj�[����8���Y�]y���%)h6�m6�a&��z�f7n����Y��ڞ#�%^3F�5�.��뚘�M�VJ��|�N����x�<'g�e�
�ڸ0������heuϒ�z��3c@+A����lB1��b�e�Z]s�rNs�c�������:m1cI���+��;!I}񥓢�oc�?އV_�g���1�sQfg{�����k��J1��x�X�����cSZ|�İϕ�[ǭ
��́��c��+� �[��Eu�,~������T�<��C�H��@��I�vk%���G聃���'+&�f���oj
���]�4@a����i��Ax���˖j�j������LLLjV�A�����S<���|Vw��l�b�luzp���ѣ��g)�;��K&��S�n;f�)����Ɣ��WIM�2��c�N�K!eP'$@�6v��`獵���P������#t��C��n9��>8%/�Đ��P��e}(��y��cX��뾱��}�,��Mw�ւ�U�jkE������C5��V��ho@? ��ɩfc{r�bF�c������?�RA%zhӔw��Z�M2Pu�p\`)ewWd����S�X���P-��]w g� �zM��ɃL��UT��ͤ�ٚxchtP~�66F��&3ǘ�Vm'��X��la >���8s_���q��ͅ�����Z@.Z�(ѱ�����o��ola�[k��|JLT4�~h��-�ҫ�=T�B,�9�g"ى�e�&��2f;�L`Mdl�����L+�����ݟ��+*�RN�^ˀ��d�������ag���@��@ޑ���P�
�v������$�#��tFWo�wWP�@gy��*�vTy�C��.�c4<3���ʹ�vsҁ�^�xʉT1Ћ|�ľ�؟��#"�����[D�i������=�z�����g;���H�ӷ�|�b�����+��h���1�X�ʼ�Dq�]���Ȥ?μߧ��k�	�C��&����o�Vy󹊖���!%v�����[*�U�*�P;�a S��h�Ym���w2#�����<>����w�	����$m��?�i{���E�����t$8��%y��Ob��\ll�O	N�j�.[�ݲU1%���/h�s��'r�T'�����D�]��<�>k�'?�~���꺕���Onu�&*f��$���a�?�ح[ �%�� )/))X^����Y%J}�mT���:����g��/�`p�1����)�W!*���u��CY*�c��rZ??&���8B#GLj����83t�TKKIؗ�ݫ Y-l�PIJ���!�n�UYD��8������Ą����i�}��y���0�諮�v-�Y�c����{Z�Z� T�DG1�6��O��?$�^Ze�O��k�[
�$�+$1M!v
� .A���DW�C%P 	�pHV6hqߴҴ�B�u��Y��l�8zG'73&Ʀ���ZF?E�¨UlD�rMX�r��I>��n���.��㛾c_8��=幒��fy#���])�I���T�0$������5˞�ȍ.���Š:��>p�b	D@O���H7�>�t�N0��L߳����^���u�� �cwT��G�����e��m��e}%�ɲA����09�,��o(�di��C<�ַ�s�v��=�?=\n�~�z+�~����0�G������\��\" �'m��r��@l��^
z�7�3�}�< �=d���`�,&�Ͽ�ȁ�A�qB�g>i��?�9X�{����sGGO@�k�]:։����C���CK���c&b:^7��x��B�҃�>��*�j>�%��,��ω�zh=|��`|�CB�?ڢ��w[K<W}���+.�����͌3��������ҟ�7�-�'�I��>"�=Բ{<���Pg+�1�ogGDh�S\�)9,ջ�ig{�F�
�H�h�]v�U�FA���^�<�Ψ��A�wY�����Do�@�Q������=eD����T���\�n�bB�8�����3����#q_�"@VfeA7O�}�TW���5�_l7�aqj������錇���Bem���jKLk�{6&%-`�xxx�-)Ȟ5�Af��_տ�=Z�&�{t�k|�g�=�����R�^��MF�bu��vЀ�1���ɴ�D��q���Q��Ҏ��=K����67=�Zhs �.���s'}���KG�![u�>Q��]��-���G���$H�+)x�(���f�(��)���Rn�w�)�1$���k�I�մ+\��:�>}J=�u���;n����f�� �k ��x�e� }��h�N��A"�y � ���1lw��Yj��u8���hC ��O	�i�ӵQ��&'��o7��nL�% ��rs����n#ɪYPPD��A}��� �N�:�b헀s�4���3Jw(!A�սE�\��?`��x������nx��72};���w�I���c������x5�S��޾�F���E����t���
3`zQ�����o-I(��8`lf���P�2���	��q������i����C�Y8.���Wo����s��_�2�Z���3`�<��������n�ޅz-���}]]��� �{�i���F[�@?�R��7'4Z�)���?G���g��=�ˁ'v� IA'�?a�JV"�.��c��p;������H���L�c�ss���x�Ԉ�x(������!9Lp�;�ZRR���Ϝ����s�I��f�5���{���ai�xp�i�����WJ1!��������������%�<#���AA�v�m��"�.{ػ�j�=��BE�:F�]H�����?���0�P���[d���N~���M�[������U���A?�1�$?���^�X�&A:��(Vk��0E74��'ï��.*#�����;�U�n� �j��"I��9ձ����k0ļ�&�И������)�˿tsl8�����TyR2��q1��S��y3��9�������dp��=x�\������}���#07	xE�6#����$�r�S:{��j�����;�K���P�9�1c��Ǚw.a��ۿ%u�t�(U�>���Aii���+� �UBJJ�����߱Q4:H���?��@�����IHJ�����3}���&Tp����Pu�9���7-e��h��1�}Dp/��N��"%&Vh�*y�[����ڻמcM^bLi�,��_���α��{Ȱ�#��$ov��IIe���d{;fbr�������'ؒ�xQ7�;�
{m�#���4�՛�����6���Bܵ�H�r0��/���!��vIW^�v�� g@d���e�P���" �A�r����\a�f݁2��3�	�I_@�/�߽���(��wm�����F�	@�D�:B,׀�=x���s%�у��Y��탶�l-��mHf|������j�d/x}fH��:���4�������~^��&˽BB..�~���aB\di<�L
lZݢ�-g�lы�7z��I~�g[��o�y������-�
��@��w�X0��V�^5�%�	��j0�� ��2��{���������������HD�t�޸�,��������ő��ِ��f�9fL"s&��Z[������/C��<���~l�Q�-��,�=(r�_ �媭oI��_w�t��)\D�#''g򂤤d�nw�K�1QI	��!=ՠ��{{>��c�x<�[��[�
�KU�C����/��)�;K�1�
���A\��3�+��� 6+ PMW�{zvVz)��Q���E�:�!�O�� Yq��Q7Ru�	O�&%�h6'I�[^��bKٹjSzpe����IJ�٠��鐤�r���hxxc-�/(�y�lw��B�ԩ|8�A��4�����9{DD���x
ԟ��Q_C�1C���f��15��<���ql�Qٵ'��������������0?>:��۷�P�����[����#� _�:=K'����+��6F}�+a� ��ˍ�: 髞#I4�����]!l(�:p����-�ye;L�_�¦$��f*H9��|���Sa'���δZ�_�)���de�����2eM7��x�U����5�۞��?Ѡ�.V��RKl[�ْVv���,kf��8$����y��_Y��Qʱ"�7�/N�P	�����.��1x�g���i�F=�Z�� mѯ�nzZ�fym���=z8�|&���q9"�k@q��}2����e'����=k�1��ץ͔�o]j��M4燹�1q���������:F���,Zl�wh�����R-�n���F����~v�ш	�X,X���5�z�/B{�Ą��ޣ"����\��K���� �Ꚛ��$�`�([9�]C����RGd� `�}���A�}������a�`D��F��TG�V��4�~�����Q�d	/U4z�� ����vq�u�n_�O�X�a��0&�fA����
`%�
� �A��[;Q.AC*�Kr�ah�q7�"E��=�[K"�����o��ꈲ��z�9�f�O���Z�h�"���'��;xmct�������Fi��޼��T�\22��\�k���n�����D�2Xē��e���i���:�[��-����H��"�چ�Ln�bm>���Q��y>��@�10ЀJݯ����#p��GD�P�L��O_��u�Ի�p�v��F�T
�Yx�M.�/f%k��|����\?�/���pK	�p �-�V&��j7nY\=���\"�Zs
���٪���
����B�eJC�;��0�=:�L20(;�|T���u��l�\W������a�<t�.axd.Ĵӥ�^6�������Y����ڸM�3"� �P��f�Bp�*���\����S���:���	ך�{tp=qp0	�(tƫ�Z�ʼ2<ʺ>��d l� ���%�_QQ�U9/&��vy�Ѭĸ7��{<�T)_��ۗ��S�5e��t\��s�ӌ���oY��d�����?x�Ů�y��S���%�r�Ue��>��p��`�0%O�ɍN	ڎ}ӆ�|ߤč~k�)q���?�R�9C�]�z1����'�׫z�q�l!4������l_"=��3Ր]A]��d1�n|�YVkMsn����I`��:%�mX<��$�J�t�]W��4�U�EwllL�k:�T܋H�6��9V�&۝���)����R���Fkzxx��a ����$�#q��9���@N�1c;�Ph�	�b'�Z�m�w��j�|����d)_�ܞї������pO��8� EM�$��j֚w�4���T
{����W]���~ඪ�o��\�鮚�7�:|��P|i۟v"�KP����mn�WV�7�5䏋�=='�ڵ��L#	�O����f��'��I`�t�*z�N���xn`D��P�7Ѕ#�4����H W�����K�ʪ� {"�{��
�v6}��#�|�e���ۧ㳯v��M[݋�if�ǵ6���p�����8Wk3��<D�#�޶N�k����ШZ�Y�|��3
ڙ�#�,K_m�C�����j�ҁ��̼t���{8�lvV��6�E�K��N������o/��'|��*n�\���>JY兕���dV�H�ka�;R�Ŵr�Zzc;J�J�pb��k5����`�����0��`��)�@_^����EHp"�$�x�Ʀ��v��msɌPL��/���S�8�`-���:���=d��gR
"�;��9�w�������wqP��C L�6���]<���v��I�h<m�JXƾ:?wwU���(�yOqq����2��(L�š@OV��R����n\⻎�]~��OT�q�!U�{�bT�V�(�۩\��;�Ǚ�Ha�l+��)��պ�I9<��2��O�ƞ����UJE�#$e����\���cz��m���,6���~���]t�/Pbh�[���g_ZG̙���uȌϯVYme���*��������g���^��"�B�Ԗ�x\z)�o������c�w�9{۹����ʅ.%Ͷ���ZK�*�o�W5�����M�ޛ���i��Kwy�څ���7�MB���P�%�������6Ck�����a>P¼���_���s
�]hPk�#�=�I�a�d�}�`{I��;�?����o�����h�_���Cx��<Sh��{��<�|����ⳳ���
���t
[ZW���4_��Rv��mv�)�O�e60�2%4:3AUk-�E��e���:��@��كG��[K�	��.^,L��f�n��H>?�L�Uou���O+ZJJIH���R�]��l�g�[�D!�}�"KCI�ck01J�%�c	��6���}�.W\%s��>�����rP��\�]�F1�f1��1���{�*��Q�ϛ���o6@pfB��n��:֬t���9�NGEG�WkYL���kk뤥�
��
�)?�$]���9r�Jd>��FR��-=P\3���e�~zSh�+�h��d��).!Q�������:�yI�{Y�7��`�� ��,�� +|�����u&�!"\�����5�-���_{����q�:����b8�Q[���hx���;�(���F�H�1Xz��9��s�"�����Һ�.�
Hv�������y�����`��#�D�V0h�Z ,�>��5��(K����76A��@���i���b�X�aVȢ%�N����Iw1���t�`��ݫ�,;��̻�[e�IT�� d�F����b��qɍ�K�"���]ŕUU��-KMK<���1Yw�y��y���7+���^�!�t�u�
[#7+�����G[�Ui<�6G������^�5jVἡ� K�T����1-�Õy��0$���/�l�毰C���� �b��������V��W1|mg��^���L��:^��h�/�w���,�|ͯh�N'�Q�ւN�P���=:���q��Z:Y��o���x�g�,|9���]`�������-��
y�=��ME�u�H�m��|mb��������B�K~b+26I<K��4{�ۻO1�uX�J��Ǎz�+y ���$������А@�

�u�v�. ����Vy���.�Vw�?�:+v�������ՒS��8à�\48XW�u��ߟ��$t�z�}�~ e�߿��`�𻤜xc���^��V�k�_��?ج]:ӎ1_��w/��ݲ�^��w��
>?쫝��m�c����/������=d dT2�pG�C2��s7���˗/�I�G"|b�&��G
tX��v����3Ul=�����뽏��Y���G��**��hu˭v�����|�M=R�+ ����g���/ķ�³��HW	@��E����S=�<W=9h�������p����������I�h��1�e�m���F�U*���~:�� |N��^k��0��g���]�
�w��Ƙ��=��r��Aj+s���$�	�_���y?4��6�(��%��C���4��ۚ#�ൔ�7gR�s�V����c�/�2m���󹕿o�����%�����0��36�hE�-�[��`-2,.�oWc��x#�=?r�w�Yk���΍���q��9�.7{�5����h��B��]k�Aa�����*�ߚ�u���*��|�����R6���xB��$��g�B:l�[���%���B	�S	F�z�^6��b_�G6�ȯO[���)�3R�<�����2g �hDF��?T�=v��۹x����ju�T2x4���We�{狅N�Y���q�ji!vb5+N�%�Ea	�X���ג��
;���jp������.��CϢw����^h�k�)0(�	�����x��%K���>T�s<X{��&�sސI'�d��8�/��K�z��Y=��w�}r �$zJcg�I����i��q�y!���:����5��p&��~U�ǫ�˼PMk,��x� @8�z��iJ:�J�w^9z
���Y#�����"�\��y�����h3��Μ�R����|������ʷn�je��
 ���Z�L�d6��Ae�AL4�]rnkٵ@8��`@4ud;�%pU<��Z�p�X8s���Qd�!d>�]���T�P��
r�䨟[z+����~�7k���'ૼi!1��>ۯW7��.e��d���g���y
	���Y;x;��%\Y��&� ghx���v��X��Ǫ���qY��dt!���_�<�,p!W�)  �7v~o�z����c�*��b��= Y��4�ހ*�V�A�tP��3����T/$���(꛴�膺{)a̍���[��F|SC?�'@1<��ϱp-���J�a�'V�\��Yo���y|�Y�����J���i���'�̑� �rtu���I���2���o;Mn�eGG���X�{q��牕=��J-9�e����՟������b/�L�+M���Y 0�����v��7�h��?1�W�B� �ƒ94�}|���ﰘ�!s�3Fv�#�p�E��p�� Iv巏�=\W��3K!$�p
��+{�ĉ����9+��1#2��$[)~��W�졮�Wl�E1��37S�{��l|ۖn!Z���7k�s�S�A���>��{n���ɦ�����f���L��W�ڤ�\\\&��Ft������WQ��J�fZ�9�V0V��)�]��Z3��;}?�tZ~f=jr��f:�-�+�YT\����/�g�U+YWhVS������`;����|�s�}��lVx821�f�#�",��.�/�0^,��ƣ^����;1thb'�%Z+���z�0�;��\U�p�Ω�1�F�?K�{fsss,z*"��W�y���1X��l���g\--���F��xUF�F�cU�����!�?�hQ��R��|�t�!o��諀?�ƾ��bbb�l�0�� �2��ʗ����Ɵ��������(�fWś�#�ֳ�g�;5<%�}��P׈��I�d9����7��=�bo�>Q>�����V��ipAn0�IB���+�K�-�s�vv�]m(Y$�sK�����ҹ��/�S6�ee!�:�������7N�9N��R�����NRk'��S��Y���s>�~��N�WWRr���4nsjȊ� XՏL�țl�B�s�{j�o윥����d`}����G%�x�I��Dֶ�||�����u{"ӿ���,v3ڰ���}��5$��i���������)0�C1��h�^W=�S��s�O�c��>�H���gKi�?���4Zo��kk���e�j���1���lp.�����<�)��6�o��9L�+�B�	^�S���b{�e&����Q8��Y�ɩ��]���|�1^^r����ĉIj,[n������tڜ	��<8i��-&�m���YWW#�:�ܣ��*ccc'O�Y�m�`�I��&���Q�.Kos*�jG �D�Uz�z�����!�{d}v���Xl�7n[n�b��yT��Bl��j�͢򒷗�������]�3hZ�$��o��&�C��R>�=��FaBI���H����J�)�ɘ��>�1���APr�V2���?�k{!d�{��U�ܩ %�C�÷��0��QM'B����uM��1�Y�c㤵*@��ݕN���龆�r� 0^W�?�
[ܤ[��n��RFx�c9�>��r[�
�΋6tQq���9����߾��r�ȗy���	���o���UT�N�����'t+��!�@��f�n��j�2���iii���[0e��d�|�,G� �d�8$2rǛ��~�xc;B�y�!.+�]0N�D�_Ѵ�wRCN�v;aXPW�j�4�]�u�^�}M�/?�Y��<},� �������	�X������|xP|W*炏�:��]ڰ^!ZmX����q�b���Ą�F7ʌ%������
纉�t�C�V:mSĞc�Q��Dے�ox
r����~��/{�Y
`7_�|FBJ�w��=r�]ss��A3�����n��浢�h���wJ%ee��G�N7� ��t�����Ip���wt�]���C�b�r�0h����Β�� D"q�D��Q�t@*:��ܝ��)�~����"�`Y�|΄
��֚Nn�F\޿����T�R�a3R%*�u�oy���->��1~�\���!�P�L�V��k6�'oʰA�OO����N��t
��:�nIR�<0X����kǞ$���dوf�O+�Q���(����Q�\]��DS@m�\]���K�^���%�1ƈ��jv.]	$��D��ՄL�a�R]��ع9�T[��ϒ�)�d'2�{R\q���}Лڒ�f�B�X�����_�=����&:���6iE��@�K �[!`���0J�̱��is���u�q��N�V�$u�uvuu��W���}r:��۹2	�F���.1,F���M���B��@�2� �w&�Z��8�i��������?b�Ɉ�rD�� ��ԝ�v��2�2T��������U��z�L^Ǖ��޸$��舶�>YAV=ooC�����8[c�Z��C#�������+eD�=�5����!5@�N�[�5��V����qa����e��OG'�8{�$ H80`nʞ�YdwGn�w��XB��%)ʼ��%��z�-��Fn,��Lw����"�	[A�~�h�`���O�숱�*.���ؠ���=]
����sso�u�T��!�JK������F��z�P`P�W� ��)�/r�Gi��##C�R�.aH�0�����Z���%�C�
 O�F��@���3��c�>ux��� ��p����³��p]�g���Gk3B?ѵ!�I�^ �x����3T����f%R�L	�D�Ϸ�K_�>x���� �¥$5��աX��F�j�!װ�&u]]B���<3��ܜ���)|,m���$\4ʃsJ7-1���_�82�BE�DP6���"�(�47��B]0U�q�O\��B��n.P��7�.΁�4�n��͝��K&�X��r�.�b;��&5:�FB;���94��V���eP���4?Aۊ� pI֝���pq�����������2
�����ա��dj�ND��']ܶh��y�$�ͩ#Ҏf�܄N.�G,��y�ݛ�t#��E$��Wy��嗣�=�"�(�#}����7��&%����m���b���#W9��ss�E[�{C��8��:�	=a�w�a���,���x�ދC�G"[�k��a�Ļ];t��L՞��,��tG�Q�QMw���4Ҕ:�P�fgV�5`������ǆ�ZhW�R����B����9_������vuyA��ó@>�VihT���! �u򤽝�)`�?c7*��^���#��������Y�=�,�:<��Q���r�;�����#0��	br�*�fo��˲Ȱx�5-�A��3C�}���Xc��4��j$&!?����wᠭ+�Z�:$v�ā_��220�J��F��~ȓ�V�����k ,ȗ���,B�~;4<[������ �2:��bзA��9P5�ݘb���@"��{�QTC/'ǚ�ĉ�\�M`�pE�����;���T����GNO��ӂ�WMɫ=�Wq��!�U6���}��˔�m5�V�Vx�����?�
W�ʕ���f�1%�b��sôw���j~�����;�N-��Z�ۻ�F�_�^���|U]]>�� �7�'+�1����غ���D~qII'�bT�^���{ܧ0d3C�	Z�%V���{/�o�ٳ>D�H�r�T���,elV"��>��$a����Z(\OOOKK' ��~�r)��Β�fBN��*��R��XQ��h��Ro��+�+��\:tamm!`���i�^�w�} Q�\�և�}΀��A�^��i�.��g���b�v�R�by��Y4�%�lE0�X����G�d�;����m��%?����W̑R�)�*��"�oox�������䪪���Y�U1�=�T3�X��ý��o;�A�s 갇2�2��I̍��A�
De�>,�"f��U�B�f��S���j��0�6��B�R[�1�-.t,|�?eDW:�b����U��έ�Z�z��N2��^�����{@)��}D�e͚%��W�%x� ���Xu��U)���GJ�` t�h+�K�"�zNa�W�y�@�����7Q�̯F/ '�h�,K�w�6��ro�֚m��j9�eŭW�9ݽ�ָ��Z�����T)�f�b:Pd��;���� ��P��ңV�:�'��>�y_
��H;������y���AC"��9�K��b�s}w�$�E�v���� �@�&&%�n�Ei��Z�vގ��*8�����M�������U�[��r=��<]�U��̥�얒���W�6�:���_��텂h3+���k`���rt�QLZ	�<֢�
�[{1'=��֘��?��R'&B%$�ɜ���n�O!��f���`;!�%׳zBlP!^� .�?���O���bh�s0��l�Qa<ɓ�)X{�ռ6�B�97��}�h�伛*�b���f��=j߼z%��-�Y���r}}]LD�[�=�����5gMYv����,} Q<<,o+���)�D5�MTcIi)2e8*89�����k�&�׊���Agi�ʲW���] f��W���u�-����|�;i�?�ȵ����O���%G|�76�){�VlEӒ��Eʼ:c�j'�5\�r�1�G.�&���V'7k#>�������x��[|E�d(P�o|�����A_�B�����+T����)�	Wˍ�˧��������!<� �R�i%Q���#׽!��f�w�T5O����8��l�H���}����K��:8��|]�������*y�DG��CS0arrr�ﺌ��)N��J�,U{PB|H�mf�����&E��Ez���rF�ѥ�oĵو�cf�Sb��1a:��`N���u�;��;������P�:����fBۧ���O�f%Yn�{�޿��xd�������*$�Ψ�BO�����=���T."��
�׸���LG�{�t���*3P���$�`pV]��s�]���0�˗u�B;��d�]�\(�{�6K�6s���-���5�f���kY�b�,� �ey�l��uvVK�G��:� �¿|y긹j6I�{nr��nטo�\^^^v�{W{����X��W�X�K^ޅ�
��- -�u�~N��|1�BBB����-ԧ.?��v.�+/:::�\ZZj�"D��俗|�4�#��t��X�N��)>钘��V�&�=p��:,���1E�A��7��ʉ�$4���ri	ٮ�ЮJ'�N��PHZz��NMc���P�q�v�)^9G�������R��F^B��OL�߇�"3������Q!X��j��v�눡|#!����g����4�����?C����5���/-jX��0N$=��M�{�PǀZ5�spa��|F�ِ�Ƿ���?*<�m���Y[[���~3v����*םP|�W�2נ�?c�{9=����n�X괧�)0I��������}�=ϑX;���������`Z�'�e����"�Jl�!�����<�K�X�=R�_�����Õ��|�:]\��/2��Kt&N���GG��bp��zTĸjn3l�5�����b&�¢=||
h��1$�W15W׌R�WqcR�Y#���3�>�v�L�0��`�闒�1�Mg்	��C��T�{�W*��ߟ|�d�`�Dr��Y�̸��>0�$���Ao���4M�<m �<�F�Yx`��'� %D,�R�������1�#����I�j�ֲ�+#s��f�K <�~͞#�勼N�A��04���~���j���D	ZvcZ��w�eo~>��C�K�bV&�r;Z Y�@5�ֽ ��P�盠z���z��is�Z��(ă��p�f��� g{;;5�=����&�e^ai�˸�UDH���-1H�No����*^�Q�Xx�X���ɮ�}AV�(�ޗy�\{?d�v���/�$8���z��'�ڒ�9**j&W88�Dl&��#>�2�{���VfO|̀�jhiu,ME/}�62ʇa���M�n���;ς�	@_+��@pq炓�� [Q��]R�1�U�^�NNzV��Ι��O�	3(]�N��X
h܃�n�����S�vf'���ho(����\�S}Œ����Χ�+���W\����2o���B�\�C�����܎F>�g�"G�յ��=7s0�5fB ��P�u�l(��M�XmKK�Z�F���} ��b���`�Zѳ���5�� ��_��z�%w�oq��qٕF�&;�!lQ7���ַC�V������	���K�����[�����~�ˇ����x���0R�W�3_���,����Ӆ��\�+1�#�"D�����`>���LjC$�YZ�	˧l7����$&�F{~p�MNN���r�Xzt���j6R�m��9�����T��ٓ%d��' s�n!Z���b\иw�֙39ӂ
�&�� ������e0��iii�K�Z�Kssm�Ly�]H��R��xH��y{�'��b`���na๠:����7�� �#Wc���K��B=��G!�8g�@�\F���T'=j^?�!��)��Jm�qG���5^�Qb���֣8��ք���ۜ޴�n>�`�+4"�L	+�K4�F�i<m��??��8@x�'�j���U	ߑ-�HF]���4�9x�_7I<p��Zi��\=�&==��N���};J�	��ydE��G[��i/{=`�,�o�\�{`m�E�Z�(�W����a�z����3	30�6yb�?h����]\L̬5�8�˛J� �}���� P|y`:���k�u��!>�Q�uϞ�X��G'g���$��0�C(��/��m��zw0�^���j�|L*�8�d'���2�p���?���0�U��.s\Z�=;�;�<1;77ݕF,�o6HMS�)���t˽r��C��4!�xBG.�����bE`u�(2E`)������~�G��hL��q"*�%a6VT��T��o��ך�le�$�D6±���9� 5�.���ևz;.q�Ĕ�M^��9�V ?������&/: �+��^�cvj�iMM� M��|��և�ӡ'_D����A�03�ܡ��@��H$i���3|�����@����C���~�Y:Mc�ޱ߳-����s���?�N���߷q�!QL�`��ʌB��1H	�G����!`[� �}]"���:	Eɹ���c����J`���逬Yߠ��������������q�+�G��ب�Hp��-��.W7�Be�7H�l(Ž����3��ʣ��Y�w���D�p����=#��SW{��~Te9X+�R��>+�X鬚Z$�[�++b42=+&����NWV��&�C��@�>~��~�fj�J�����7�(쟦)�?~ �F��qq ���u�=xp>g��ۯȾ���p��F��Fv���$����ɞΔ��Y)��x����щ��ݺ�R�l��g��_=+�X�:5��tV��^��а��m��(�Y- D*֚�*]�
�dW��*�*��Y=��������C�?&�D��*���-�
2
|�~��F� ]gZݷ���W��pU������;{V�6���:]/�z{��;ϲ)l���^K�fG髨��Z6f����#�����2��$i�#���1�f�܇0'�}�&�r	i�r�Ç�`���Z��D�_,�h��̙3E��Z��Yb�p�lL(�R�Уߪ7�`)��r_E
[%O��;�

[\^������ʜ��/~
؁	�P�p������[�I����]�é�1�DE���yN�� �O�
��<��H��?^v�M��uŎ(�;F졘[��fFF5��u�P?��������� ���N������?��S�G�Bq4����h�����ު�����1��JWQl�-�SQɑ�j���LKg$Οp��#$!�TH(��w�<��IX���#hi�Hr���藯ױ��cRѥ��M�������g �ݚ�_�ܽT�D����!Ӧ}���[� j�9����e8����>Xɼa��K��)d���jg�#{i�Ct���҂R��z��uz��sz���9WR�!���لh��Л�B�[�8
r;2��p���ل,qfxr,(���M ������!uZ`��h�;�i��KuEB_�D^��{�0KT���@��؞㙚����ю
qq�\�I�%&&�?�*<�W]�W?�?'"Է�*`?=]0` лp<�ւ�u%%�i
%ɖ+xl�|��''����v��7z�3%�lT	e#��*�N��l ��ӎ8~����*�;{�ZX$5<�����L��~��tu�QfJ$-	++^ ���@�J������\���`��T||���oN��8�PPKM�)� �2��	�l�WV��P���,�B8͉ͥC6����e��Vqj(�!l�/>ڂ��Zrm�+�r��ґ�����ʎ�
뽇+ݶ���!H����<G���S���0%Ƿ��ب>X�sB��t`6�e�B&tx���XOONJ-;�X��)IdJ��z�b�����*f�y��}m�O���7��ACV\��d�	�:߱5b��8 [�?_�,�ޒ�{�����2W�R�ck��V�l �D9y���I���\���L�d?M�&`Ĺ��4���JA9z��F��%�`i1�rtv6����TW��)c�ӽ����}$�%�@�k��y ș�U��� ˻���-c� 7*j�\�;V���Ԫ�
�Ð�����_6H���R��8#�"&h���9w,���>�yP`g��7��X[[��k���w;���[Y)���H�C�He�\@Nb�i�43��:��?�s�AC$����e��f�e8��È��`�Eμu����iG�і(�T��u.�����i�fck�&��fi�5��	�
�#�D�dڰ�����Z�	�����y;y�!���D�ʤP!���'����}|�������q�ҥK̓n��6]Z�I�����������=:�_H۽*%�#�����?}�]���^�5f
����uj��&F_(	�i�]r��e�צ�kK��h����#�6M��ț B��iժ2,��������-h�G��/��Z��:�A^�piX'��v��������>��Uy
kN��� Zpt�Se�F���	��u��%mٿ���m.S�2\A��������;@Ę�p��^^՜/|�*�����K�	ي��D�q}/�+{N(>��1E��-�_4(6�l:���v]�(��72*� ښ���iZ#�]��xW�dM�l��D<�fX�9ڳ�=U�/��N��3��\�ٮ���h�?�*�^�.��>rH(i��pQ�Bp���'�PS���2v|�	cK�*@V�>~DP�$�?"�&'_V�때��"ǆ�땳d8�8��>G���������8��WKHHp��= z@*z�	�b���ǎ"Lu��5��Q����,��Aw~�Zy��x]`�}�����};�㡊��$nlЉIK{�G�fU�x����|�E:��?���͛7�	I2���3H###ˢ<Ժ ���q�DɎ��˧���Q`@�~�x�1B�8������FO�s�p�^���w"�NFZ��e>VU��l4S@6�����1?�J��?��L���?�Tw�A�ς'C��
�|������{`�Y:k$R�Ģ���GV�!VwwD�������C/Oc�_���C�T	���:���{i�mN�fG�H�l]�1'ln�j��N0rM��u6�����f��1�{G^M�xIG���>!�BK(��w��o��g�N�<�����	$xp!'�F�^"o$$"r
_�Y=�������'��)�XOr�����`'�H#3~���U7&��\Q��z�'��>���ϋ�b����Y����#YԲ��i��⋠�u�u����^��������VUW=y�Ϡ8A�r����9YYV�����+�"�8���C�������yS�!���愝�לi�*f�vU�܊@�b8R��+�Y-���2A�ڟ�Xj�F����zpW�RX�����E6h��l��=�nڊT-`��|o�e��ez�/0�[�%%%�9��L���t���*���2�V������y-�IG�ť}�N�c�O�F������/��>_�|
-�_��А	�2!�22��=�	��n�=�mݍ�5(JQdU�.#����I�r�{�#�9�Σ�x~��	��,@d�ǤD��zZAN�3����������G�1ފ�2d���-���v����5r�u����MP�E~�Oډ�?
����N�#�݆������]p+%�X�,/�������TS�=M���
@p۰�q�EAU�g��&7�M^^>K����2�����_�,P��K:*T{1���Ç���)))q����5�������?=�p������	Tf?Ƚ3�_2
���hAr�QW����#�����ص����X��������Q����F`}`�<j���-������&{�XCSɚO�cT熉�y�[M�h f���Kƫ�w�� +�2����f�%�s���R�Z����(��SEqT�3A/D-��H�M1Z����r�u}�G|�"{��%u���gFbg���Gw����M�h������i�Z�n�ö��SL�?���|rz_Z�Ҳ��)hx7�Wy�`��Ƙ��##�N..�k-��Y�����/<褔+��7H�@H����=���LD���|vO�^�w�wy`f��q	��F���]Ȇ	9�w��-�rv�8�w2��,��QO��n�h��oҼd�6=Pb:D$��f��9$��$aA&L ���z��c��"����S}��.8�*-��j�-��LLV�Pl�������ޠ���<F��	�T��:uL�!Ï����g�f���V��j��,�m�7e;�i�F�333Kϙ�95�!wq9?�G��C* L� ^L�2���\���nD޹o�0r����*�@���;�{�3�:�b>�e�����ʀQ�ʨ	�޷s�w��0��d}Di� A��<E/�!�E�!p)!ezj
)Yd��>�m����q"�+����������g���9��uy�eぶ���?@VB��sz�6��L�t˚���G�]���A�L�u^�eĳT�{y�Y�^�mz���R6$�9��?N��6�|7���R6eYn�gw�NZ������M��@I�2G=�����>̌q�Z`13J����}X��S�>��mYl�6�.���ċ%�� s�����{o~��R`X���CYn��TQd��A�](6u����.{�h>*cg�=�J�{j�o��)G3W׌�o�VnRZ9���Ӽqe"�}7Mپ3�q���'���=�L�J5����;qh��o�k�|��	�������P�+�puՂ��^���6���*1�Ť�#{�����+�O�W��o��iqW�=�L%�A�y�b$��b!dupQ��v��{gԺ�.7�E��{ڝ��H6v,�Tȗ`�[����n�A��h��]�١q�j��w�pOZ?�$��g��^�[tC��a���}���69�n�������tx�DƔ����9�f�^�2|3��j��[��Q�<V��>��G(�2}��<����¢׆e�� �׍���~\��m������&w�f:w��]��{+�o߿_��{ �]��%}����S������|�V��2k�^��S���d���r�V��O�S�E�*������^iۯn����.��X}ek��=p����~j˧āCD�P��N��~ԡ�P�&��t�gO'����D[�ۯ=�hٽ�����45�O#xJ�tĊĖI�Ǐ��t��u��a��s`�5���7[�y���W������Q��Z�XWZ��Ӿx���0�!K��x�����|<=�����&��)��Yk�%r��%�q�Se�7E_}���HP=���Fߗ
��ӷEm��V�������I�b�#�y�4�Cw���o/�X�4�R*i�ׁ�;��Y��H��ȧ$Yn�9R�5Y���^J���o��3g��5�DFvh��M����15�Z�?��|�c�m�� ���soǷQMee�>[}�MBr�f�&>^o��{[G�w����t��$����ނ'11qt�ǹ�v>�۷;���)��yxZ��T�[���{v�7��J��貀�鎃fBǋ��zS�<j3�l�}W��%z4�va��/��:�7��O^y��5LȚa��^�?��|���TOXx����p��p�7�inN���$w���|ģ���4��54��1)�~���ӡ����C�^�tH1o�r~G��i��<f�r���7Y�H��gEv�E�n_lcL�ZJ�����$�n{�|n;���ܼi��%vq�#{��~78OH���q{o�/�H<�5��td�����W��_3��~���}�Q��	3&�eY�5�~�$�8�|��	��k~���J〟9��m���UEDc����W���������?�T�-a&4s)V6�#�7t�5LgЬP���&-��f���֊=)�бG-�?�<��3���Y1(��n����m������e�
�p�r��s�'��=<8�3(&33��������K�z�||�C�,�q��س�|."�R3�O��9~���QX�Ya�'<M��Oc����g�,g�;��Jw�9gn);38x�V�M�p�����~����j�)��,C3�n��1�$�3#_'6Ϭ��&��֮y)O�N���@V�՟F��b� =�~� ;�^�cn�H�:C�6(`��������� �/�B��n��((:���RC�C�Bm�Z����b&�юU&%��sñ*Ԥd�Jen�#�ee�-,�k����>�����x��sٯ��{�2������y�u^>�d�f�
�:	-���"��E�
�b���E.nn���ZCG�������u,�����lN���BB�,�?"�I���Q$�:�WI��^�ɖ��s䟉|~���w���.�
��v�w�i�w»�ˑ�1��#�N�(g��uƈ�m��	HH�x�RK�ƨܼY��}
,#���o/������g�og���A��6��v�rMH���W�Ep>�*RY~\��>��CrRz�"�a������No�J0H�hCv�Ԩ)�yY٦�an���g�޽�����fY昹�Z*˰�Z��(&���y?�y�@�:��Z |��Q�&1��|RGA�~�p����Z����'��@.����P���N���@/��b���r+=s���@��������x��]�R��x0�{,e��V���9A�Ӏ���Gz�{-1�����*��V�JZ��������?�1�6(����x��ϥy�F���/� ���;��0�fBUR'�VEaG��,�}���I��w����E4���D�_�hI�La�ȜY�"��m���u36���ϐvXŧ��4��{�b��#7�;���?�7ND�k��hjI&W���-�ѽ��[���I��	�l��K���f2x��]�y�4��K����Z_bL]��=��1��dxee�8۵0lic/�\�1�!_�^�o&ًmmO�4�l.�!�q��:,#[�����ޞ��R��(���܏�.6�c ���n�U�LJ~����œ/�ki�ڞ���Fj��Z܊k�ԗ�xrS)�jRx�36�Ѹ鷵���nxj��U�54�v�%�/��Tn�Fe��ӗ�(��\���7��ך]/Կ�`1��u�X����w�o�~|��&�����k ��ॎO��О�yp]�qK	hT�O�ߓ�\��s�2���^X𙙥\�yb�B���ƈs���G�F��E���et[c�/K�=w���1Gr}�H��>�V�����S=�p��"����	��cimt٢̽,�U���B��k�L�������a{��������"x� �*�t^$m�y�9~2*��SCj� 	ʅ�~�
G1@"��uޭ���?''�!��mL������i�������q�4�������5x���z"d�A����q��C��Y��ߍ[�T	޾����޸Al�  ��!��n�̰T�j���HLy0p���˞���u ��eއ������r��8�x�C-d��H]t�a��fc�! �/V}3g��SH�y�c>9��2��ޛ5n��}w��7�
�jHV�w\|A=���s���>W��n@����3lwo�4"�n����}��Q<��ɓ���o[;;��k&���F�[�bk������W���~=�eK��6��Na���&pvu�����F���^Ʊ�����+Jm�}m���!T�qlᮣ#G��MF����Ǻ�}?m��t^�_�A��!���Ioh�8p8Vz�ܛ^_�x�78�����h7��$�'��?A���P��>�<���-��we�%�bv�"��
�������~�i�6�z�잣�A/Gᤎ;ƾ��t��%_m��+��,��|7,w���F�ł��r�ذf������ě���1%8�SJ���]��--��#��0�)+;��y fP��tP%��oa�g����ҊG��4X�n�ڻ�����.��T��Afp���U&���W�PT�7�t*���fW�f�W��ܛgW���@8������	�,m�E�苇;ǟ?� �me̪��𫍛���I"�ˡC�����6MO\\Kmn{��������ya&%��:"{�����|��B�>	_��;0�t��Y^���L)�T&~ϣ:z���D�\��3.7,�g;~�}���mR���Ǘ��h�f74�)����o���N��P~��nΡMsҿ��b��{�,J�&c�ڄ9H�#�8��0�2#Y�?�?����y?|H��ᘻ�m-�Z�@;�IӔy����;n�ftE���4��ue���q�{�oѤ�r�\ �K��Y��@�f�P�26O޿�x��|'�	OП�]]�2\O���z\���{�贸v���H�!��u�H:��y���+@u�	_��>P�9e�O��s����/���	V�3Au���+��|D����j�<��,�O���fЭ��)���ƬE�06ߕ�t�2ɷ>Jr����v$y[J,M���.r��k��A�ϟ����ʮJ�D�k��T�P�+�Q�c����>H�U��~�@o{�FG��eT�����3/y��t�3��u>}�.�s!�����.g��۷�G��0+>ZvG�����4�����xr�Pv�p�~P �Y�o!V��q��9~e�¢C�l.5d�=���U�l��⚬j.��'�;�т٦��5 ć�K�|�y���_(1�8z��;g3�s���(�G{y����(3,V���l�&��\q�~)��6�-*�� �<ls6*M���xƳ9���z*��:��K�ΰ3Y,���_�fH��py�}����>�<��	W]�������:��F�֎0���#�i��}�^erc�f�V���m�Ko'ڮ���؂#�y�H2p��z���^9�y4�x�ax���W�%u��R�}4;{闇1]\����33�ۍ�Y�[�ۭӷn*�?�~yY�*�2zW��"Χ:�A����$Z�n�h�wc�_���y���$nA�0��ks�;�NI �C�ɦ��޽{��A� ������S I�ըy�ϻ"���d�����v����y0�$���_M|]�E	,t�n�?�afBa�t�dOT���c�c�9�t"Z:jvVW���:�2%���a��1��n���X4��9�-��i�j���;l��QTt�e��\�X�h����q1���;O�w��"4��z���!w���4��Ю3gΰ�4���b%@����h{�@�&�8�}��,9t��aө{�7����z.�eq
?�y�e���x�����h$"�5D�	���D�����cbN(�����V��!�	c/x�Tx/$�������S�XE3!BʲߦZ�":��C<�c�<�u���>���2�yi�*ZV{��F����ҡj�����)��s Mi'/Yݿ��Q�O�!�W��jI��4[!�׭�?�������W	edeoB:���HBfFd�ʖ�Yd��|#�!��:I�W���������o���ܼ���z>�������z���a�%�B >�۲����P�s� �,� !<���6�].H�/�a-���D?&���t�$'#�@��X;8���+�������������թgOk���LM��ξV��ә�t*�����ވ�~w4XY����f0�S&o�C=;WV�|�����n݂b����fnn��^�3;3��Һdh3h��8hd�U��z ��0@Ɖ��`���++Hk�]�mo�m�(��B��R�o�v�ѣ9���=�B���qh������S�z�iJ.g���}� U�J?ԣo����tV343���~L%�thH_�����f���Q����C�#uѱu�;�`0~EV���{'��~[�2ַߤi
�/�֌Y:sPZA�Ze�4���x
 8}�+�G��_Q�uw�8nke�=����/w5+���X�u�ӕ5��9V����rJ�
d��_'�re�KH���$����f� 7�bx[0�o��X�m��=_��܇Ů��o�w�z{*��X�D@u����#诤:�ܔ	z��a�NK9@R��}V�"��M"��K��'�P�_q��J��&�x)$-��U��+3W���'q�j���9��a�3�]� '����g�ɕޙq��r�{�j`c�M��Ж�`�G�NWrWj�#�i��\*!!��@s6���==�GF�o�U�&]]��L_���G�3��@%�0��Ě��b�,p���i��{�Er�l��E�R��II?�[zWS��e@�4�(6��I�8R��$�?�Er��ru(W	2������Z�}Qq�`���Q���!��7(�P�*�ŴM���ݮև�z�G�1��Ύ?	�.G��!�1�_�O,��଴>Fs�H�� �C%���ɱ��)���2��,��� ?>X���a����;��������i�N�8@��v-+s����]�����5��ۍ�Vo������~Ŝ�Jӗ/ܴ�r�q]*��˼���""�k���P����n�EtN�⡖�`��}����R���?� Ӡs�)R^�>9��C?�Һ'D"1������m�MNe^�&�A�!�����ӓH:�x����Պ�ʮG�4jQ�3M�^��+�6L\�Z��w��A�k������� ��c��}�r>>[?�ǂx�n�ä{ֺģآ���@(�l3(���1�� M�M�|������Z9+�T���1?���[l�j�Uhϡ�L�Y�h.�<��{�I��'NU(�Nr���X;���%%E0YР'����J�/Ts����Q��5���8G�I����B!���({�ʡ���%��ALq�5rC�a��T�5�&�0��A����G��"�o���ᰥ(�k�1o��GoK<�L�Fw�8�n���\�%"ϵ��ԩ����mw߁e��l�!�0�z��ήT��gB&:3D>>����oz	&�g��BCgr�\'	n�TgQUE�֧��2F5���CN�葶7��&�̖WP@���P�d%+��Dx
���z�����R�;��{��ȯ��Fړ��АL��̮G{��z/

�n����om�����C�� ��͍��d)�Q ����r���lePP T��fQ�<�v���)����n�L��p���c��&�W:	a��n�6(w���"���U�ԭ��ͼNL��Z�=����k��
�+5=;��&姅��_z�D��Fcc���,����3���47W��]��NQ���i�&���KL>��i�9��o�iOOv8ԞԠ�/x��Ƃ�`�1�c��j�i�ő�w�~`�@��Q�N[��}��z�8�v֓=Q�����
�EA�'�pm�$edex���f��H,A�Z�ܸ���s ʟ�ΐ�N��#�:�n���}�'�����JJ��[����5m}���i~���~SSww�۷��~C~�SɕX'=`�Q��ï��U{�������>�뇠�d�����re�ژ�$�&4T�2���oj:ALӥ�<����c��!i�Ew�z�%��g3��Amm׵�[�Œ�x�d�5r^ۀ_J�K	9����=���R{'�������5n�<G����+s�Lu_9��wx*�
wG^^^XT�d�;���C߀:��E��u����.��#-��3�c5x�=��}9!a����
��ָL`j�M��<%�ׯ_��tjA0�uo_nϪ��Zh���f�#�񀋋�u=�x�wM*��%z3�ޏ ,S���߬Ӭ��*�KIO/(��C�,�p�P�y⌜Q�VO��M+�vVQ��_W�}�4z=""⿁hC�@)111�B��k�!G��9���.*ڀ�	���*� U��Qg<��F�j��o���n���X�w������Q����!A�0�߿�(�[�z�=O\�p�m�!M3J�S�� P�%_F��[/gJ����r��w��hv�}xH޽�L�!����78����cܜ����K���!%
x��u@߼��Ȫ�bpp�I��c7�i[��";��J�J��p�~�qe�s���t0�]����hy�,E*��_2���'Cg�������#u�����;��Z��3�N�H���٥�9��6�$�I�2Pdsϑ�RB�QE�R�7�����b��Ĵ[���L�l׀�ba�x���u���Z����,F�\�|5w�E��ő �_0k '�%��I@nu��� H����SS�2�%��[�Y8�|J������n��q��j$~�n�/�w���j?u�1��NZ���(o�U
���ׯۜ�;j��N%''�ӑR��#<�0��f��#;f�뛍h�M��ؔnUt�lgn��,��f�?޶��j_<%�D~�>8O�[����iJ�~/Ýә�������[�3��g��3@�v���'�|�B6��hÖ)'�����������b�٠HǝN��yҟ�����,��w��x��2;ղ�{Ɩ�Tz�����/��i_����ĉ<t�UKo,�`��h0���?Y�N�0i���6p�@�M޸��BT�����뢂�<ؽ�V@,�IE���V�j9B2rrS''����+��**�>�Ds`/��'B��&b�Iy��H�
����Éd|8��$O�(�����w�.P�CQ	ķo�Z�L�K?ϯ�<�'��^��Q317gM���Qm��6��JΚC�����~h�(��H�W2�x�@�� ݫ��� '��ۤ�	�A(�$'�t��֟����9�R�x^���6H�?�00��0�!�(��?�{{�.���UU'?On�Y�Y��蘵
�ڊ1���.:��gUqG�-OQ0q��g~��C{���kQƣ�R��(v�e��*�K�Ǐ�.ɼ����)���#��e)
9v�u�I��EJL���6+�>#g��#""J��PZp�<w�*\��ל�����erP�r1ErQ�J:Y��X!饜�*��>9�UQ��M�=<�Z�̫���� ^4�D�u�e)���gdp�'�L�L�"E��f�~Sܺ|�������*�?�
'��xv�d��|ae���0�\+�Q��<�/��E{\/c,�F�WԔ�7$�E��a�I���@|k��qs0��D=������{�	"��w��l.�KSQ��Cm���K��b�v)�5\��{b��z��靝WIw���=z�?8�X~�Z�8��@��"�'/'W� g�٨H?Aֿj�o�OT6a�Pd��-�/��䱛"Lv�ަ�������]C�FC2���P�f��*R���K<r�q�7������.�m�[W ���P�O�^��>>�,Y�f�����g�I����~f��I#D�A���8\^�t��Om��`�D�Ɔ�-w~�Bssw!aa��"�o��8��%R�BB���N���G��F5�k���Y�5�=��JJ�<~e!��
p��j�a��	�Y���_�6⏸T�^DTk�0������4��/#)��cU��E����122���ʽ������Ķ���Pu�d>$�������0c�3-�P4�3A�J��䖷�׎�����^��T"۔Z�l�RR���V��yc��o���_K�K3PQ*Q�I��g�4v��u��^ryj��uF�٫=�L���F%��ؚĳ�'�#�ﮪy\\&�����Vc������o��_�������s_BZ�etTP�bָ��� Ț�M	��q��!3�)i��\y�O���d�L�\��z�ӂ@i��ݫiBr���2�&�Zװ��jkq�81 _�B��5C�㿝�#,��x�7�H�`�T���?O�ò�(�>���ϺT�4B�HE�i+Mt}�a��tI��IIo�ּ
��-=�~9��_O����`�f���z�n�߇�BC�6%���s&wL���k�NhV	s�Bx��Urr0���ZZ���6ށ1jn���&�r�8�/��{��{_?sTo�����<���#��
׳&"�Y�YyA�s���R�K���~o���h���|-	z�]T���9�>jjj�jjN4	!R�˓U_�*HBx�b�[����'��2�i��pӅ�dM8��a��;����ij	�'7�F+=�43���&����dEN�=�_���b��T R�H�g��xm�}s��=#W���P6�Mn��p�ۖɕ����Zڈ�/
C�8��y��𡰄�EA�Q�DWV��ŬF&?���͝�RX �<<|C�5��g��3(K]c2߻�+��ݎ��l��v��ݔbk�����Sl��{��鿺J(.|�o~���ޞ�-:7�1�b@K��󒷽��t<�N�j��?/,�H����i�g���q����pV0h��j��H{s��Y���uI��⫢/�ZO�C�_�D��mF<�op֞��PH�� �u�GR,@���Y_-/��,U������8!�}**�i�7���w��d�Z�����������3��753�y?�M\��c���n��}�Qׯ#�l�� ���e�G�O��/ܚ��m�iz�\K �[*x}l}q��D��5"Г�����xx`u��F�c���f�Agu9J0�f��h(��ޤD�0E����P�eQ�w�����l��oo�����0���R�mW��kN՟��%
i;)�%�쯎�#ћj��^U��#橋o ��qI������.���iC�az�����U����[���tD	9FfQ܍��j}0
{�հ�O/;�84v��adѭy�Ԑ~�,V���f��ǠN��&6}�b�@��ɤ�-|�Z��`O5x[𧪻�E`L~��FDF�����5�.O��E	b	��� A�� )�����ڜ��~��J0�ˋ�����*28<�z�3z}]��Z48V�2֒�ΝM*2"�^��i]cc�kT�G;��K���_{�Z��N��Z树^Xڷ�G>�E��R]�)k��?�U>T%�_u|$S@sae�6_���f�ձ���;��G�ѥ���BBB$zuk�CdM7 �p8M���pӀ!8Az�"at+�t�A#;;�X@'M�����5&?��Űuc��Y�<a����maL�PJ�Sa����s�r�k��'�ĎTz�'�?�<N�+VZD$��n���r����1/��dj�<sڐ��l��a��iM%w
*���a�݆�&���[�!I�8X(L-,���$����o>2�04\�ܶ���-cX��)��?��H"��o�{my�~��izU�|���k׆Xx��	e?����؋o2�.}�	TxӉ��A��0�$)�@���h�e횅�����D�"liD��hO�����3~�彈bS��߹s�$xA�2=5�MJQ�>��Ī�&C�B���W�
k�Y���ۭ�n�չ�b�}@���~1d��?����BO�}b"&���yo�,mTT��iWrZaa�И����g�f�^�l�E
;+��@:N���5��H�S�P�oݯ��#����c�t���+���,���<D���U�^nؔ|�w[1�yv����빹|@�Ǔ��� ]�p*n�:�UG-,����_{��Ɨ�.\�1G��'��g0ۓv~�74;�/��]�{�$�)�LE߫���ZC���"�#9H��7��W˻i {�d�7�5�v�w�d}�@��L�T�O��$%%��'��<h�?��-�~$��X3&�'��-����& :_k�訓�Y׸y��_�J�͕Z#w~Ʈ^BY��vui@i�X��c�t����Z�)R~R�}~p��X��P>==�@%����6L�̃��⡶�fU��S��0���h'wN/o	'C=T�}�ܔaÍi�Y�#���w�Vn[<���/���˽����V������!��6qq̏�������1�OU���Pf� <���]OIy�)�>V��k���11T(��ё\���G������m�g�n&�R'Xfh	�\[�E�Ʋa~�&m���f,a gDDD���:�@�B�1>9V�{R�������\��i��6����Z�),��9r0�&$��	͚ ��KQ��}���������,$��"�z�֙���NwD	N�qE0.*�b%��0ٚ=!�4�ޟ��qt���!���Ujj 
[�b2����7���}�#�ݜ��f�++�
�z���א-~J9��GdYY�IRmӫRR7$S���C��>����N�`����j�iT�NIi��yU8hVr;��f_�H�!���[g�R�S�QeJ�w�CP�r���v֋�n�K�
W�>�m�c]�4��iҞ�\�'�^��_����7 �f�|�=_��c2&^��-���TUUA�L��Ry����op<�j���ڜ�2E��� ru������m;;����0��#�h�	J�*�)j�i��J}�G����7�-e+��;�}��suk;�]}���� &�a��Y�-�� ������C��]5$6L�l3+�� �Δ��T/!`6�7�)pq~># D��f�]���
ٱ�##`�`T~�@[,�VLݳ"`��� ݛVy�0�ys(A(,"��%��E�Z�h��T�B�Fy�X48J�Vő�\����M1l�{1��wE�2ńU�4^��XI�9
?՟��J͹i��r��/]��&u�{����J���A��ƺ�[�0�:�i��� ���L��o⽺ T�**����L.g&����8�7�35o���
���ne��0�'G��/H��)EZ�����1�(̤��*��Bd'���%d�$@���Y���1� �[�}�E:&��hB�L~e\�8��pexE�LBa���!�0P�Q���Fk�fO��~�C��sΝ��5��?[x�}a�""�)a��@x_�����p>��)Wד�D2&��'aP�`e���r��Rr�����Prۃ+BdYr���3����ԡW��U$x�7o3�=|L k:�*��EV�0��h�У��}3��,l�į���N�?����[��"��'�:{N.�$K�0v5��@���8͇��N����^kvC����Ca^��Ҍ���%�%�7�||�ݥ=[\�����+n�������8A"p����)(Î)'S2pM/��K�7eh	�ZH���:£�2>΁`��ǝ��Ut�HG6���r����ֲ��A�"˃tt�Bt�R������V�H>×ܞ2��rRc�[^��־��7��S<�fL���a��g�O�/��v7\^ZV���R�7��J�7L,��hl1�&���,ٯ���DȡB�%7�Bj�}�Kd]���u⑾84ױ����O`�a�˻'*�f��
�y���lk������3/��Iyo1�H�QR]���$t�8�Gcd���I ���r����9�7$3��w����Xv��S�`����;*�3���w(��p��"���o"��2d@��5z!����8o��n�D��@����i�26��w�g����yWU��V�'���%��`�N�Ğ�3ɓ����E�,��ڟ��|��L){��{�%� H��f�s�-c�n��=��t�����5���k�VY�`��C9^KM�3sq�%�U�־L6٤��V�Z\��̴�u���޹g�z�n=/�?���1�긿9*�օ��:.��1	a���p)
���TW�E�b,�9xӒ��༏�ET�G1��>7X���-���0�����ݖ�8s|���Q�)�`�(���-�|�mz�EYXY�p?����A50P����\���N�#ǲ����說�������]�!'kzt�2W��9����;���ڜȈ����BQ��['N������Ρ(����&�'���$k@� :��rP��Ʀ@!���s�I�JP�i~}�H3_D�ךۯ6�P���SE��J&X�[L��z~U,�)`	Tb����&�L�̀	m3�,ņв]jņA�Q����f���<fܯ4��V�Ūh��*'L��TL�k>7[���ih�w2E���j�$��6Y�	�7v,���p�{�����_uuQZaM�k�!��SNFq
<�w�=G,z��B���7ksČ������rmꇐ����Z��?	b��% �Pd=es�G�K����������H�U6�R��,\s5�
�Mlө��/S��/��lū,��a(���TK�*�Qة�*S��]��)xWR���6O���>8���J_���fY�Nv��f�cӬ*��M�s�K��iO���щ��x��0G+K	��@�j[ �.�U����ﶴ.�����ih#q��O��"���ϻ����s{�G�w��B��1�9����O9��%������>��Bl��8�M�[�������f�?�wo�Bp��_n�>�fh�.�kH��KD+(���W�sNUM�|7h� �8Y���*�U���R��WB<�m$Y���q�������?9��ҲxC���8�@���j�ӑ��A"?�1%���9NEjo�x�2��a$�7";��mٲ.$b�XH+ҹ��3aq���H�sT�iݓ�D���h����l	p�m�,����^QY������8�T�+�2T���������� �[�8#�<�g}B��#�h�����
�����}]�����Z����+Sɩ{� F&'i�v�]R��?�U���������Г�� ΰ�:Q�|��gqq�,ll�B]���О�ɬ�����Y��{6m�KNNn���7;H���ӈsa�"�X�X�8[W��\%�QV�$�x�c�r� ͅ<��U�k��'�D�6�o����!��s������A�<�Pup�(.ʹ��L���P��͏SDP�Z��К�}�I�#�O�s��_�z�O�|��e�e�VI$�{}�.�<�2�I�p<����{ך[
K	��W��`���L�������(eS���qZW?Q�GZ��%0d�F_W|��/ ���J���/��fWa.��뾱r�kt���ĺ'�R�S�|�VW�P�c�e?��7+��IY���,�LJ.����PE��!�~`P˽�������P���n^E>��bᑑ�R>����ݍϑ�'k�!��4;+�U3�/�	,;1aJp�y$?p٩��+��gv.:���� |1;�i�y(O�I���#������|-�XH/6�H����(�y���|^y��J���ᚡ�����N��Յ/.��A$�#��W�)	�vtI�yC� W�f�jО\]'	n��{�=���[����p��ӭ#5�Tћ��ڨ78F)��f���w�&�(2��4�^sO�ܟq�w�`��i���5�Gv�H��4��TWW��(˧�໕�*�iB����>Mf	��F��o�dJ��9����;Z��/��d��Xk�6#��/,�K��!���w�1E��fQ�dA#&�#Z)�����ץ�Ɇ�NJ�~�8�4����\L�{�����4 <2�;��F	�p����җ���qy�G�|\U5J��ob��h��%
��d``xn�ğx��M��9@!�Ӟ�W񺁠8q����@MY���kj��~��{|���aw�͊�Kv�s���2�/��P~5y�:����2�'�8n<�#|E��#�����󏍇��T�a]+#օ��\��[�z��K�ꍳ�ڤ[��f�ÌoX��;���$�U�?�9��V��yu�G��}��u(r�R���{>�2�ݿS#���=��4)g�3�̦�a�=%�������[R�o_��okm�t�D@������ͦ�4�k��榦��2u1�*4���%����_��2�4�����~{$��B�;?(D#��i]��\L��������㓧c
~Q�x�U����"��nP���9;*�~�Q��N��!�����V��ˤ,�։���Ndiha�/��~�Q.��G�X_{��Rbv��"�뗘�7e�>s4&'�� 5	��%>74�"c��n��y��K<n�]^�k����\�еk��X��V��%p�H�Pu���s�L��ڻ\�W��6S��+F��MSH#����e�j.%Y���%R��dr/��_����
��Q[W]�˳��YH�6!���$,	���-Rl&?�g�wԁ:�WGQ32Z�{����w�[����ǀ_�Uv�33��d�ls�j�
_��_)�b��.)�K��]؞ק��9Ԩ�1y����f3]}}d�LD��S�֛���;9�+e��\}�"��tpp���'Z�t<��`w�#�tz����|�bz�h�v��A��%8���c0�]	)�r6�u�`hy���T�A��pJ�� �|ᙯ�Ț\����aIXq����	�↛;~�ylс�^�ecg7uw�mͣ��
<yG���5�h3Ҡ�S.��&&&�01���a�N]�����J�{��=�B�0.���U���-?����meo��%6�7'+Y�Vn��Z�Ą~B�y�Ӻ���ǯcbR*�~zzv�D�T������|����  ({~'8�W"U�{��q �BX/ �)ϭwȮD���(���7jjj%ee#;�=n@�X�渋Qu�r�HI�!��W��ʨq��X��gώ)t�
Z��F�W&��^�t����V���� �S�Xs���%�*p�n�%Oת�Ɖ�(�j&R��0o00/:h�k���;�o+�!�V]�ٌ��,��=$Ğ'���E޴��P����+�����3U�;�L����)���4��PUV�ΙB����&��G6ҽ�
���F�bH�F����W�������D��_������Y&�=�-�@D�YkU�F����c-ܡ���x0��r��b;��#��}Vw<�(�`� ٶR�J�X��������Urr�k^~��i�)v�H�<k�Dl��O{jM���U#�~�:U�������m�����d����w���,�?�"�(��+6碨
:�!���~s��b�����I�����Y\k�����Β��RR�����Ƴq�+����^2f+-��{�URۃ+W��9eՀ���#�h�V"�B�ND���IY��;=�	GB�����aqQ�f����E�~ݳ��J���R]Bc�d��\(��~`�Zf�L[��N����^`���ž�a�\�+[�ω&c����@ϟ?/��跢���p�U�V�d���2W��m�Bs=��.���2�(�z50?�<�桴1o\KK���G	t��S�1�+f���z��-�����C�%##^�d�ݒ����� d�ܮ��L�H������X!��)��:��i��{UZ940z��KetO��pŀm�\u]��6n�Qo��Y�����'V�;P��[+.h��\�eVƖ�5��$X��:9��9��o��wٲ0�T�Q���*b������ܯ����N����IG@.�����<0�̭Bdo@x�sʾ�fB�][����L�X��t���>�6I�Ut+�����5U�!���~��[�`�_|��AKE�r�� Pm�U�᭣
�G����o��ZÔ����OB+�J����M"Yt�l��%w�T�A$������LD�f���A�)��gl��)�*<������RʕLL^�?5�	��t�MRjj$���(�P������N�:��201�7M���4]�e�K�Zj�� �R��tc�->��<S��LyK���I����,H]���"�U���v��N��T�Q���4u8��N(���5���y㽟�Bn���d�x�����M���y�����6�>�~��`E�������ӌp�	�������>�:M���_���i\Z�b`O�9]ӽ��3�~�A�9R��W<}>x��Lक़�4�݀`��>2G��h�JY��i<><�`Y/>{��ԓ�I:6�=�0�����G:Y{&��9�|ؿ��A�wK�L�����{7��zV�uN����K�ld��7�9kw����#p��!�4���ء�%OO��GN�/Zq�j����a�1�B������z�� =������{_C�����4�>�2�����AI�Y\|�ך����+��W�[���O�[0^V�98R��52e��m�ኩ���`0�!�u��,�����Y%Ţ��dM[�G�k�G������F���s�t�{�&!�J�g~�FBJ
o�/kЖ|�`aUj�ˍ��������p�����^��?�֢�˹;������@a��w�o���0��K�d�t��G��D%J#_*¼Xҁ��e�Z��*wzg���sK�Z�+:KC����:}���c��C��8�h��|-j`;Wz�R���])$$'�2���LS\�ڭ��ëN�J�WY��3IC���+�{o��Vfse&ɉ2ٸ�G� s?檃��s�i%���)�>��:����/�{k�$99YHE�Q�0<����|09{�R6���9��s|#�-�t���DT�����Y�X2��mB8E� ^PL��?#x�rq�2X����c��*�O�Zy�۫1�$�����ln�9=?���2KG���%��I�G-E1�����m�� �X����t��Nw��T�kkٿ4	�����
���`̬f��|�=q"H��%
$@�-4Kُ�9g;�wt f��S���2m��[:@���7E�a�3�;����&W~�.Z��ҋ�x������ Y���_� ��>5#I_���o ��x�9
�_&�/���mtO�2�L �	*w��U5jT�%؋�J�b)��(s�8}=���}M͵���Y$:KWVN����^Q�A^��g� �0�(��7�`"/'ssW>O���e������B��Z^�>�|���,3ٛ�Ib�++`q�.E�	����v�<���9Y���E��9'@G
7Mؘ@�	�	���}�;/�@5�����>��չ��L�֔�\0<�"NB^�PMqT.�����o�[B���U22;��Vp龍v�B=�.�;N��,,T�l6]H���\�,���%w�������9}�4�;$��K_�&q�x�D9VRQfuM���[0�Ohl��+�11���
G9޸����JJ���/䢻�9]��$�y�(CK���~�.�P�?-F~u
�;5U-1ND[N�1�Ի���15�_B*�$E��A�W9Of}+�[�LML��x�IoGEG#ۊIy���ee�	֛n�]�J�#l>x�#l�2����e�����j�N5#�b�}�P 1`����D�
�<Ea)	���d)�
�$/9¸x=��n�?v��[q6��jlu����
Nzu��-������&I-~W2��[��((Ƹ3u���J30א�U��>wf�KR�9����9�0�(��ԕ+�$�M	s*�O?~�fv=�jU�(����E�$]c�[(:�'�\�F�οS��T�2���<}u
-�R��[C�=u������㩚�A��wO�޿�������R0�]�kdg�?&|kD��K |�3�z����ۨ��~��m� ��(���
˼���F�ˉ�g�����i�}�����S�
ى�"Y�ˣ��ߓ?�Df�����z;�rUG�.0�����jt�?X:�Lڭq��˝����b�*��C�Ρ��NG܄�iP���=�����>��k�֐�ly ?�|����L�+�~;T�lj5f�o��Ö|�X_b����q�����iU�}W��d`����upW��p�몴�Zj��-�~�ڊ�7��-Av�~�zE�b/$K�F�V�����ΐ��^*�'�Tdv+���p��ޘ��N@�=o..d�0 �+{d���}������DG΍���ͭ�uT
&V&o�Ӆ���^�P�&�����P{���Z݋�9����uv^ս_�W�p}a�`��������b̋c���^��ddff&�h�0�0��ں���m�J�\O
b^�\JBf�"*)),��&�I9��T�����v#4M+�� ����,��M���1�ŗUh���+Mi7y��vL�́:U�K
P�+����a����j��D�tiְq�J!d�{҉�Z����uk��BH�ޛ�p����hv�V�����.����!�^s1��#j�wpITelJ����|�L@&?8�2����C~ Vk�Ό;U����;��HzR�=�Pҭ�}�w�:j}]�'��l�0j(H�11C	�j�	Pqkj�J����{�3�'?ٻ�����˴�y���徛�k��%��{�%���_���P��m��M������n�3N�N!���C�.=�����q_�T���O˃i6�p��s?~;]�{�R�������',N�~?ZC�9ȴ��Lx������{9i�Du��K\��.HM~�a0�OF葵�[2���0�f�k_�� ��F�MKq[HX�X�B�fI���ْ�� �0R���Ȏ#��#��O;�ږ'�������_ݝ�ZF��ji7��L�,�?�������t��*��>opӳ�fKl�I�)��f�����^EX��	d��NPu��f�
�5?'@�~���'8
s�,E�ݠ�[k�E���z���S/����z��s��pRB����i׽����߃6Y��!���C/;Z_��%�X6�OQ��OQE�wģ8�"U�I�t���f�:|��g������g$�n�AY(}���@�P��m�ߢg&���Z�-:y2���aۃ�yYC��3lR�޿���V_?��^�r�c6�2�G����H{G_Z���D,q�UXb���'��[�^����hkʨr��(kk[�B�+$�Z��Ϟ2���ݒw�Hc/���]�M��l��p��$�=kGj�Uy:.��i������V5`?��ӀT3+	1+yz7>Cnf���J�uE����؃��֡�v�J����;�<_�}�-���kk���-�\��<	;��Ɓ]Oפ��x���}G��.OI82�D�{�I�#8Ů�k�Y �U�����R5�g���-�w,��0!'
==.#����	_�妺֨�GTU=	��m�8�l�?l0�b�C����g���.�����|*����J0�l�`")�}%i��ݽh�+&e��"!2��&!2��c�}�ID"*�&uz[�;c�K%��ȋ�VSI��5�P>���Eޞz�ڸ���ޱS/x���[�+���x�ض7|���X�I2uEfaĆk������raaa��9��7{�P����<0�{�sB�6�ԕZ�ʣ��
;s���i4����݀O��%`�~�Ђ�D�L�[�X����:��1�e�K��Ho�
��@!�zټ͊�σ�L�)�O|��:�o��;z{?1$��� ���QH�gĳnF��Ֆ����z�1��)������\��v�C3�Q�ìˉT
���T���z���Q�Z]��^����K��^�QB�q����v\1v��|�q0����%+#W���2�ӑ�M�'�!o<��XH�c�; @�?�"�,jbcC�l�q�=/��%o�v��R�Z[S.��:i�I<�\8�st�>�f�+6��'uk�~�"�7�d����WiR`�9
Uq�n'FK`k�uL*�-��[4=�9z�����iik ��p��w��DT�,.|Xoȳ�VVQ1�j0�LmY\;}R���Jp���	��̈t����\�]�B� �o���۔��Xe��/3�Zn�\�������~{
���gq�6]�u9�$�3������7���8� �7*���Iz������Wii%C���xh��녪PRR�:�b���<��",$Ͻ��c��࿷�֒��]�)v�M���L�M�>kv�����[k��K`�<���l.�<��q@�$������%c����yQUn�&�9���?
c����hK��?z9�@#���:���Y��[��2쳰M"��89�4���5���	@��ĘӞ�.�&K���n��.�R����݀V��F�޵B���Z+��WR�T{�n5'���H�n����ӂ�'
*]&��o:�1�4D��ol�ܓ_����\X�
؂<*yK�+sy0D�P���hf|؎΋]υ�O"������E��4
�G�M�`�"o��4~�<m�𻶥��&c<rԞ���	yx1cSΤs�^?�M� N�cҾR�%��&�bh�!��|+�W%o��Ċ�A�B���`"\��;#��g��_`0���Y��:JJWؒ_z3���J�b�9+�}몭\s��44q�<�<����9`�f��d��������h�꓁z_3����q ��A� `��-�x�NZ� ���sH�<���C�=���A��tc��M��ֱ�������Aϖ���Ť�]�jЂ�<cT\lo���勦��(�{���vv�Q��,߾��+ѵ}|y�(,��̌��g��=p����p,t �O����dv�k�r�Så��{���ϔөx��3��$��80�.�]c�
�IU���\�� �wrЦ2o \��ݳ�h�۱<�U��_�.CU{�tN�eTu�}kwwiv�>��=�6�}CB������!�w���O���_gP���$�V�9v��iy��g% �����Y��Q�MNղ�Sh�ƽ=)���;Pj�����#�n��ɴ��e�'�=�'j�����iVV��s�O9H%Sӭ�G�
zN�2E�a͍��n�n/,����BN§`�j�v�:R�P��q�^`�cBޮxH�JJz6�`�����U��k}QA~D^[%(���Ţ�QNCe-)�e��,������)3Z�4A���)�����ހ�Q9V�:W��"�}��zj�>�6G��;X3ť���W����)�ݣ�r�"��C� z����>��L�nIC"��r��du�{�H]��+>�M1v|�sL�W�4�z;]��:?���Y\F�z��ߩ��Q�o�x�{ҵ��"9�����'B>`����H� �/7D��丼��$pGHf����k��CZ'/*���s��[�>{r)>�l�u/���c	�~��h�
���<싽�| ��+�48#y��1����H�S��d������9��Vie)�;d��~C|�Io3����KQ�?{&ո���
XwS:��L�<_O6��f�%5��}���e�\ͮO����������t�������������s��iO�M;�M9AQ��m���V<ݟ�+.	~a�b˳��Թ��ͺ��ע~�T�No�p�bzv�	s��?l�9/���Ae�d���\J�����Ks�����'�i�ro 4$d�+8�Ril�6@�6ޜx{�Kct��JQ2]"vۥI��罗'ʡ�JJz����C@os|u���G2�c��� O�V�8�(��O��,�?��������i�8��&��RP�z�r�|���N�좲�Z�����I��w�[���2���������MrO����n�u�i6}��Q:7��)�Rf�$�(�������f��B����@�?n�A̩�h$�՝u��� ��D�?G{���7c�^0�t9�{Pf�$����(ɱ�ߣ`}G��}A#���NU{}��ma���;W�6����&j�O:��t��">#�^$才�Ç����� �����U���{K���-Bv�^�++�쑄�����G2��d����������x����]�z��y��|����z�^��~�n�z��|�&�n�	3t���1�5X
F��:�ʊU��Z]w㤉��ׁ7:8�A�l��Ħ)s���B|= *���(S�)5L��K�{�j.�ӏ������Y>3�s���؛JcE-����~Qo3wy���@`4�8w�V�n��ߵ�ˠ)�7�����)�-��,��7���УZ�0�P��]fH�Z��ĤOGB�㍍����Juuu@�H������^���?����1�:����������{�P l���C��21���mDZ4�R2�c�T_���r'U:w���|nre��r�*Z�O��:N�Q��.�R\�R*��"�á����l"��?ɾѴkl�{xE?>YN�̌̑,Hs�1��Y�W��uz�6���I̿C�wR�:"��h���v�.�Y�`��Ĥ�l�- S�( �x3�g~�L�#��:�����Z8c�b����'�C�����%�p� �TEm���~�O��X
��@
 �ڥ��4L�-y����g R�t��K`�9`�%ec�E��\�gh���sd�]� ��V��ɯ����.X� ��9�����]=��5D�>����t]���߱��.����|�-�睹����MMW��j'bq�s��Vō=$�H���2���=�.���s=�<H�wmep��������eD2DB��� ��,�h�/��/���|��f8L ��i?����sp(G���+d���E�����
���D�>o��������#�/�p��P�o�0?⣩���e�����ѝ�w��Kγ]3���hXb��뗙�Tʿ��XY�nk��@�NG�+)MA��fhFWhjd��"^��T���ى�i���@'H>��L-�Ő�{$,(�����Y�k��+(��������9Z>}zeii���
:	�A�������!pQ11@�y���vx]U�NI�.�w�ir̇��tO�n�hVd����҈T��֥����ۇ�[��q֓_Cer�2�8ȗ���J:��t***�?�5)���A�%�s���γ�h5�11�6����2�p��g� �ˠ����a��틍-1Ƌ�-��U]���D�n`�y�2��e���q�I�����������e͑)�H�ȆD(��َh�Y¶����Z�^�׋p�Ċr`T��_&LuV<�./���sJ��1E�����D��(��`�s�amړE�,4L�8S�8���r����#��@Ɖ,L��̸?��n� �����IZ�?;H����t��N�#*�N�>��\ %���aEjP��ѷ�m;��R~2J[��V(a��jE�6���L��3ۊN�À��],E�]�T?���?���z�M��t���Uw���j����ը����Ǉ:>���f���=V��5:Jm+�-B׊���/��)o���E��郗%�T��t
\�� $�z�#*��s����bO���u㖇��6��_3�r̦VaajC��"V|����q�	uuw��,r��31=�K�\k��H�s&7���	����EsQ����0���N	:��
�.H�r�X�께p��UņO��y��~��j� ��T�FJ�������X�k�[���Wę�ݼ/��������oO�Ggq��8�L��1��s�����Z��>C������0��[����i�������HA@�R���?�`��Բ��/ǆ���H1 �Y}_}o���(��G	JK���dJ�@�0�����C>��>0,����VP`����'7����n�<G�"x�7u�ʣ�.y`��|p/�����S� &��vw8�OGsdg��
vyXuC�K96m�ޅ{%(}4�;V���9 H���)�#�@Pҡ|���P��������{h셜TF���9���/����{�1�Dl�g>O��v��>'�}޳`�H)�{K�`@��Sr@8_�۷o�B���A譭�wX/񫫠3 ���O���X?���gO/�_��G��.c0U�!�:�=��tm��S�y�<g���3��\��@:�&*hiYH-y�"��뜡����K2�;O�	5���!|24� G�邎�,x��0e�����������]��܈9�OI�Y�_{<=b2[�z�}. 	�'Ř(�y�����@�2&Vf��F?w"��g}��#Ihxy�7Q���U���|����z��]��V���;�#-}������y
�����ҝ����/��(��Y��j�@�ͳC�&�].M��EеB
wSJ�,�ISFF^i*0?T`�ghs����t���pqO�0��!k��o�j�X�8��|�����Wn �l����C���F����'�9L�=>�À�y5��~�%Z���j��rmn��?�9u�T飒����d�>(~55QA23���f�eq�f����c�HY���[�]���o`�cx�[�������x�sV����:�Toan����^���(D��	kc��I�+�i�
:���e��S}��a�߾���Qκ�du�r$bS�w�CUaӽ�^��j ��o�;�&s�ҦL�E��\n]'������k;�&��mqqq��|�f���Κ�׮�KI9��8I�'�Y�?<�h�:����*����W ��mYY�!oj�� ?+�ٷ���)S4ظ���e@@�YR��@:r��1� qdnsI����%G-�����TW�vxz�*N�H���2!/��e�C9*��n�̨���\��o_��dk��L���)���ze+�ƭ���Έm��s������?�����(���L��O�?~�n�	{�
et �Q6���޴��9/���'���B��A��y�noo���B��LrJ;�@��!�����؆�M�����	�{6����D��G
�Ϸ����J�k'�sMinj
��/�Л+)�N\l���!�"����<���!7)fcCX����,@����S��1%7~��↳G(X�_��U���f[���²�.8b�Y���@.i�\[4܀=������2){��>&��Z��EEٮ9��s���p��s��n�a��-�dR��ӿ����gv�˟��E���Y$��r�L���|}�**�D���7&4�u��^��Qʊs�����6���_�;��.i�\�$�ɕ�_��NOO�9a��@���M	ـqS�h���V�89��H�W��=������u�J[�/��G��Xn�?Y��g�X���_�[xV)�}@􆷵�!|������!�:l�6(=�Ur�O=�x�N(+�@}
�6N�am���3Y%=K�s�熬J�f������F(C��Kե�L5`���Y�V�=!w�	�����ɻQ��_��?�Q0y�����4�W�ݸ�z�\k�Kd7�E�wnu���8�{e)�#KJn�]),����;B���:��s�HQN1*丢�b��*Љ�/��&�&m��7�"'�j����!�b��߁�����w�o�鲇ؕ�%K�bOU�ggy �1�=rx^�Z	���f+������.�-�"���m��w��BC[��=E

0k�캟����}�����,8j��-l0�G��5��Y��h�	��)-�P���bL�ܹ��w���bw������"G��1�8=�����)�Db��{��
(�ܘ��g�2��+qW��h���� ^�ҒΛޅ"Y��$��Ç�iԽ�ː���TR�%WWW��Z���Z�FG_� Q�,�!\�9��OZ�x���Z��v4.���f�y5z����{d>Ϲz�%�X�Cك�kq#)q�!gu�m	B:p�l���x���4P��-�ꅚ=%�xע���OꌡD@�#E	�Qv�O��������x��.����l���ɉ��f~��D3���P�j똚�jk�l�*9y�b��<oj��Ѓ���Ҭ�g)S���! �0�}�h&�����F|�O��z~���<��sl[KGx���5F��Up�+�5�7o��¨U��Ռ���@]X�<5/`�8)r<�7�B��|��.��'�:?Y�}�u:�%;�� ���@��O�~�6�K�!��J�i�D*7��t��uZ��˅
?�'�}�ś	TT�l\Vpێ�2L�	�7�4ܜ��n���;���ə�z��I1�4���H<h��4�XQ�xQ&�W�T�����KP�G������ӱ�F�}ij�E/l?�XU���$
�LYF~4+9"�m����ש�C���a'��0���0�e,��R�@�4�`)@ɾ�E�d���'9�|�h0��������øn��:P�����5���%;/�oM=ܽ�\��^�Z���	ʼ��pq�2�{�;?o������d-䟋B����%qiX-&�D�; �͓C��=�$��xr�}^j�5&ff�-�^?�����)��Y��r�T|P�Ql��O�K�(�ݿ��'��Н�V6�μB<�n���W"r���=VA�yC/x��W���a���9/�)+k����oғ��	j�
y�	���Ŷ��^L��(��`���o��6��rx#-Sje;�(���/4�6���\������I�tOL����HJ>il���D��AN��QEy�\\\�R����:���C@ְ3��U�1�8�3���&U#��S"�]��<ćG�Ľͺ�Q[88�B�s�ѱ���j+v�{g	2���m�uHȥ<�o��{{�Z�e��I�$ht~�wA�]��z"m>u���1�$�rݸ�����Ѕ�̡�;ZP<L̄������f㈿������_Q9�x叕��]�h	��Э #����o��gM�>��S�#-}�8���:�{su�P�К��ܸ�Ljo��8*Zu֫��g��1RN�yv�|�ghx�B�^oz�w�{2���i��%s����*=�����\���c��<(a �A�!��=��/���x�0yP���fi�(#S,R~)�	����{��A�c{9���xP�/xe%���A6���>f���%~��I�U�K+��M�J:�!�I�����z�LHXCO�/Z�9�V}%Y����������}y�.�cඉ��oK��G;w9��y�fd����\LA�k%ā|!**��4:kx�̄;EE�A�ϷI�#�Y�� �i	}_�v#VTx����g��HZ`�@���G����J��ϟa�9 �̮a��z�����W������h��M~*�S=/��	5�<y�2Ug�N�,�C��vB�5���w��(��*�U0|�pʯ������w�
>�ss����N-���hW��[{�sp|�����6@�d�tKg��E{��Ւ#^���<�m������{�A;;_QU��4�$ޜ����aw�:&��z�êo��$*�E���_��L�����HP���&�!ߑ!��Z�*��aO\�ґe��k�"��'�G��\~���^���G#yR�x�ī�3�8��S�Hz��R�a��Bj�H�O��E��~�T�K�Ջ���>h I���B����9�w(��x��'������E�؝�
���:)t���	�s���D�+?��f��IJ��cl��V�� �^\ģ��V���ua�����_T=�
��l�Ƌ���0�|.ךxv&�Ńx���r����t���P'����&t�8�������'� ��)q_���KA�'��	�̄���D��P&��1�����Y.01�$� ����X�T��@�OZ���@�ƂB^��	��B�99n�Ԏ�2��hDs��A5����,,����~w���-$�� �蠂�w��K��.x��?����=E��wx8��TTJ�xW@R���5�l[KT��ݦº�����F^��Ew"�oP����^T��L���?;���/��q�ܛ����B^&W�T�IO!�uś�%��4z~R�@��
��l���Y����<VHA�u���_�{��YJ\v��EɦS��TgζbW���:Y����*j�`�����nH�R��Ֆ߸K�ᠽ(ݧ�����Hԩ�m�{t$��m��������I�-�?wvh�%|2���Q'�ez����	��4�d�֯��p	0.P[�c�XR��Pyue,Ql�vC3Eo_JhB�j*�{���s&��G�O�~9��w�`6��UVH��a��<w���G>F����:E���Vx���FY�03��R�֖p�^���b������)7�nF���G�k���#��#�e:;7A�0��n�ʌ�+�������K�Mh������6KJ�&W��Ս��@�R}�̮ޘ�|��8[��m�QW�;��/�7P�j�R��1�-���t���'�7,ͷ��PlZ�Џ)r��~�>ˊ.����/2ά�M	7ZA�+W�\�E����=��0ZͮRSR��R։"F�JbM��.\�"q���4�s=we�z�&�����q�řĦ��y~���aG�*��8h��٩�oG#c��7u��?�(}����f�ۺ''� �$U�v��&����yNr{D�!NN?ad�?�Q��CT��������φ<w[[�n/h��@]t�7W������[^�T&���1C�t(�t��n��w�束�N�p=���d�4��iK�Á�����Ev��]@�鹽nA�gٚ�GLb�6�4[��9��&~��u}��p%^-�����N�q	�X����`e�V#������o���W`��ga�����[��geq���<4��\d��	Vnn���6��wh�`�`�y�� ��*����B��,=��,�r4���r���b����s��>��XҋI�Ƨ��G�� ��x#��9մ��+��h�N,DCHo�wB�n���4�-���������=yش��qh�;d�o$I���c�x��t�dE����j���E�:��TA��^ ��+���-O by�RI:F���a�Z�|�:�;�4����)ǯ�z�����p�q����PQE61�6y5�b0������Ǹ�:낤�ʭ�,\�8����Q'!�8�K�l�
h>��N��F��8��vu�<�quv������.G���Ø]��Գ�'
G�Eu ���DD'�o�>:�y|�ʚ�g_]S�����Vi���VWwwMuuDM͝o��5��fA�T�뤯�()��/н9��C��y2�G�����h�D�p�e�?0+�H��dH� ��q���P��0����G󾚽���wY�x/�s��Wز�ڗ���;�^���m�Y *o_>`��>����0�Ɨ���汍&���i�ts�����<�
����\t��*{>鵴�G�Y"���������z�k�>� ��8ƫ~�q��x�B�U�:��[�K��"{��MZfO��w�݋<<�
��Q��Qо��uLO���c�Ѫ@�;���s�I���+2��ױ``!��(�/4�8�R .֦�x�$�����b���̜��P���Vl����i�j[*������EZ�55
�H���r��^�ٻ��载A�T�Y��Q�zE3�m����!�3��o"���2��2@C�@R�K?��B�� r�_�;�����H;;j�ܭOn�:�_���!�G::��\_�20�ii�Q����b����`z�ID��&��g�	^��\4�ZOC�wG&�$O�5 ����� ��$B��a���m"hl�r�jn��T�����?� p��ws�AyGG6�Jd8U�x�Q�|q����XQ1�1*Yl����s�.p[�����Z�8�`x�ocZ��J�f�f�}���h:65�e(�	}���Tͺ�N��=��e�R����bȚ�~�i����Qi��ʗ��
�����+�́%��d]óm@"����H���rw���Iq	�2Y+��K��
EYRF��{5~�^�+��{�s���j�x���;��"�bG�X\%���%g�Z���h�za;�>������+����F�
]2Ck��OשB�����d�၀шB�8�!0,��B}�]����.������ʇ�C[^��[�_��(���ߖ9�*�-EC��Q++�H��<'�WQ�*%����
t��(�?�:	�*:9�`u"s�\K"�kqQ�1��9���}�]��ZKׂ��d��ß�y�������먃o�_Zg*]P V�v�gz�u�<���w���yh���2a�G��<Y}���lt��Z�x�~��*�>̇A����:�{l�AJ���61��{l�?x{��$�Fz�U@����ʧ$��۬eͫ1���4,Nva׆ �v�5h;=&��tИY[�c�t��@݊���T��ɓ,J^k_\P&��Z��׬���q?�&���%���?�#%��	͝L֣Ňn����\wuo�5�E]U"���ż9��LIDe�>���~�)M2Whk��%@X� ye���;Z!��N(�2�\�����p�{#�%�0WUt�̌Q)�B�dk�X���[�Fme�H�����A:��?��J�q��� $Oͯa3��l��ͽ~N��������Vw�t�1�r~)�����b�N|��cc�Z..�:��4x�0��蹎�<��uV�aa�noϟ��QR�����ܼ�%� }TZZϵ	$:�P� �9	 D�R���0���v����~���knS;��b��]|�������1a�d7��Cc|��R4Ԃ����G��򱧨e�y%0��d���bç�m
�-��������&z7K c�4b���3�H*8ӡ��r����Q7�+W�FTW� S���q�/n�|2����,��������q� �yFF�ی�q�y�z���.�Жu��#�����/��<��V̝��<�>��)�@��0Q%�0%�{��i��w���I��aj�g؇��̢�f���v�:�ƴ��;'�Ko-��.��/e�#'3���TC�
�\���Z>���1*��c��9�?�
�Nf/N|�2��Z�x��tR$v�'��EM�.-�9��Ң\7��CŁ��b�!A"@��KM�������?y2���j��]f!���DD����X4��a�J%W&��G@�1r!N�2;
LU�.z��v��OX��2�j�+��jddb�Ax�[ª�|}W7�TX��Q��Jx���E��x@�a��7�[l�M@�k���1	-x���Qҏ�^A��g� ���[��4u	>9U�?��oX�o�x����Q9��4u^6����	\����9��PK�,s��8��B3�]��Һ�e��Y�0ց�TnS�"�ؔ������q|-���'�/J���6]�&@��[$�sf�	JЌ@F��]��� L������akg�R*4�5���	�#�Y ^ �D��tg��)q�"P�����u�q/��u`�yp�g�����`�+���ˏ`Dި_�L�����P��慙Y�c���%P�#5Q���Dًh������h���Λs~�_GA2R����p]�OrC͞��tdk������ݦ�\Dkjj�����1�VϞ5V�<y�����L��-M�LbjjS���h����cq�� H. !T5���ڄ5@	���|=��M��� eحS/KI���e|?����t��WG>Ua�z$Q��Lͫ����&�Zf� ���F*�S�J�ms�oǈ�k3FB=����U��0 ĺ�~�Wq����>G���d(�����>%x~�>�	�L�&Y�
�� Y�#5��0tJ�/���._B"�����QR�5��}��vu6��i�g�-���'4�"��dXnecCr(Z���#��6?�U�	�b���`����^��i�S�$��NQ�M<�BS{b���t���?.����,�٫"��\�7�p��	rl�5�I��_�H� u���{��T > gi�l\_�܀<V�� �i@�h@�h~��P�Λ�� 6/f�%�%��6�w��VD_#c�
8�NM�,h�s	bN�t�-Q==7� j��;]J�ƢY$�����T���,���u]�a�� d޹��nm;U�=1!�G�����0H�gte��Md�,)9).-=���b�rH:U�ݺ��_��>{EaEA:�f��glf&��X��ơn���^�!a������y4IGŻ��+]�/>a���[=���/ŏ�b!���B�ZOL�Q|%���*��CHJ0_�J�h�w�UQ�2E�XBF��9�ZN:o���h���ޅ�߿��HV�k�OM�y���}42k&�F��ٔ귃2P�DB �Ld��˄�In�J4@�ҦU�^625���P��<(+������6� �b-�<|}���s_7��IZ����,?��c���^P����^��TvX۔�/�o�o��_���>~�B�`rn��N��h�6���� �#�w�U�Q����' h.�U�5*:Xri�� ãY=��N	Y^�(��#R� Y�Ȉq}�*� WXH��,�� l���&
�a "f��`��� ��z��`3���o߾Ex�֕M ��������_��q%�yO<y��Բ�] 2@��j�����a++��s�Y����m@y9ڊ�
tD����sZ�a9uH(H��Ľ��OzEi�y�h�b�c�Z!��u�j��}&�Ӡ�uD��Ec*1�'�E�Y�"fXo��r��R��ffe9;����_
��EsF��0c0���k�W�Z�@F]P SSS
�"p��j�7PPL,�Q��$�@>�yKH$�I�u����7�t7����￢���X�B�$���>{�_ݣ��C"����P��Y�#��J�Tu*B��i� %�1n��=Rj�'�@��5![c���|.���E�V�Qˋv��5_U��Q�\�ʚ[�5���;� �a�r��!�8"�1"��CE�DGWyz{�*p >.�����14k�I��~�%���#�;��������mݸ���&�@���1�VUu�&�]D{o�B������}vv�m�)f�^�\܍�zg4��a�e�|���b��������ݥ�*9��s�Aa��!*��z�
�J����`7o*x���yW�-� �K�hBh(�m�{es �#�{�~�P#��:K(r�3�E�
QE��B�U
�0<J;�������3�=W�{p��]�����Fr���K**H����ﴶ122
���G�A����Xb��5ו�ݮ��5wZj��[[��P�;HIE���� 8OVO*��à�����q.2E��ꌅ|p��>�jS�Y��3dv�\�3y$�%/�p���-P�~Q[)�z��ǘ�& 5��ԯw�n4���7��.��2��\�D�ݯik�{f~g�A���M�AC�$����Y>{��qٽ��f��v��-�v)G��{�������M�G8[[S��g�O�24,SZzG�u>���b��7EԜ^`!�:..�5Ů���-d�R�Qb�u�4b*+t����a���@:(Q��A�1��)b�/{?����¸N뚒�m-6�\������a�	��Ɔ��g|>~bwx]�]J����K�NDq�u�\Hb�x��\jG�� ��X_X~��X�߮c�J��`#*����n��h�WJ����d+Ɋ�N:0
�x�b "%�졻���T�7C~/�)ll4�Ѕ��s�ܙ)rd�z���"0X��|��Q4�~1
@�wAӨxZ.��< ��� ?�Wq����+$s!�@��{��l.���U䢸�$�����d�a�H�I4�l ���U_I}���%a/%�d �������xibn��t��g���=�Z������l��[�Aosr��n/�nA�p���u{�y�����-�э�h���\��5��B����/�y����4�{��&��V�9>�$-�8	p�� X�Y�{C�z�.5!@!OBd�/P0$���:�������'���b�}A�l4���4���v�`H�{��9�7[� ��T�� 1Y��rfX�D��8�9�o� ������1�R�(+;zo�7մ#��'�d����Ҡ�y7����ܺե9DHS�d���b.���&?+�$�sJ�;�g�
����jj�hCZZ*���ڀB��H\  ��\��?�=����z��z��b2 c��k�'�]E�C����dH��� �ygY3�0œ�v���hp �ᢈ���e���g�.��+�CENy����e�LJ۠�*�|��ue������!�)��Z3�і�>أ/���8)�˂7߾�W����8\X-+�,8�
�����X`��/6�T�SҎ�x⌌�#']Q�X�.ba���?���0�ǻ�&��3O����
��)U��SJ��ӝܮ<w��ڢޱԑGB�(Y�h<T�<$̪�]��oc='���䩔��~��6�",����H�{)O?��=�'��+�ͬ�Vl���u&@̓�-.^H��xp�?��B0�Z2[���ʛؕ������c�8R7�A�]�I2�J.��
'�G�T�YԎ%���'�hs�q���32"�
���;�5?Y��"��Ġ�T�d����{|; ���]�L=(��7�/���7�L�t��i�NO��7(;z�Cf�y��s Aк���L�t"f6TA�����2�E*����i7T<ծBa7�:���hq��龶��ћW��؆�nˌ8�wD��߄O�;ՇyeT(	Kx������k����_�8��Do��M��������Wb��?����;�vS�R6M�(,�C.�kp'��?�.�ך5���[+���֣#aqf�9�z�M*\!'77�,���S�-&�K�C����d���OH�6���>��b^����zǦFq����C��_��R�s��f�A2��+T�d����| ��dfib�����l��D@�dr�,���]�Z��W�9Z5����Gr?m�t���P�A��{e�Nkr���Zh����o�H<*���_�Aߘ�l�*���A  X����|�'��u����}D;�Ho��j��]��<�r[<�@MKK�M�/W�>/� �3���_��6]����g��D4(�����A�(�J=i�a���^�?e���,�a���~MS8σd��������Ө7��'("PS�ޡ'�q_A��p�,w�����<���]V 	!i����A����5��X�4ܠ��o��%�РC��ڪK�>o��	jb�;����M�ȺQ&W�&�����m�K�擗�����bT$��q++�?���^~A_�D�����}A��2�Vv��U6L�!�9g�Z�|9YX��yR��z��ˇ�::b�d�_.���iॿ��p�<�H���{�w��S@�:���.+�v;M,�~�\Nظ�0�s$��!��UN���&��u}�E�=�8HRM�U��B4�!w �uFrR2����o�G e_X��=!��6�V��Z��{�H)+��rzZ�իi��?�Ԉ����q%\�%�]$edځL� �[B�A����p�d��������r�{�Nf���e�.I��hL����G�I(��j���>���1�MBA�_̄����F�T]���bE1Ȥ�q��>gı�ˈ�7\+ڨO���@��[R�_�z�r<�w�sUmN���Ag��|^�:- ���d��B7�>O�?UI��X9��;�Ź�t������
:1y�[Vf�=�/��q�n�r,ad�+�����Z�������$�m���D{���Y�˷�_C[�|6.|� �d��޼�K�	�&n[cK����3.(�
h?`9�t.P��*Ε<�,��x�`ÿ|��,�^y��P5�GN���s�Ms�����A�7ڡ�OZի�p/e���)�a2c>��3V���j\�:q!H�:E�埰V8-�� � ��z���'��d��E]uu�}��Z�~��h:t�Y��Xbjj�Q��e�33w٩}�y��b[�˿��<}z�P�,+ͩ�]%�C�k�76����zl�V��:��� �����ꇦ��Ŧ߶�=8����j�A��Ukv��
ex�)�<���]��n,U���
i�@V�Fӆ�sv%c�{���,E�|H�x6��)�l����( ��!�#�ҟ���D��n��>�<a�v���7�Q����w���2�;h#=�[�?�-��h�*�K�������T�7���\�Z}}}�L���6����1�6�KGǫy�%G^�/ww�A�C��[�gϨ�,K���쏏�x��!Si�[�q���E��oH3����X
Fh��j�A�k��є��~{Mc,�<�<AE�|ԟT���/7�l�'��i�d6���n�]�Do5M��L���?�ȉQ�y���wx�|d�}�Hd�\�]�� �ey����*��y^Z��4��b��]�%�e��Q)����aL���{�SY?�5�B2+9���w���}�إ2u��Ʊ��V�=�����z��Ւ_��6m��.m�sq������l@楥� U�Y*�WW�/. ��W)�5p�鱥�mBV�۝���d�F����.3T�׽�IE�(������7��|��D"GE�.����xɫ�Wc�ZO�Y��%@;H��̀����R;Q������Ap�
�&&7@u>8��`e�G���쨏4��pZx��Z��e������P R-�ˏa=��RL��kC�`�Gp��b��R|������̏3��-+�(f��VV�=��11�V;�
mڥ�NA7�B���8(1`�@�-7���jRl~�F�&_�R����R`'�O��vE��	�AL�E5����� � �F\��(M��q��7A���f�`��DL?a���]���r���Ce��ޅ����؞��饋��,��g�8�_ �_�я:-�����[�>�4�ǀ�%<{aw����e���Mc�2 � �t�����_�ܹ���zw?�;�;���T�k�QiDx��+޿ק����ո�|��L쐀W���-��b�����gg2�_��
��u!U�z�7���hv�~��q�O����+�~V=Qs*+.�:R�R��t�������CP�+�/埇�;��g]c�+�l3�-��6�w,�Ot�.�$P�77J�Mp��YT`Ra���!SԾn�졁��0�t�\��g��\�Lߵ�*���g�hb�l���x��j�!������ޞoU0?7�2NS]y-َ�oc:����d��������gR,��9�-lm����_�n��w�1p���	1��Y47Z��sjj��P3�֨���VKojf���_��1��[ʠ�a#���,�J�!�Z�X�꣊!���"��Gʈ��S��e�7����*���KM�����b�kh�����i�/3%eJ���>��ۀ���{Ǖ�шh7��� ��M��8�L�Ԕu��<'j���}���L�G��D���ٶ����/��?��O>��W^]_�=U�R�]պ �v&.����W��������bm��=� H	�i)�s�0"���~�=��^�2vqu�HU�ՁFuZ���{�i>��_^�p�a������-�5�T%*��5_$�|��[��px��[gj��k�`���!*3޼�H����2��тJPE �3޾�9J�r��˂��0/(�<%�ϛC�
p~���^6���:�\�L�eM9l�n��H����>A{+7����QT��F��l\�����h�h kfN�*���^��?''E����y"
����Lk�V��~	9-�4:�3�B$�h� ��Iz3C�;q`���
@��}�l���C��b`)�'Εչ^=���2y�.��v@�7�B���*%���D"�k����EN��n���^h <y�U�X�Q�ܢ�Dux�44T�N�6�,�Kf�eB�pA ���yՆ?9���p�0F�"�pf�;�
:w��\����UX�,Z��2��x�d���|] ���?;y��{?@hC�)⿺$�%���C��ޮ��O
Q9ߓ��͔���Q~��dw�-!)a���:h )촮�X�	=>�� B�Y_��]78c�O����Ԥ�Lv�"~��͸ny�#�\�ɔ_�is��oQ��^R�%�+���/����GT��/� �ɇ��P%g}!7��A�`�V�K��N�P*^��O�i)/CL�-$�FM�ݹ5<8�Ü���n@U,AJVS[{��-��J���
�D�9�}�v�vǁ0�Q�H��5)��\_'� p�\J0��=Ϭ)q(��
�{�@�$@ہ�8)���d�	�����9P8%e�F�59��w�G!�����������v�|ȇ9C���� w�FS!R��1
������tt�*�����옟o~��Xˇ�Hˊ�n3)���)v���d���vw4	wv�Ǭe�K���z�162̿���ՙw�q�P(h���̮.�������@v��k��cuc)�^���<9�~L�o �(�P�'����؋R��X0[��5A���\�����2Kо�L٨����6O�5W�%r��Q��w�A�e<�rswV��ꋲ|����b` ���y�t��i��G2��R2����\��E��<�:���1�>�L�j�x>�x���s��sCFN� �}�q��G@6�5�����	{�u熄�S�v����VW�X�m�{2 �`mk�T2k�f�F�+��"B}ȁx{��UÃ�Cd��� dq�Z��/q��:�q�A�S���t�޸B Τ��s"�29�:!-d�
,}�u�7Ksuo��̙f�����0��S#/������'��H���
���xi��	d�z��X[�0t���<���12�����1D����M(��6p �Qm
������&S��e��a�yXN`����s��&AJ����L���Vf��W#�cВ���|i)hkt������Nn˟�o�G~N/d���9=O���Z��^�\ĘY�W��t�r ^��W�A��/:9�:���\P�}�D���m@�Y$o ␉��7s�c��� d	j�&U�O������,�Y�C>�]� �?��RSS��=qIX�犘��5᳏��g�C����ie,0/S��-�w�0�F�EC���О�o��o�UO�&�;)t�6���.�΢,.�sm�73�O�ې��'#��M��1��sUv�gb���@��;�����zpy7���ȫ��6h�1;!zPR鴂�΄dBH�����&���	-��K�V��_J[�Q�d�E�o���(��-�5A-�->�5!kO{�Z���/4���/t��d�ok�,h?��������Vܿ�p��J�^�zk�E��[[��������>D.
�fFF��!/��*Y��ch�Z���GI@���|3a��ܜS�il����>��g������&���hY��>)������34N;�U)�:�V��v[>�ܾ�HK߀�iS�7�-{X�iH����\�@�8K��ѡ��7)��Ҁ	�}7AN]���b������V�F�K���Ž{�z:-�����X[_�1���kfF�PwEK��/��U�8[��OQP >ǚEq��H�ԅ�9��I���X
}���D��d>" �1J�m�0��@���;������uR2�6���Ҕ}[�йq�g��29td�@�����9D��nSn���1�<�Y;%�(�n�	�b��;�q����̜N�g�eN���!`X�R����ѳ2����ii/��V��5�C��y�՛_)���H|�v�ʠ(��f�*�ץ]�E��w�h�0	�<$2U,h[��Y�=���,+�=zKԕ|�V|�妩��=��ɵ=��n��+*�*4�9�̄��o�Ǎ�ߑ�&���i�+��v�}�]��Ɔ睕���nϥ~�OO�����3̄�Q�\}w<����$Tv������QfF���{d&3�C:!������qp̬����~�����qz���z]�s��uߗA*Î_S�2�͝V)��s :G���	Co; ��x���ڸ�� �ǫ�w��y�H'�N�-E�с�#�-�*K�z�=�sʞ���s��N����"X��MOs��U��%YA�
����-��?�9�@׏b섳�:��!��Y�h��{��.V)U���>��T��˭����B�J�	�^���E�_�V�e|�W��=�����G; ��'-䵯�r����.!�3k�r��������Y�vt̼��R��y������/��,vq�{�sT�_CDY�a���è���HVF�����DD� e&`(Pd4$���n``�^W�����Xoq)�*���,+G��wO�D 
Ϝ�FZ+20 ��|h�CS{�G��%��?��|��P�H`��v07�����e�`��y�q�z���<* x|-j'����<��aWWW`�0�78s\*G]%�\�3]%ze~�T�ԉ�f��5��WG�W�z4�.�w7cZA�����c<�Mp��b���9��U(��N�b���������,���/2����?���"�l,�O �L��C ��(��T5&�z��$01����$��Lֹ�(��z:���>�����O��+&;^���'t�d�hbPӗ�6G
�d����H�E���N~�%�<���K����ڳF�s������݅_�A� �E�3�c٢�ed�����[ncS .�ۡH�`�F��D�yD��,X���@�����Ig��=�@�d��߆,�ѯ
4l��6�0v�G��:�ׯ%�uӳ�Z��ǿ�ml�����=��4+���4Ӡ_�r.�{ֹ.�r,��Q�Mi���D���8�VO`�������d)��JM�;��ݯ�W����h|��<3��o�Wֽ���a� �1E�ܼN9\N��0=6�(�����WE/4��]/�]	���f��Oc����p*�.Kʚ�Z��;J)f�>5�jl5|��s��p�mb�sJ@�s��yO(��/�qwR~"O��ʵ��t���I0[�����N�M��B�EDkɩp����j��;lji�
j��z��eceDZ�ԭ�Z6�$�t�{�\�Mu�Wl�^�{x���p#�cq��JI'�������A�2�<Ԣ�$��nݐ>ZIʘ���]n���k�*���ª+��S��CC�f���M���߽k������������#�1`��w�F|-9d)��k�kR��~ڻ�]Ž,w����F�S��C��q������Q�S5��� �k�'�e��hnȾ�a�"��E���'�o�k�����=�sR�a�Z�ǥ���b�g  ���mY��͡� ]��s����p=�O��+��C##�h�FJ4�N�s�K��'���:�4�u�me�DV�7�Ȕ�0�C����@	�������֒�Q5O!ͭ�?,K�n�9e:(�jE)��D�nLq�g�J���q�m��|�|�/����S���/�#a��;W1<:j9;�hE5}>s�>u��oJ��Hx�M�%	��Y
�]_�VY��ATy��8d�]���ZT���sV*���c����\��(�y��y�!x5�;��<�_�+&0HeW��y\vF[
�'^�&Y���ϫgߌ�O�'�Ϗ�U������Ĵ��F
]�W3�Ǥut�b��)_�'@�U��:�4퀽����Z�D�$9t�HʣK@����5�rNE����-7��.jj�VnF?W��2^�����Y��2�v���c�r��e���~:�\�6.��NA���|��٘;��c\�Z�z��AHh��7r���tj�Y�s�.��:�/��#�n���Z�� ���V����=&2_)P��뷉�!��C¤ �b������}'�Jy~�����*?�VTN:n�>���C��8~�%C�)����(oK,�������G
;�F�����%%J�����D���R z���R������-5E@�;H�+FHD���GG�a*-}6����a�`����P3Ƕ����UT�Dw��_�φ�$��x�p��,��x�Ĕ���vg��;/>��`۠��>��Q��\ZUh���w=;�غP��Cj)����w�����i�_��/��!��b�̒\u*�w,ohh��G��am�<3Z��̌u�<>���W(�jf���%*�!z���������+�^�O�&e����O����h���}R�k��QB���+ޒ+ޝ�������GHG�e��c�m/Q�� �^��ݽ(��%�g�ߙ��K��F��t��i����J�Zb��ƀ�^����j 9s�DJ'S���[�Ul�����;Z�ij@��rБ��7�
��������yyfQ�� d.)����s�����ܰ��u('�����9�r� ��D�=M��wW�ր�C���N���@P����`�������e	��C@&-���F���"���^TD�e�)�_g�'�F�9�ח�|����؃W��i�P������#���]^''d�̢�Z�^����]ԟ�an�OPR�� Ds�������ŏ�O
�O}�1P��j��E�;8\[���^{��iG$\C��/5a<�-˻�J��\ިQE1�{�1�����FC�� �fB��?�Rm��~��U��_�wׂ4<�,-8�Qt2KP[�ݻ���Ǜ�y-��j֮�7D��B�Ot��į��D#jk�Uy���E$'�=T����\�zqZ\����j/+Z?A��<k�n�p�9kr��8��ߝ@�Jw���R�ՌM{JL{�M��O���v����J'����is�\��������ݪ�rrbl)T�����;��=�<�ۨ�q�).k| ~����(!��E��=�����Ef�뛘���/7h��}A"��եb���j��'X�(D�:~-2��o��[v����"q�ؙ)�r��I.#��{}}���O��3^���B�~ �KV�&���V�y�0�upw�F � ��+�N�����]^����7#�`JE5�� ��W�KV��\l"^�Aj���r�ו2���b���z�� `�̤M/r���pE�4�j�U/����>a]���6[f:;��ͤ����KM��o���hxX��������2����9Y�;:����T���=;t{��S�����:��9�ǥ������G��\�] ���I~֭hJ�H)s؃ؙn�ݨD�}P�{�)c��ta������l�ݳ���;��{�AK��Nv�41͘��ഇ�<�>�C̈́�%��Tڝ��]<Ƿ9�6���SL�Mm��e<�z������f%�h���A�^�^pչ�~��$�����aj%�V� h�8�v^����խ����Р����|�.�8��d='~ [)�a
d&�7ʇ�f67M:%� ��XT�}q<m�?�	r���j�w��Ϗp����Oaj*��e��D�}�e����?����|q�~�	oڕҥ�5�_��; ҳ������,#��A{Hsf'����\#� p�L�߇�S�}^��]���{�S�9�,L����#�HX<)?$;�QJl�K���fJ�(�|��x@�,�.��_���뿥&����o�8I[�$�2�5�,��E"���48���t�����!�k�������N�X5�^=�K�b֑���V�G��_��g��yeO��Hr�:ryO�m��6���Y��j��;��|����g���+W���Fi��v�&�����E풒N�!���\k��gb��&�7�ꂃ/dkڎr�OO7.��$��╦rrp�5G %��O�*Zo�d���=�A�s�@�F{Z�}�T���㈏RR��Ώ��jν;_�R	#��t�����%�/����)�d~��fNN��n����>16��M�<; %f..DYd���=�E�����&�#��K��H+'���{C� Z|4�AA5.�S��O��+y�P���Ž{�)\�f�A�d����U���	4n��BJ��Lx���EeX�7�~PAԊ!�5�}���	(+P!�J���R��f/�fD<)$q���]5,����6'k�����л������G7ڞ���x�]	��XB/��3xI�?��V�O}�=��I�W-¶��ϟ-K�q�aI�e؟W,uu�c��g��ޑè�:�oN�Ţ��d?W�po��''u����ޙ��B���!�s���%h��4NL��%Le�w��� �X
|DP�R�6���+�K����g�o��V���$������s���8��m0)+9C���
3|�:@OX��Q�J�	�y9���ޅ�I�l_J�NB�kb�FAƦ���v�܀��~q���,Fߧg6	��b#F�u�B��BW���wg*{�#��H�(��x�9�!q�dnD��|h�݀��e�mtTDuÉ姽��.�������$���tJ���`����uꚩ�Օ�EZ� �O/��4Nt~3y:��K�e�0�	��̐3,���Y]'������S��L��D���Ү���'�
���YY���i��N�ȿ|�Ni�_�",)�8O�]\Kt[���G �:~��{�<�B�9�(�*W����@��Z�)}����Y�|�gKo H%'��Po�Vґ�J�$j�{Jdm�(è�L�˦�T�><a�9닅U��Q�EF����޽[�����m_Mc���S;�qеpܿ{��w�� F7��Q^�Zw�j�I�ϟ��&s��P�k}O{����`�rT�=y��J��'��`�X"PDiC��FEE�}^��[(ޜ�M�	�$�ɺ\��>��A�Fh3�\�����u�ե��.*����3�/UL�[F���T/�� �U씁Wj�bWW�So�.|�7�Y��x�E\Q���1DǞ�U����ɑ���D�Y�$yt�q��r�)t.Te�Rﳿ>�6)�	�y��2��\����V�.zջ�!¹��_C����G��N�u�zc<�ؚ�:B*#~1�D���u�4��ܛ޸���,y&t�v����H ��Ԋ��Fj��UK��M8/��m��z��P�r�f⇶ ���ڳ	���>V����^�z���Pm�U3[��0�����f�7�û�1�(�jNr��G\�fC�͎ �z	C�?�����dZ~������=3#o�am���vu���� A��ϟ��ǜ���l�9�3���751Qc���h�}Ë������.	f��^�WK�X*�r�Slp2Ĳ��4�җv�k��4.|�U�w0���R�	m�s��E����2M�7�<�^��e�xZ��YW��O���������	�	�Z��:7/��M��R@:���ȫ���0/��s�*� ����\�(W�= ��k3��t-�wW�FD�% v6����M#�\;~)�/MHٜ˂[7�Br ��I�G��bݩ���Γ���X44s�wה�|w�q0]��]h����\Z����:`�7�g��Q�y�<a��:�WVW7;`����5�Y]ݸw��1�?�<�\c�T�i��K[������P�RE嵐�}|�V���F�J�`*đ����XRSSe����B��q�=Gy���߻׌J���"$�^�%c��gT�k�Ɯޢ��S�YY9�db�eS��JTy]W/��
�����ꪗ3ˇ��~GQM>�+�g&������!��	�1�/Qy�B���h��'47�xRl)�NMo��5��U#�m,�� O[׏��_��M*�P�S� ���b�f��'������hs�3�Z"_�[H�H�M{z��JD��e��D����K�0����fA1!Q��4?/J�(X"y��"W�כ����8����w��t��s�WK�Ͷ��p���^ꋫv!t�� J����H̀|���g�3��&O��ʪ^�}e��8謋�(��J��w��2������ �m�[��k4������$�~�@m�Eb��:;�^~�M_��m��]���畒j1 �E/�a"���5�����c{�tLB��#9S�A�����MDX��JKd�θm;H��Ꚍ� ��o���BL��\��ۯ���ѵ
=��х��!'�UJ�n�M��%f��#pK�b	3�źF���$�4��EF����j����L7#��_�+��Y��Y��2C�^�23�zU 	��HB�t*jx|\N��������ȋh�Hmz��lQ���d� 01[e�SS[�u�O�ҩh�S��[X��ݞ�6�7Vw�9XA@�5y��������1@&�����,��S�+���1d��S_��W�#1�\�0�� _��#E:Br���Ն���W�Q[�h�P�\sy�C}������d$��2Ԥ�z%z����5%7���
 ^tRUR�����Գ���J�g�J��G��1��
���ۻ[�O�;N��������MM���KM}������V;~�Ș#�nm�2����	��qBE4��c��=��3��bFڅ����,�g��v�2Y[[�"+��W�.w��_r�S��J	3��Y�H�?0V[9QkD�>�l�ܤ�_�����kp8CF-.��YW�����ux����"�T�Wr e�W*�}z4���3�=-�z���0���-�gj�&�aT*:���*^`�;�g��E~�E�1�J�:�$���s������"��A���p��KW�r�ХP�?�,_n0ps��'�F�-�1u�G{N�-U�d��}Y��2����"�춸.4�����,d�+
/��/2�H���-z#�����������4s����4��d�/.u< ՚�9�-ѫd�>��j%�Wv��Jr?]�8D��2��+
׺g7͂N����d�m`j���܄
������@�����á�1�d�`ɉ����Kk|����ϝ�ɀ� @9����9
����f����j��2���_�T��ԍoFΨ�^�<41��%[�M����e��8E�t~�p�H�Đ'1�2c����(���	^����ش
�(��Y'm����@�,�W����$�/6���:��KY�e{!��#f6N�sX���ު��us�4������/l��T���@w�1R�;Ȏ��CI����k�8*+zc�I���Ӵ�U�/��(�a�L�K��b�nii�x�L���q�I��f����_�:�j���W�}M��,�K�u���� 7<�~Kk����Y޽{WS�4K=��S�bvM�?���eS"��π[�	�Nr;��#z]�}y�k�u{����k�Y�,���VF|Q�&5wف*P*���0�Y�#�QGu(�(p,p��ͥ:�$��Q�u�C������sl)@w�T��S���U�1A\W:K+svυ����iW3TŽ? \�q�����g��L��ל;��j��E@�[f�Е�]s��
�@ƕW�W��E��{{{�Tz��ַ�����Ls( #Y>�P�\��Y.f��;xH\ZZI!_92�,�����j����Ο1%So���8̒� ]�I9h:K% �djo  y�*���qH�����̄�?�W��L�������S�M���E��x�����a�[<Xu������,����/�lF�䙡���F�pz��*޷�ٷdԸ�HL���k���� ����#}�)R����|���tu�wP��ѕ���⧾g�8�v
z�Ƞ�%H�ߤ4��Z880���{ׇ��[nVY�o ���J��8^�2�444�^�VX��޺k@ I��6U�� �_{���0)�n��
3x�R�,N�)�}F�Hr�TI���Dھ�W(]�b�XϚ�p��S�Ì|v�נ�Y��� #0�zH�T�H�P�eXɁ^P� 4
{�OPr��T��a�zc@�Vx��P�k���Y#��seďZp��w��#1ji{�S�=�AޓrAz���]�ior������`*�$��w��|Ũ�s*ڸ�~ꏗ��f`U�P���j2����g��kD��@*�8�Rș����H�Iw:YY]y�W�d隴EeAL����AH���.�{4���Y�o��RӞ���>Ɇ��5�{��$�X+e�ue�<Jo��w�w�UDop	����_��n�L��VN�p0�0x�`"/
o�7,ႩD��6�Z��$Mm�&*���:�����7�� G��n��t����l��pBҊ!�������0N�bڪ�1J�BI�o�l�R��{�gǾ��I?>��_��l�w��]]���f]]`G�N�n�}#�Z�8E�23�<�Ia9<�Eˇ�i��U���U"��ݎ�\Z�l� ���QB���z�������X ��
��`ޓ����S<Q11v�����99L!-�R���cb����z�^1���E�s��������=�U�l�\��ϟ�����(���t���r�y��3��~(�phg͜��A�O:�Q
9��]T%��
O���mr�Q�E}��E�m��":�4��B0U�:#@��_�Y�yOB�/��i�^
��� ���u��
�#n{�������/�P$�%QWW���,x������YρϚ��ο�#:[#�W~zpB�2{�C������go/|�6&��m�w/�X�Ei����b{4_�S׹�qlL����-5����cY \0�O_ }��zqQ�TT�w*.v ���.7�vhN������89�K%B��qr%��m?�����0C��8Ӹ�X���F��g=���������) �[���	�$2�j�&(���%!
�b��}	ޏ���~? S���0����B���'c��Ն���\�9��l�Ed�M��B��4��Q��V��9��B��.�Doy~�
8=�M��\ڳ��a��$D��x�W}�������45>'�#�kU���j�I��V J�"oQ7���𦚓ఔ���Q	&��dM�w��Ltʟ��4M�̌<����Lq$^6t�ތ66��3�c���j�
��u���¢w�&�բ��]�v��,@������Xh��-�]��O�c�K�(��&OB�ë ���@�E�j��R��כ�ƺyO��h"sx҆����^�\={Y�T-��5�T�$	�_��wY;�t��o>L�-�9�+O����.gȁ��v�=/*'�<��겊?:�z�uP�&��v�6�4mv�vb�t Pϖ���i�����ʥu͂��1��|�_��I�6ϊu�kjP�L1�����m--3}��	hJ��3�%�s �w�û��kLSAp=	aׂ(�&~��S@��=�����j&�2�.�4��P`00((E�U�Ȳ@KFv l~,�]��,u�n�IP���/̵�f�z6�� �:K+A��)���,���S�C}):g���;�{ar�ߌ�����wU�q���⠒ccjܡ�sB��
�cw2����a����m�d�g����wt�b���1O������y�=~�X���.�E�z:��0A�iW�t���X�UGA��Oxq�u����s�����5��#�@$991���.��R��&Vђ� ɡh�w�#�J	������X����(c����@#j�q���[�:�k5ת�W[k *�."���i���(�2Lb`��1v9�Q{D��=�J��W7}��h[����4���)Æ��Y�$%{@W	���/ kUV�����\;�8�sz�$H�S�M���)a�� n9ӳ�?c��,���a��4�ǭ�/ƤN}��)Y޺����'�f7X��r�ۣ��mIIg���]?�^����ҿ���dT�IY�M���Ʌ��n�C�ǲ����z�&\���C'�������	�"�Ȥl�ϟ�qq�!���甾/@�R�Q�mQ�eW��b��nTc뼆[��_��y�o�`�{-ӫ�s^/��)�X�A�æ��������r�έ˓�c��o�Js���HZV��]����P�X"��� �\q�U:A�3亂��8�����u`I�c�%�T��þU/ɚ]�F���1��ͻ�2��M�{�o�OFWi�N�M���c���rp0�8�@}g��� Â��UJ��R��^�����G�<J��Jɡ�K�rN��Vt�������]��[��JF;-��B�f�KK��UI'������^�Lgw������#:�-�A���4���p���E��#�=y�qs#�V�jƦw��{�p��Q �]��t󼜸uje���|qz���%i��NM�oh9]^+X�M�91��H�J�d4�n����Fδ�J��
5�j�d��K�?�	Ϸ�I{�w����8ch4��!N�F�f���m%#�&�h���%�.t0�.�_^fL�%G��/G{gBA�	�ĉ��G#PE�V���e�/55����F.іBỻ���$�|./i	�ј�;���˳EٵU`RD͓vR�q����	ҹ��('�"���;�	%P�|�g鉰��V��+���+���.� �+5Ռ3��7�{2������?}�/q&��]s�R�!��o�*è�@��@7���p����]�`.}�!�|m�M����7#D����B�C�4W�+ot��,VT	҃��K�����vκ}.qN��KJx1`7�,k�;�ag]1W�5@:~o���o�˝!�#�ց���@'m�:������%P���]c	�+Pk�T����MMh�j�d��;wLE蓭�+,R�/{��\�{i��{�6�{�%�"V782X@Ƶ?����Y��p�H�pNp�5�*���Һ�;�P�*V�9�=���'��z�+���\�{P���FQ��4�W���J��f�8�\���*[�jÍ���RiC�Ld�Y��1��ɔ�'A�h[�q��hԜ\v�؉�J���d|���vSQ����0x����l/I�J�'�� �7���BC˚1�X�=�Ajym-���F|��E�	(k�A�����F��zpdr���R�L�?������S0�q��(��͂t�R� 	�w��v��6*�ͬߦ��c'��RȎ:��˱;mh��
�*�DF��C�̓�^����"[5�+Lp۵t�=�����beu{�j����o�r)��@\�D����T��[�,��>	(~�{�2?2�$hR왨/]H�Iy��O�����V@
cؙ��������yD�G�,N��
�A�u��)@H�n�R�M�35���kE9_RI�R^n�b{kuL�'�h^+tu�+C�0貚�565̗���-R<@߃N~D���6v��Y��A}����u�N��hZ�L�3̋�( A�54�|��;���x����r~�QVY�]5���h-[��IǴ+�� ����'Ag�0Nbt$	(+h�f������-��:���?�	1?H���:��I�Fs%�։�޽�9���y�5�B�<�0���o�l�ۜY�c�1�_������C`�;	v_�d��	�b���:L����N<~fd���h^+��K>~~���1������d��}GU������<�
�0T�А�,���ɑO���a9����5�<�-��39F
i�?�Mf��C\J�D��'���/��7h�/���"NuǄ)��M�gĔ����}��	���MӮM��;��d��II"��K�P�4���'#~"�TJ��Cz�`���]�ڎt�q�tU�,b�>/�jÞ|O��&eD� A���J��c�J��9����1Hd�f�D�vG9�9��@B�F����ꢥ�g�m�/e�bT�ΌD4��|(;?/"}�7'�K�*�>'�O�
��ݭ
ޮY���U�5�]]_�G��u��
���:�hRV.�ǡ����O�I'�IF%�� KJV�*����I��=aq�� �JCC����
�>�vzۿ{�b�$.���ϯ��/x�@n�!z9��"'ϼ��:�|���)����բ_���)�a�aT���:gAm+ek��/��>j-��}�͆L�����Z�EP4h�I*�<3�t�2�7�)�K��?|����)���,4,5r�I�lÒ��.��J'�d��k�/d����A>�ABJ&�(��u���oJ4t>��r�S��-�ۺp`�

��l��Et�\�mcly��OO�+��--��?k`xηI/2>A�*s!�?W����,pd�w ��%��ea;����`��@�_	�����R�z��v0�'�2�g��7 �9@�����}��\t�aI����=4�w�L�Z�)tۭU=%lk$�:giR�r�t����Q��^���� ��~M�?N�J@TM�=P����N���)9�`�2�J�/�E��|_��*�HU��*ް�H����ߜu�=��W���}��K�AH�D�ɓ��O��{��"n�Ѕ6N/f�G��ԍ�\�_AۯC̬2@(��S+
������!㳲
 g�~��ʀ�;A����M���w<�֠y� ����$ؽ͙vJh�ʯ����zƑ���mYIO}��E߆��ҟ>⺊f6�=�B=w��O���Ks�7K�PՆ�'����\�j���lEt�Q\����eۚg���L��K���i-t�u89��o^'gKC���'��QhR��L]>�VI��Q#��s��*����Y���p���]ÊlYod���q2�oQ�=e8�ol�i�������]"kxt�fI7��nm��lF������D�ڴ�F���mKSi�}���rZ�,+�{�� 6���]jm]]���Z�{�Ғ�н���������E1���=����������̓���&����>�8nLQV5��4⿊�ȿ����ڻ��	_������'0��fQF�(l�e�=4`j;�|�2 _�L��\u��V��7�`��?ۙ_5,#���GK��i`>����nK�!S}�
���~��3f�Uuu
�-jjjb�g@Kr�L���N���?t�o��F$��A۞��u̹�����&��X�3�QMe�75=���3ڜ�E����=7�Y4��=<���Ws�򂐑��{��)"{����^:�ׁ���.�K"r��1��O�
�\�U���\F�S�eXU���Ǵ�����sRV����X�ձO�ֈ����I7ޔ+I����D�^��5ⷱ:l4,���q�b˯��-������ӛ��v��f=%ж�}˻�%�r�6�.�2_&�-�JZ4������Y(�%v�4� �5�)ʰs����* ���v d��!���H���_�u򵡎����芵��5�k@@��uk�I����@�O�����a����B/@�0��f�q.r?v���y�L��Ռw��L0��?{�����5DTV�r�'Zb`g����&�uW���Y҆��/����Ra�Ѷ��9tx�� Y�p0��hlP�}0,}�&���}:D��+`�̼H� p��l41𡃀  (�O��8�u�(Zߨ(*J*]>���u�؝k;��Z����jP'���u7��殪ި��>���Q�1���QA�9�ތd�Oہ��[�y�i8�%��g�ԯ�*�˟��*�b�~õ�~v���O��#a���%�~7��^Myt�)���	��h��Z��
�h��rt@�&��<iUO�����K���f�\A��us6���e�r�)����0hG�R��EY�}���
��)�[=n�9�Pr��ۮL=�-�QKS�P/U����������}|Y2�z�4��5�\����jG���S.��э� o�:��ù;}�ޝ �:<$�R���3fWɭ���~�tlmQ�m����{M�]{{$	|�w%���7< �~|��"����薋n��1�7����� EL�h��}utn.�@@:��O���G]]s	V���O�� ;��=w�6��XwO�X��@���3U�=�o0?&��A�r��x@�v[�o�p3�f��bgE&U��$(�TE�"@�E�Ղ�Ńm?~�Sc�x �5_-��HlN"�Ư���tLQB�R��)J2�gv��L���y~����nD��Z�����;q���Div�9Jd)I:ksf+p����131���	Sɳ��Ŭ�9����6��R�����)O2��B#~���{�݊G�k��Y�6��!M-�=�,��/*��n�7�Q��J�t6z⵭p���c�=��ҏι8Gռ�i8T?��J	�ȰVφTpM�>��!�
�<[L�!��>)|�t>�
	��fR�پU�ioU��@��ظ�:Z�b�@�ʦ�����B�,L�K@�RC��H_� F�F`߼�腓�oK�2f�yB�Ԏj��/�w�SJɿ ����9<WD�j��"�镕�|�7fa��^(k�V�/��$%z�|K�	 �DEEo���tY
:��%#�Y߳��"%g�k�s@��=��OO_��K��Hr�"p̀���L�]6)s�d7*���D.��n��&����DD�eZ@G��3V�mK��<˖���~�Y_��C<��P�˺2sXF�i`n_�n/�E��5�~���̤���zh�D�b��������#�2ktڭK�9�Op�+4��^�
���r�B���u����o�ju���a�Bi`e����C�����,�U�=pl��]��b����8�<:��.(%��kk���3ZP��d�Ak��
�Ά����X5KY�������S���;9�C���%^�+6�F��P[�̓�X��� ���j:�׻-�$* ���'�(��e��� r�����B���Լi����Tl��Z(�viD�Mz�\���,ʉP����vtX.�'����Ϡ�����4�r��н� ��w��xJ�E�?;_��č-@{�{���=]Yo�!"�Y�yw���}�o,���1��1��� m3Y�ux��}֡F��u��7q&�����1�FcU���y�kk_�ݾM�u�1q�87����«Ԋ�L,��O���x�2�E�O��PA��EYA��6�6!�r��2��|7��K8iѕdN ε~b�/0uW��ڦ/~ʣ�n����a�I��\�����8�L��f�^��Ȳ���tx��6���1����,��6$ض���D͝.fԀ'!W�/0�xS���bY�[<
$8�a�����سT����fM1�E�2l�������
;K0���B\#���B�`��끈|����
G�{��+B�����O.;��X޼�-sTV�u]�eyt��κRh�ӕ�') �P���r�"T����DD�]�}^�*��l3.�k��Aj�fxH���5�2��J�>�d��=�G�!r�g=̗��E^��~�	�Έ0O�0�ZU��]�M����؊¿���k��\��I.��8Ĥ,�W��pa��EOB!�&�������0kP5~Q�iJ���w� �7�C�����G� ?s���Ɵno��;&L��ǎPo�w 6ؠ���(��G�
;�˩DKh����3~5�zxx�zU��N�M�]~�%���~�*W[�m�JRx܎���F�u��)�k�h��@~�u�qp<f��z�[S�8:y��
 �D/����AZ�/ȺD�
�T+��0�T����9+�V���fP�N���!(�+N�޿��wA�+�b��%Y�Zot4������uN
bC�k9Д��v��[N�q������mTuAٔ�s�����tz#<F	����V�<ޡ�!5F�0���ɹ�vA��o�E/�̂�ɳȸGԢ���˳B�� ��~h)��#%�b������F2"Y�
�1�_��_��w����Sʱ�{�����U	C/�>��^Z��F��e�B�{n=��0h��=<9��ZŃ}KU��|Hr_���P�S�Ǳ� <4w���(��i�>�.��V���1H�4Tx�t`��VX@R�je�;H�t�F��J@���ɓ�Jd}�./�P�3�eRȃD�>ϧfݓ;^�g�8I/s�e#U|	���j��}cbbRi�a�<���)jA�#�OO��^k6��al��璒�}K��SU�V�b���g���7VF�Rari[�R�Ƿ7���lI�>�Ft��J�C��/&�G��׾�<d�;���vb��;����E#�9h[@��Xb�A��3�./I���� T#�����.��'M�@ٚ����#�Ts��ۦ���s�`�K���y>�$P���F�Ӛ�7\�:ʜ�@疞6iH�_�W{�)�L�e��^��j���X憢�s�"�V�X<d[���GlTSӞR���w�� .�%���e@�_k�J��\]���M��J�,��ʱo3�,���H)�?�[|�P��&&!����s5y@f�$�#��U��T�S�X�$�3�䣨���?�}  �EL�N��\�����������9�KA�ޭʲ��
�A��|K�<�v&�t�u rY�j�� Do]Y����ir��(|�_u�I}?�ѭ�CF>pN�]avě���	'.���7���/uJr���TY�L�xf	�db����z�2l�����O:���L�4*5P�Pkg��6oEE]�����X�2+B3+�Q?؜L쬷����S�$44��p �O��	^�@#���ϼs8 Z����&�ս�||J�S[{�[m=�$W�]���5�㣩����@���H���1nZ��H��HyP:��E����jH�	��1'a�c2�K������ t�k�P�\U��U��6�:��#����z�^v�3#fSD2P��7�.�P�?��� ��S;�?C�C��KM}̓B�5:��I�/�|h�jWϝq ��S���@I�{qs�߻��j�����cwL���/��܊Z�����ɧ|4@�^m���>�v�!{���m9���w��w�USJH X�|�A Kޓ��56Q=�H�$��ԙ �0�.�<���]��@L�m䵋�� ��U�3��@mZ�UA���{���eM:��w��XK�Nb_-A�F�X[ձ�����aB�G\�#MC�_�іע����t��<b��|*�;!|�|	��!�\����|��؀VI�)"=<�JCN���P>36�������VB0T��ms�fy�ƹ���9{�Za��8S��V�\�W�zh�Oc���ny�	�ɺkqx�	9���
�sv�H[袡���c�	g�2Sd��&e;%zx��ز�^��t?@��S揫8�k��
h{�ڔ� �$t�0��S�1���.��w �@�
�RO�
�c��4BfP Z!+*26�u�P�[� �����S��¡�m�S8�Y����ָ^,�D���ja�sIŦ�u�_�|�hУ|xCgu+�a�Ȥ!(�I�6���� �kcM��q�S��.�_��r�	���+2q�����9�5n��M���|�����.t��4�oW�J���:��N�9֋wQ���=FY9����5�AAqzŗ�E���u�0��,���sYl1x���P�����I֗�v<4���owU@W��B�Y��պ��w��������Rx���.���7�t����7�:~,��p˭~���!~'[�rĺ��6u�� ���%;A���1��~e���뒜j�'[�<�z$���ɩuk~X7�k�$KGggi���{��9=R��4蘟w^���E��<)N�.�ɯ���LΆ'i w3X�Ʃ�����[xx\�:���/�C�PON�S�\R���y=d/���h 5�U����z�(���R�.�����
HHJ9��t�HI����R" "�0CJ)�w�������r�Yf��>�{?�w��
vk8TV�ʩ���t��ftx�����,�[
N�� } #��$|g�Ĭ���r�c)ly��2�أ��6=��pΔL��m�$�GS�ߋU)��i�)��T$r��[�_$c���eΐ�.��i|����[]��1��.R@g���
BɃK�j��������H�>A�;ff7F�N6�y-�7��X������4��3e���<A�l��Ѯ�� �j��f���o�G�0�_�vLW������Q�V@aK�k�T�|�ᶛ)�@.X&���N���ѡݹ� �6�v!�!�I���-�s��ܩ���k���/j����+5�k��n��Zq����;���ds3G�׽9����+���i��2��o�?
����G}گ��se��= M�o�Z��f?n�����r�o�X��;���{�����H;QX��Ύd[��}���d��pm4�3�����1�J���wʔAZ�;����n>߅<g�S��9z���W��](������8���/-����
G0�8�D�.gqH��m��U�ɰJ�P_�5j�w	�||�T����c"@h��'=!�5%ހm���7�\��b~�����X���a�V���2�QD��JǇ&د%�D�t�A��۫��fF�MY�=�j@}�e�NN��*6nF�8��1S�Ő�d�G�#��ˀ�*�T^/��F�d��<�����8 ��q��Z2���+O呕4\�����O�&������ɶ��:��� ������8:2�-�߬����<�r��9!-@J�mRq�\~B��z
S[��Ӻut�{z��V��:��ٯʘ�;٘ݘ��]{�l��d�����}R��7���B�$���R	)k C�2��8��X$��]�!�C_}��?�'6N7�*[����m�e�P���Y��՟]�����k�g�r�(�j�r��_%.��M
·�Z|��$^0ίR���Q��w�ٽc�R�ó s�����&� �͖��v�[jJ���Y��Z�����)-��T@iV�ܣ��~~Y����>r\j���s��̪�c2�e�c��2�p�n/�O�ڗ�U��M�'�Ky�*==]Q�>�	<ds���n׵��*~T	��ME�$�<j�h)-M�����2������EX��C`�S�o�$� �Fv[&<QT���"��K�<ї�	r��`��\$��f�#D��ߥ���HAV?���\�5k�5V�p�:����E���9I����v�
;���3�������p ���j�����VVV>��L(J�juO�)x-��0�^�KaqH�t$+�9n���r�=Eo�Em%F䌅"��ᴷ�UA�&��tq��#]�z�!ul��U�b1 ߿-퀘~�UBSV�)vl��Y^N�c�JI��߄e��˻�{o56������}Ƥ�[l)����rd���q�d��9q���_x��eh0������D[�1�<�]kt�ѿ��/��l����M}о0C�.���F����
ʣn��W�E���9�[#S�R����َC-i��*����&��O���%V��#JK�����ȫ�4��_���_��Ѝؾ�s����:n�~����l�J_�+Ji#��8Q�;k"&���Xx�^w|�� �o��Q��BP�Hr�c�"n~���AWW�&
��	B{8jobq�/w`}0�����dO��T·�����<<�Nl�U���5ߪ�:�;̴�M�����3��]����:��@Zh��Q9�4��d��*-��q�lj��_f��,���Ϭ����4��ci�=Gk"�u��퍾�Lo�������⌎x���3��_�>��Π� )��u������ҏ˲���� ns�ׄ��t1����-��!q��=��BQ��GGJ@d"3����C!de媡��1����~w�?�h&�&E,��G����m����M@��fM s��Ng�s�:%������ڭ�o<��ee��ml �%�� z~�6�p8"V���h@���[瞯���滈�_��r��� �pk,'�S#����\��!��k@��� xc��L��-���6P���RiiҾРl<����B��4�<匋D:�.���wp�0;��l��f��Ⱥ����EtY/��@�М��h���Ғ��������w����o�w�_A:8ˁ
�F�ffpp�����&|��ƍ�:����r�Y@'�k~�_�[�A�VIhE�];
.����us9]�~c o��q�>�)�D�
����y�)�NMz~��\d�͂o��hph*ڣZ� ���	����z�)<�eS�>=���6L\���C�@���B�I��|\j�u>ݾ�Wh��Ӛ�𒎈 Q�$�M/1� ��B2��Ǒ5���Np�|�XX=�V�k��v򆍈�������J8����щ��=qs2w�p����V1�0�]hx�[�(K�Y��ۨ�ZZx�I���P���{�k�Ѧ�R�ԥ�_o����͚��u�%5��]�h${[
3��/��J䲧&�����bh���@���S�3�:ԉT&��FfOD��C~9J�P�~��^|�D��'k�qqZ�ͫ��̓�1'7�e|hp2�&�4���(��v�m�X;���*�pKKٲZ��o�cPű�����\;��Ԋ��>(��݋�����˥�?�5E�/�+-=\-���=r7��8���I�S�d�}n�>�Wv�����1G������:�c������W���>hj�e0!�}6��8ܾWT���w8F`W(&&�4���B^'�����V�����Mfbjj��9゛��@��$��p�c���M
�QǪ�ue�D9Ą|E~ɠ�G��rn/}��g'D�u��X� �L�w����mo���|�y����.�n'J��r����*m���p.7���FȸJp�O���������C�R�um�u-?������~�#�9��{⵩�~���)"[���"B<ى癿?��zn�)Cc�X㷶 }��k��GT�����s�{����ZU���QG�����\T���W���������Yn�y�U;ق<�7[��fB�AOZf �!-���a��_+���m��X�ҫ��9���<1!�C�
¢��@ s+��su��=��'�z�^�C��Y�CW��	���o}�����ӌ���m4T��Ws*.�y�=�p62}X��<�F|�S������hDt�2�!{|m���}����4�b��|}�[n?��)��%������#�h�<��KҀ��ʨ�'O�eɱ��i�G�fEB�z�����:�"��3j�<Wu>[���)��u�G���{���z|�Jx@�}V�_���U@%�ra�k	/1���̠I��G=��8�ԅ6���w(L���`�bY�x��C��#Wl�=֊��]�A(��k�(�L�RM5��u*�_7���Aw�<��	_{��<�}~������c1��,Yv��l��4t�{���"�j��}��nB��@��2)�JE.��n|��Q�l=�4'Ue�pޘ��ࢢ[H��y�ҪkkÝ`$A����m�W�ۻ�'fm2(�͙��P��x��������OS�%��������0.�9�y��2��t�{�q.ք�q���A%[�ڎW� C�$Xp$b��,j*�{랄Ն?ܬx�I6WMF�i��LQ^�śڗ�V�g���߸���*�:�(EȌ��fE�أ�{�3������4���O=�GK�}��X�����q�8௴������^6�Y_�V�	�u �R�2.i@h5
3����7oȇ�=#o@�z7��@����:ܺ~4bk��5�T~�1��)'��|	&^�XWa^�!?u�1�;��|A ����FB&օΘb8���\t�׀E��N��nP��`�rr�$��*��� �8t�z���|���_��ڛ��_�d�=8c�A��~T(��?��wI)
��d���啕�'�k"�����k�qs��ww_IӚ��·oV?�J��_113����Ԓ>5]i1����v
���q��wu��]��w$B�p)��2`K��	�R	7�=p�cy$~�zl5��)��#^��S����j� �L�M�fb�$L��.�	4�|�;���.�XƜ%�p����Aو�L����Z���a�|��B,)�E��]�����q70������\1s�C�Û�z|ፍWpJn�;�X��������.r[=���S��W���kۼ�8g�w�`�jRX�=��/���#*w>�*p�p�`f_6��v�������.]?^B����բzI2�u��ݽK�DME5,��� / م�]�����r�;�e��L\�u�O(��@>��ө0 TV���1E~u�������dlL�Y�GX��-�\6%]`�q��$s`��L�C�B�B���k����a�����)����]�*�7��v���%� ��ϥ3[x��7e4�7���0�l�o�O�Ă9썑N0h�g�+��--x�ӧbhAҵ5����^��������g����,��ݯT
$'����%500��ev����.+�Z��s�A��N��������C�]?:�d4�p�ꜯ��QDv���Ӏ�T��}�C���#�6�(�^b�����o���vf������/��w�s�zIY(�>sG�;�e�q��q��0��׸,i�,��Xd?��'�v�*^�[I~�1l��a�[�j\ɋ����n|���Q����3�H�K�3U�[HL��5����� T�7l����F�]ֿ�{_G���#�*WR�t�` 6�`��H*"�.�<e�B�Y_�
�}
_�����Q�W���k�-E��W0L�w�@�ݱ��@�pP�k����eQ.7(�o��I�f� 1�ߙ�hVE���B�K{�zx����*yј&C�D�m9\����]�iG`��/�N�e^����S��o�oK���m� �+��4��/=��vln��O��^�z��ys��՟?[��d��=<�V�����!�!.<���|j�@>�zC����4���� ެ�N*��	IP���vc��8���cm�,|�\�R�/%2;�%�D��
E��xa�C�gYM�}Ax|�<����y�5��6�%�>3Hew‸�@���&��)	���A�;Hw�1{X��0�36q%�.�_MB�Ç��@'+~��8- �&@�>�v�UFD��I��6J�%��U5 �J�6�/_�
k &H�-����>����d�O���c�����1���. �CHx_�#��>F��11���ޤT���!145�&ڷ"�����Ąb��bw\�n�����ov0��׷���K�o�[(^��9b`jJ�8<Ħ�7��|:�w�����A��T744L:"��m��&@l6|��ر>�q�Y�H돫���f�JN���F�=��,��G4����x�m��eX�{�qY@|3��o{!_;�g��ϟ[�H��a��� K�ګ%�����rFĲE���}��\,%--_m��2'b�;�~y��'"�'�Nk��^m���22�[����\���(�3o�?�!�ӧO?�I� ��GL4��E@���j��[c�*א��L�|.k� �h��ꬻ����.��O�?�B��,�!�@�NOZ������� �Љ��dk�r8(J����Z���)�rx~{nu�W���B3ZY�!���e?������m ����(;��_��ۼ$����[��������;��8ɫ��"22o�'����G�e��'''�"'0{�<!��_�|IZ����y	S�u��f�����}���.��K]J�)���Jה��J����U1G�٣`�C|"�P�v�<!��o6��{�=�֨�O7fr��5.Q����]ܼ�LN�f��M���r7}e�����Z2&!�^oMY,��A�������6R�[i��B9զ���o��v�i.�ŞtܾlG�*B�2�f���l�?��W#�%�Qj�oi;i�`WU���Y�W�~dk����o̞K�Oe�}5�G-8�����o���̪��U#��W�"���-���"���f��ζ��}(��'(��L2x��8����@��CE�]ŷ�6~;(Ւ*Y���6A�����
���X��e'Zγ_V7L�_B��fW��o*�	�I��u%ف��ٶ��bBB�����1�~)$R$o�fV����%�Y�k���3Su�=��%��T\�rL�����M��.r�R/�'�./_b�@���ӏ�ŵ5���h":::�\9@����%���e�3�-|OĚL+�?�tR����bFōD2�k��J�Ԥ &���_iz�D� �"�<����{{��������b��{���F�&��0����VX�A�XV���8|�4�>�� �rҮON>;G~v�v��P�$Ƴ��8��d�(G_?q����~�J�Z%�n����:̡�4�/*WFӹ�����4��-K�}�?�R�w��V�`{���Tb�׶3ƌ��|",fvw�!�e��
�뻍�4���v�z�j1 �[dr2��$�7OY�q���������ڂ�&^626�y&��1�^����H��1�j��>cv^^p ,*|ိ[���Zi+i����'�[(���m��P���}u���⥦=�qq!y<GT����U9av� �DE����=����^+��2S����&6��^���k��?�����C=�Zޡ%Ξ��Ŧ�h:K�p�Q ���O�ޘoQ��41�O���N����1��
@B�8�=��U�굯���3�yP{��Fөb7T��фne��,zy	[�x_�V����,���Cž�����ag��4��
���E������\}����f����AlQ�S@��B�����=��%`@I�3GC+�Dɚ* T5��a��4�D�� H�%E�V�����%eX'�.؍~2�PiC��՝�zU������'�y������8���b�ru�`z�~N��uP��u���Ο��7U���PV���H�5 n������k��JF�4��iI�z����Du�-�������{�ӽ��kNU����g�Ƭ95��c�ۊxO�Ͻ��ُ4ܧ�%�L��˔�'#@1r~MzXc��h/����&��ft��l0�/2��ur{���66�P�I�h�q!����������w4I�LE�rrb�K+���C��/{^�l��ܳ���7x�+;/�`�~1��9G��;��L��p0������]///���F�+G0�92��n�L��C�'j�K���r��l��rx,ɠ�ig'.���V���ur+��f-����� �߱��^RAe�}��D�E�2mg�?FBt�İ?`��G�f��Ȝ�+��	ܻ�AQz3b��tb�Zة�-�)�����^a@��I����D�`�c�$f��#�.��\w�z{[�',n������ň���L�倿��'k@�F�epF��L��?|l�����J�D/A�X
,�S|(%.A^I�
Ǘ=YX���I
�E�@2��牯�]@luƚ`}�&^��q����-R@m����DDuw�"�Å�*؀�VTV>m�����5�1H�g|ʑ(Z����Tm(W1��O��@���7�t�\[#�2\*j�|�X�T�� 6�%c2�4�=�d�Iخ )��q&�@ 9Ȃ�%����/p|_�8����k;�v���4Z����j8���}��晙���j�[p�#��[���F������A]-���ל� L�ܦP��f�1��j���8ς^�o���T0f=�*�'��wTo���G�(.C6o��m���a|W4�	ɀm���"�/Q2�J��041	�"�\�΢ݱ�c��L�����v�фHe���s���J���r��T��A+�v�٥1�mG��*��P�C��nE����gS�MLL��+]x�����:coR�7�p�����BJ��r�Iti�yX��(�z�֦�4_w#�7�B��6o���'V�����/��q5i��$G)�����8X�X��"��]�o��E��R�+��苡�1gg�Y��� .��B��������W�yP��N���ǜ,1bp�����n��+$Ȅ�j��^�b_��A�Ȩ�K1�
�,W���]���_�?��ȥ���TxiCP�3	5s���jo�N4a`����tR�j������n�o��r�ջG�����WX����ZoD��� G?1�<`�:!fs`˅��}46�t�wt�	�2�����U�J0-{6���9��f�(3��k<����,O�������#���ͱ�5�N�=y�˾b{�w�9�͎�ȝ�=U�C�հ#]$�����Lv����C����1��!.�gT�*�9��t���cJ2�o:(1'ggׁS��o� "zX�e"���w;��&�JJ���Xz��EDj�W���N4Fn�s�#m��P�c�W�4P�Q�V�ܽBbbq�۴_f��W�ڄ���I#M���;C/y�]��3?��8y}}Z���{���l��8�b6�UR,��f��s�s�/7Y��a�$z�����<%%�s1n��_1�l�!��iii3��'H8�*6n���@��a��G8�_�� |�q�lj�+1�����eUlDg%�C<��Z:U���\)e�fgg�{4���|�'��Ϗ�8�8����9�
=����� ��.��c�,\���;O���9|{	�ڃ�~���� g��}Wƨ�� Ui����ss;''��^��|F���P(�+K��@I@;����m�)x俓3��}#Rk*�FՆ��f
LB9ܧ�ু�;�!nf1�}���:�_�;��G�3��uQMNZN���#���"iʭ���B2�	q�8\����+X;��\�H��[�'.�a]gQ�Iaeݸ��@��g5|��1@3���6��c�	��oqc��W���Z0�?H����^���gFL_l Z�U��	�?e�L����t��{��FB ��d?*�\�+�g&M����}����Ȩ�Q~�2I������������9���O��=I&&&�7Tc؈���P0���]y_�~q��t�c 3>-�L;��~�:\/q(DÁ�}�\���+�'Xn"����ݕҥ�/]� W���b�����{�z��*O+r�/:6)H'M��KB��h�\�u{H[M&OA���t�^�0^0��\���qo�ZEpݗ(�Q0R��緕�ݵ�3{|��XO�lDHF.ԍ-+���1��tx�;m�e�D����̽lg��<��B�C�周f���������罰�/Xۤ.���%�' ����;���8�3�Z��2̺eh:4�<���~���	� �`�Ŭ�/ވ��32RO�,"�S{{�Y<2r�>��Z�v ��Y�`���|R��h���~��KM����b�^���y���[�Iн�*��#��Ԛ�܈�+�/@����|����K+%��$tigN�/�sM�N���Ƿ�i�����l��PRr�9�=��)��˾z��eO̡t��ݽ�$Sw�ލ�Y�15�	u�� �77?pr��>�&���W��)_�C��y[U����@	%��h��+y�t͙���5#c�Ml�a�ׄ?�7tMB���E�L�+
�a�ڏs�}7qS���.//�c
N�ʔl������'n���z}�ݠx�%Wd:' ~ȶ��N��ɗ���	Ω?,����&�eБ5,lJ���ۿ��s������T����Ib�u����>��T+~�t��n�Ie��xK,�]y|�OSp��Hb-�M��,����!�͚g�9.T�Ƌ �D��*�J���-f=W�ua�'�oq�ѩ�H���"�+m����*�.�� ��{ו���N�$$%�>��)�X�|����o�ha�_�+�ƽŭ��j`Z��H$*NWK	**��;�c}gOq������/��l%�� ����V��NS3�g���v�\||2�6�a�C�E�~>��d�lAOn�z1G�,]Z������3_�xm�A����Gf�3�K�6�2�f�?D��tRWrIG'�x̉��Q�B��e��?8��0� �a���F�g<�R<[�� ������W��@��HQ�����HI!#J��7�Y���f�2�[�b����AE|��$����JET�ah�W	�ZZ��K���B�Q)�w>�w�p�z^�[c�e54Š���k�δ��*�U�Y�׻M���P�®:m�_���`�ퟲ?H
	E����FR�����Za��x?��)��nT�b�sW_zf�";u֮�������C�s\����t{��(����'AR,�h���_��\�&(\�'��6�X�pÍXF�\�ѣB�W���9:��J=)h�� A:�Y7#�<�4S<�C��q�	��~�ɴۘ���]K�țGT�����
{�� df�~k<�4��uӰz
��^�`���̳���YcG'^�*��N�OK��V��W�;�=�ܺ�=��]��F�����~�AY8v�L�eu�V�t��b�X?������T��j"�텴��$�#� V�KG��W�nk��Od�;`��m9\�n]4�>��E��)���+��Ȅ�E_>��֦���`�R+�ҥ��K���55H���Ygkhj�v�,��`���~��w(�2ɫ�E_���v���G�]�s D�&ܶ�o;���:�N�L4�������������W��$$$[G~��5P�l�鵋/5��21X��(x�E�R=.� �{y�lR<{��F��qf����K��������Y9	���_���pN��61���d}QN�%8���KI\�XU��P�_�������&y6K��z�M�)s*0�x��3Ym��7n|n,��N��;J�$����$.�V [:�����7H�}�U���m��U�"!<4��K-��Ʈ��@{���|��d�⏒R� l�r�Y|�K�r�+~t�o���@��;{@ɼ�O9�����e��Pҝ98`U|W��}Ax��
]�<��z`���Jcm$��t~Y�+-��"�P������������MQ���{,�y��G�����zO�Y�� ;��2 �X���%٘J��Q���`C'�__�uX��++W��wh��W=L{��q��&$S���<���V��I���oQ����C1�W���!��B�8&�7Z�X�dX�Ym1�gm��nք�� ?�+PR�x�:|��3YR�?v��C�]cF��`���-
/)OꉋdNz͟��jԣ(�u��;f��r �9@����ń��_iyU��J�饫k������!9@@,���X���n������vihk�͍�<����ʥ��u:�W �B���A�v�| p�±��E3����������7�U" �}a�� ѫ�����䃓�����+������a��0�%{=%ʛ7��`�/�5T����j���������8v�ŀ���"�M�"��KZ�<��g����Â�>��B�v��	}~�l�\kYѶ�B��}n����?���=޲:�a>��R0�ϟ���Um=��M+��Y�����2�eq���ەy�����ʼ=��Pah��¶��V����}�k��]C�n��8����s{�푝Q8"Q�y�ƾ�g��
['������e�����:���6���mV�苛A$r��:������%��~UD�VL����7��2�˃���|�(~�宀@��a�r�N������Ώ��j�G5����SFG�����|�C��䡀��d����R^Yi���7�y;E�ϸO�m�A��l��V��ss��cRV.�Ý�@���v�����dg�t��\O6!@�A�@M�1�0��_4�b�I���w;�Đ~?��|����)=c���5�^ˇ	�d�����de��釣0�˾R, c�å��q���|��er%�� ��[���5��@9�h���0�E,���B��D`ܾm؎��3J��/���(��ؠL�.v�<�V[~�$���l7�ᗗ7��T��¤���»��λ>��6NK�!!=K�Up2�s�=�J�C2缓@��2%E�C���K���tY��=��ϊl�gGFn	ܻ礮J�Dh�66���\��o|,�L`|Ni���M�3;�--��,����n�� e�d*��,7��Ȟ���w޿� ��4u�����\����x�5��#T !+� �U/
�#H"�����"��S����_.�D^=}%�����i�K����o1���n�,�͗��D 9�ܻ�q�l�:q�OF֧��t$Fs��G��R,�of\$��Sū����c��vKq�i*tb=�y�,
|�L��qXz�EwOD������ݖ�����14M��zv�'	��*G�/�k3�/��˓_�lV�hV��द��n|�ՃV����`��=�BB�Əy�n���Btw��9�E�l�������;����ik��?j$����iȒ�Y;�4��2M�}89qvqu��k���;�mii�GB����$�ܿ�0��[��0`���������]3�_:B̨j�܄X�c�w$UY)��e^h\Q��W�U�V#�^���1|b���B�1����z��8��A��L䘧>�a��qWy(dݚ*�6-,چ�f��/FJ'Uw��#�W�Q�0^��ѭ08l�f7+fW�r����9�g���V)�90�]���g�߈Y�&B�v�{�=�_�=���@iARN��v��d�C�/%�3��!�3�3���3��ȯu��=ր�b��9O_AYY�ڬ+ckd�UU�${���d��NW�x{��|F��CB�*V8~�mI�g���ҠJ���ߊ�c�uDȢۨ�x���?��G	�B���ܟ>}
[Y�I�'�o_Ѯ�=,��ԜxƇ�A`��*�Y�oVU��;s|L|��oJ�&�J�n���[�� %{z�r%�_��4#�����H#��>%��!����"6(��N�~�g#�R����sں'Wg|�7/�j3�	��"��Ӝ�6'�i~�k����Q5�h<��Ƶ���(_�;�R�S�=��n�7-��C�&%�"(G��z:/���`6�!bsp����vCN"K�WIIv��{���T+^P�-��z_��%�ͬ��I\�!wrr2�ћ�����������;�Vܷ�����4��,\]�gV�Rԯ<}:��CM���=�xv%�sV�~Z�����&!��R�Y�D!�g�!ߐ��'i��-^lD_t�n�% Ǘr,1֊��}�Z���29xb]����"�}�h�'���0���^�DR�g���.�$`�|�5
�/C��ҹ\jP�#-1��sƓ������	�C	.�̞��0{X=+��I�w�@V��T�Kr(�ݒV��[u%dEo��j���<*ݡVxT�r�+�\�f�yՀC�^YՌ��z����uq��lZV�� ?�8���}3�?�GnLP�Lk��$b�{ٿ\Z��"U�,�	~��T3��02>�dS[[��X[������
X^�@m �h�s��D]�+���ѥn�u3A�
3_�i*��ttwEF�{�X�=��[��������=@��҇�ݾghMO�"nʸ��C������Wk��B��	Jx���������ʗB�u�K4akDXV�k;o�-���r�@��� ��_V�p�C}���+�4
��hۧx
肍2�a����wb�������o5N�)��{P�s}[<c�խ�81i`�Y.�i��>Vb�W�.���ey.��c��l;ٯ�f�{o[�t�4ɔNm���k������Q �3W�b���+���0UY������'��rSӁ���4�Xʚ���R����FFJ%<�L�D�/�d`�g]b
&O�KF8�>A7� �4��j\��������A����i�XV����ˬ 7q8;^��U��<�]�#Q���]�@I�*��_n�K5@!96����y�	&�Wl�t�Z<-f�]׾�r;U��:.����t��J�*�m��w�uω]�(6"J��QjU%�qo${
�Ԅ�ˍ���?z�J�-X�<8Рk$-t&\��on;B��.k�(����bV6�B���}ڬ�:WW3W�>�UE�;{6Oڂ���/�Q��N���n����;z��k>�0<<�:�h%պ;����pGFCI.("��}���IIX�9���}q.M��<�Ŋ�#b��.����?����J��ޤ[�*Z1Q]�c�M)Zg,ū���J2J���i��G;��mJ"i�#?�j��t��Y���9������)��s\/�n}=�8��ס*'��u�0F�z������0t�ڶ���G�c��ԗ��4�My��Z0a��$�b�xl��ݿ�a�sz-��K3pS�q��0�y���VwOr�c@��b ޠڎ[>S��C�ʎS����nS�323?KE��{V��0�S|:�`8�Խ��OmGo"p&��;�C����16y�L����&�A�'�[�r�I_��l`����5;�+�!
C�6�^�=���--rᕌ.��Qsg� �̪nD+��YS'q�8T�q��q8�89���.���|�n�Rm('���/��\E��hM'u���7���Pj� %[��6e� iWP%��)�� ��ZE��V�5�?,7��U/r��+(�/�+V�ӽ��`a%�$�i��A�\�S��m/��^;h�.(�ԁ����`A���++N���j���΂[�:k�v4�*�������7+�����N�ґR��R�kk$�M �rr^��H?&*{Eܙ�hP�}v�@4+���pI��૥Џ�� �g�x���G�$����rk�,0�ʟ�Kp�Nj|ߣ��yݷ�')\׀�/�<AR�[�@3{o (�PK�M+o�:�P��@Tl<EL(UtA�������ط岏>;r�@��p[����O+�a�M̝��:�v���2�A���EL��b����t�$�k�&?�l�a���Ɂ����g�'�ퟞݿ�
_oS�q�I���V�K6�J�������ihb�9[�t]R���?��3m��'��ܦ��� 	�H(�ʬ�<����N4bo�L�)T�����s!j��KZ�Ǐ�����U�,�uZ'���#& �r�~������A ����zx�3����jb� 0�WK+�g��I$�E��[׊c�@Nלﻌ�c��k�����h o._�g�e7��Ł[Yp����ae����C A��MhI��C�.|"�!���y\j�e?�N�qt�e^m��0�<E�;��������v���.��!�.z9���^��UnS2��U++ī��̀~n�ߚ���؎1�vVK�K;VSu��v3��Ŋ������SF����
)��Z\]j�]S���olr�G=���~ʰsM�i/���P��%z�Κ�L��[R��sD� �ӵ���'&��3y6�߻�V���Z��ߜUmH��MM3o�֑=�6;-�<�C�Aӥ��B~B�=Q�C��Pyդ0�j��֢�#W :A7R?��i����$]Y��Qv�h��Ika{3�OF��rL��'������k2&Kk�)�C�|�޿�32R�1*W@׽c!ë&W��6��W���Û�V���.��B���N�t���c� ���ǂ�穚͛S9�f�\���w���.��|�?�=����<���qu�<姶sj�*T���2Α�T���4�v!./_b�xA�����{KIX��h��D�Y���J	�H��o��b�],Ñ444� *�wi�>pK�^q�cT�O��v�X��A��@��N�hc�}<�vY���ݘx= ��Y��{ ����.���]a��F)���1	�0N�S� D��@�➗v㤡��B�׋�q��Ƶ���x�7m�Y�E�%���&�&���4A����k\ޤ��ש�m�p��Z�u�Zq��oR?�cOp0���>����`zӆ�����/nU�B3A~r�5�i�a㮸V߾�>�Sɝ$s�g��4!}�)��fT1���~�5��; J����Y�M�@l�v���7UG��+a���c�7-���===��9��K;~~�u:��s壗�22��Q� ��_��5�+.�堦�''h~���������f�2L���r ���d�'����>�9���Y<{z�DHx�g|��ѫ7J�z��GG6վ�.�39	�_�`V..�]]][�-v���?
��W���m:>����X��e�N��{0/--E)[�
���l4��0���[���+J:*�����%��@Z�<C3j��H{��=u@�Q��U��+�ŝ��Q/,�<z��m8f-5�����6�RX���=%���o�A��R�n�{{���Đ����6���k��{��~�3I$"��כ*Ƒ�MĐ��#�g��F����A��u�razz���;t����V�Zy�� ���\M�U�|O�$�`x���}a��o22n����Z��~H(�|��&�g/_��^�M�:�h5S�e)�(V�v[6n�*����H��<T������Y&��5��31���k��;S/��Öxl�5p�_ǌ27���(n��J�9S�������%��^�ȽzuR��Ow+��4t�6�Yo�Yqg���"��C{Efzƴw�d��qCU!Ƈ�#���O����D�e�idf�cN%)�Lw�e�է@K��x��O�����<�a�����^�GtmR�>�z^{���4Q8&23憆a#�+H�� �{=������5�7k�[&�<ʳ���pw�M���Qp�v_�l�b�β��i�����Ѓ�\xY���@A�W
^h"��2z��{PTS��DY�?���vݓѳY���Q�m-XV�D�'4�_���������Gf��Hߕm�Ev˱m=N|pq����J���9 ��~������T]9*9����`!s�6]����{��+�]�ٻ�k�t*��Fp�s+(t�jd�h�A�Վ)J05�+�S�9}A]�պv쳾�)�NV�ƃ���3��GȺ7)P�[/��w���q4]�lf� ���K�D�Lc�{��O��UçOm�qqq���$(@8NN�o����}q�~ci�)"%e�����<C~:~�f� ��z[+H��L$����B2���/�N���?���3Ԍ�zzAW��q�,"?��:r¯NO�"�q�v�r�Ɯzff�""#gݛt�F����J�~���Ҍ6�L�[#��Q���.�6	==}GGG�Kr%��K+ ��[u����f�rz�Ҕj��ݔ���M�]Y�����|�yV�XI�B���n��u��u�ؔ��
�>�?���v5Rt=PHJ.��]�,L�9��_��\�+]W�&�O�{�]�����32��I��4Y��/����Ĩ윜���N�^m�/q1ۻ����ѧ�Jf���xSt���y����ۮ��{M>��3ss@��9l?x]9��͍X;O&�iv���v��h:�x*����B��!���#�Yɱ���cdfo�압d{&!�ӡc�8f��]����?y��u�������k���m�Jԧ)����"��yw�<�{�8��k����w�ֲFuR���DH�1T��������R�lT���N����C��f��X�ʾ�j5�,k���2�@�H�M�W�ډ�-d�z��Ӣ�y�g�|��]8��Iĵ;��P�Sa��sqi�Jk�a��]�W��u��JZҋt�9՜�����@VX�$�"�e��E""�&m����h�[�##���34�Ty��	4�y`}M4\H�uE����n��!D�m߾񇇇�㆗�nl0��i6؏P~Q�fl��I�+��,�ֶ�ʦ��#**�{,�=�Z'��ח���W����o������IIt��鮸ջ��θq�Dqё�M�s�����*߻)3Ʊ峩p+~:��	u�����i����ӫB�Sc^�.v�o��B�����t�N%�RYt���+�q��V%=ŠKoP�θ!��<)9S4�=�����	f��.Q�7����;Da\k��<F��9m���k[;�Sn�pYG`p��Ke��,%V�d9�R��z�<����afe�z9=�t$����:�LŮ��(�(b��Q�BaΠh~�26-��n� D3F�oA��hu��F�-���G���?UTl)>��2�@���6p9�Q#f��]�f���_����J\Gj�A������:��ƥ���
��n���xE��Ot����I��h��Z��@����ß
m����*3�'���K��p&u�yh��Y�vfvvB}���%3��8���f�̄X8�>?�^��e/�B�h	T�"�V�p�����dy�������ȗ�Vh�%�m�8��4�2�}�[ƽ��o_U��<��0�Հ�
����+(�a�O#��a�H@O�үyN�&d��u���l>�\'�@��\S5Ӵ�X�fSh�0�sM���2��ۣȾ��������O��^B��㝔i`�������@����Дd�ۢHeKK���M:��_:p����B�f�i�^�����]^P��/)2_:Z8e�7X�GEF�y�p�]$E��R���b1E˔�����宮0ꪢ����Ծ��q�v�]6�©�E�S����_嫪���nlZ�Ԗ��p%Fn~ 0s-�N�?'�ᄜ�Ǵ�!�D��jо�����.|�Lj|mo
���TM�6��k��`l�K�T�M<����̫[Zz��	�#��Xht7��e����.������h���+�&<�ƻ,��0�QvAA��w������v�a=�e��C"��W3M���H��j�{�,[[���"c��wɑ��& �!��Sh��$-7n����ù�1���?B�Fk�C���AoRp����^9�dB3�MOrt��̘��������}�|�٭�͍����Y�/|^�u�.��m�>ZT����QP(���uJ�2�K�HRSD��H�s8���q�@=[��v����!��!��v�*����!�%������V���*�luo �-��*�{�b��GoC���keP�	*	�!~l�1��������k�T��_ut�薹)f�,5L{{yED5��R����%I��dL�G䨓۪���2cC͐-���b�/�М��L=�A�o����}����`��z�TQ�nұ����m��TxhR�DP_b�ld��yH�f�)tp��>���E#ߍ��ǌ�pӥ孺D����	���}�c٪�5i������5�K.�rbi���S.�(	��)��ʏ��i���3j_dӵtg����A�+���5+/g��XR����9�Eu�v�H��`� �&�"eÜ���2ܟ"		y���C�UL�<h|��.��5�ς�p�8��%��Eb��]]���yGvk�������W65E��Z��@C��x�uXՌ絘��J��Ķ�k:H�����WJp���d���o
�N)��wG�A�:0Ӕ�q	�k�<oE�8�PS�n�Ȃ� =��^�c:a5F�o�����IRdZ{Kg�!���l�ۋ�w�*��T�<b}u��@�cx�ו������e`,�h"i�	a`�;(��J�:���jE��$����n�<�n(..�QgN�^��_�qKU_TNNď�ؑ����XJGw�D�=��s�	k��q)�������n���F��9>(Ywq�����KK�����v�=���O,w��ma���&($��Pཐ*��t�D�ľ+�8V�oZ���n�ݓ^]��y��q�8B��C���ʶ�ë1�J���@��W�w{�(��|�^�+si��C1����q����\�ӥл�Vj\
��-l�׾>���̸���5�%�G��?��h�Ԏ���5O��4o�(��:	�N2�\N{�A��G�-v��.�ywy��P *I�����L�����+M�U��my������������:Vu��K����D�#�iO��R$�g|�$Pi'��M��63<<#��Ɠ�0	�<~^��?E8Y�<w��2�~t�bP̃:�j��o��>]�@/����~��S�N��P���J�k�)xv���z�>?��.�\c��O��"�����gΠ���
�#��P�N�������&�4�ʉ�B�?���93��a�]�%�u
ݦ�-���χF��ǵ�c��qо�+�Zwň������Ԑa4��O�@lԍ���Q*����y4��_x��Э�;=���׾Z���A!*)���}*@ղ�\L������b�(ik�/����7=mű�S��T@HDTU��X:0�Dx}����9��l���^��J�>����� )�L�+Ƿ�:wr�����Ӄݵ�،��&ip�M�Y�$%��z�1)ƥ ǵ��������3�������;��շ=�Z�w��oy�=HS�V�ֻ�d!%��0���c%��\�R��7X����b�͞.i���)td�P�n_�����@���N�9�C%L��6aj�3P��
q�9��T�����
y��~���>�+��<>Й���p���ϘO�Q�XZwvb��ʝM>T+�fP�߿o�D䙧!Cڠ~��=-��n�y�r�O��.2�� C�*�ƜN7Goo��ǅ=�#�ӣ�����I����k2U�b_eJEF�t�����3SVM8u��;hX�I>�]|�=!B��A.�%-#!a|QRr����_�
"`.!��zt����Ǻf���?�1�y�(�9��^�(>����N�f�d�K�+)���-����ND��:0�
|,wo]��g�~r[���,� �}��h8�p�Jf��Q�-���+WWe�ˠ�A�vL�զ��,�J�u��� ��}�wո���*w���?>��=h����5!�By%H���{�%3��������OdZ"��D G�-BH�-�i[cFM��V��hȡ�;8 �'wF?'ٽ�,h_t�D�,IV=#���;�^H�B�����zs�b�I�3Ow� dE��3��kj)v��0�Z#8�P<Է@�X�XIPq$��R��Ή�8�sR�}�k�c*�6�����ts�"��+�'CyZ�t�t��(X��E���{��ɠ�U턜����ǵs1j��]����nn�S_	�G�g񀘥m�=#--lp��|��Y�n��(�6�=�-�,��xH�ع���T;ji+�u���� -\\��	������TH9:�	[�D &  ���N(h�?�42�{B|9�.JJ�_f3D�4;c)9W���wr�e�y�Z�Y���|򭎯���U#@Xٞ�w�a��z�)��2��V9�F�CfC�#1�����Z�G���g#mH44�����/����g��~ީ���f��������|Fژ������\��"p:�[������K��N{�`��f��@���}���|�[���I��/N&�P;|k�r���,�\��9�b��	���b�7W��;������Ā��w>�j�!? �.�gܨ��G>�b4��㡆��e�s�WRh�|�zն?�MZp�R$a�_��6U��{#kG>�ZvH$Yt�X��p���0A���/#5>��s��<��C�x����}8���p�������Ǹ�r�UH�RL�`��`�@N��3�����^Q
mJ���k*����g�[�Hķ�A@��ܑ��.z��|	��<{.�055��	���{\U�q�n?sb��Y�p��t�0>|��<�� ��dG���S�Y��
1��T�֛�6���jrh�۲��4ҧT�9w�'����;�*Dޢ������L�$��ȸ�$�kp��S!ޓ��5f��x�cr-u%~:����@�@�Ix�@M�\�u�2ի@�o�z��ғQRާ�uK�����Yg./�e+��%M˸�Cw䋮����)4��ʛ��S�l��gTԽ��١�ˀ��/��DLWpZ������ϘؠbX!а�� 4���C	�̞���`T����^Z���qq��L���ꠅ������?�Ro�Z��$z<g���I�9Z�G���4:\�b�
t)Q����"�3��=�������̖w�I��X��> �K�|��E8~���?F	������yJdh;��
_�������^�����fN��O#��{ ��������W_:����n���E��x�>���ˠ�{��MV��I+^-�J��m�6Z��<M��ށ�k�|�2��"����N��ڰ:�#l:�<Iz9x�[VI_x����u�7�o�bt,ʥ�ߠP7}���JJ�:�1HNFv2Z߄��K��������)�%%�15�y^6��^0ۗ�r�W{~��u�O�ࣖͰ�C�F@@>� U���l�gd̅M(Zk'NA8x�,���+�Ag+���RR�5R8�&�Fȓ�LFQ����i �Ϋ,rd�O'�?4wݗ��휡wʎ�����o��g<�G���I�Aֶ�AV�ʉ�@Ĉ��B�d����M��>�:����k3��I6Y��H-o�9�=Ar8��[[<)��8p�������x{�֗���&_���TR����D\A��ý�ۀ߻�x;��w�:���_Y�"Ѐ��)죦�(͢"���&���dH��
�4'Y�Fn4�'%=&���L�w�SU���zxuk��RU��A��7�_�(�1D�0%G�%V��4���
�:/�&R�`�7T�|Ñ/ܙ�l�����Z"��=�H�P�C����PS���ʅ̂�@l�u�l'�F�?����Ύ��;WMm�~����7�V䑙(�������f�,ll���A�
�M��KemoO�S�����3F���e�E��7��2���g��k�c�SH*b���k�dq�p�AS�C�DC��A���|_�6E ږ�{khh�$KJfA������嫠�=:�딀���������P�J>#4��2��v?��RzҤ�$Ǭ��%���!��R��A����a�1�q)���#����*#�B~�1�O%Y�/���}W���z>���Qndf��lBl�=�c�0aɌ~�3ʋd�+��Vp	|�d��1�E��EQ�#����ݑ̐�������g���`�"�d\������{.,�(�Ʀ���!�΄�9��'�@�����f)}�;M|!�ijn���ε�y�bi)İ�5G�wvB��YOt5*�լ,�������2�cE*�yt)��D�_���;�� [�����r܉<z����-H/4C������=�ݨ�r�ڹ��%O$��;фߘ�j�Q6��:p�|�(mB��tyX�[Ф���_�@x���X��_U��vw�`R�m�����0_�4�5i(�£�����?��`�j��ꭙޤ{��,ͧ��˹Is!j���m�|8��n3�Iw��}ĺھ<���O��śĬ�Ak�x#��ۮ�e�9p���v�+:S�\� ��f)Z=~�\3>���/����WKK�����鞒1�3�y�s);�G�uu�S��k(�b��W �ݾ��r*gPl����en[e*�x��>�T����uM��HuUCK,S���;8s��x�wq�!;p�u�%,�"�@��/�ފ������� 6^�dMB#힘&Ĳ7���}�������NJ���P�!�?�}�t3�w�y��Ś�?�fe-�~�al�j;d��v/f�	��i���2�C�P�����kFFС������p������g��0�(�|�@tpb���f�3��n����(��(P��E�D<ˮ�P�9�{G��`��w�''a�koݴ�? '��G"wTe�u$�߸
�ii���G�y<3o�%�K���HNLIq^(w�r;��I��#�d~�
��׻�LӲﴙu�N������K����7O��4�)��}T��� �Ȕy��
��-j�A���!bCF7��no�nz�ה�`�X^Ǯ�Ft��\�Q�Z�?V���Gll�ۓA�EH����X(i&%���WcV����b����;�8Bŀ��F� ���hfU�m��/6�li�C0&�QG�Ë���(()Ü�Tg�]&�`!�� ��$ ��J�(���,L��n�2IN %�O�rp�M�F��@=6�.�=ͳ�[\��x����d�\n.*��(:g�_�!�M[,Mh���$�>�?���0�D����L:S�������@�a���-b<.~=�pff����1qzA�>~��Θ����c)�	+,v���t����~ĸ�q�SS�C��/(�eQ�Aw��	��Բ�g�y|�Y�d��=��[8��u}���97��>k1WPXh]喾���M>%o�J���㒕�M�Ѱ��C*����	�+1�y��H}��kd��o+�"�"6�җ�m�&�|Gp�mk�2k?x���y��������j����:�&MM�zHr!4
�©�e�>fP<��>7���k�;��iďZ�-(|BE������O��A�.���es{���a��_�U_�FSrLnYߠb/1.5�8���6����v�?Њ���aVt'g���
�.��Uo�z��Xw�Iev�RU�����}B3B�����a�be�* k�i�§=�
��v���B�����5UvD�I��.@��u�Ɯ�_���W���w4E���US]v��+t����ܿ�}��A�mȰ�En��Puu���I|�������A����w������GC�H,����rPKqD�0f��bb�芖TϢ#�Y-�\ǔ����o�B�����k��ލ��O���_&�B9j|�+rm�#ǋ�B�M�feл�|(����6�כ��>�Xp���P���\\s��U���)�n����3@6��A	�.�Rj$��6�EI����Z�rn�|a�����A#RN`$n�N��5t�l�m���7X�TE�ƺo�zV����C��&N�h^�Frh�*����樽�G��32X��O"����o������iۉ���r�;�<��J�h!:��u,�MLxI�����wd�����[cu�^��W8��z)Y����Er��=�T.�et@Gm?tG�!�\8fd��rÓ�kHj�-_Q(�G`{�a���7��  ��}�'<��Pp�O��S���^���4�N��� ��5.�����\\o*��Z��������e:�����W�R�����Ç�;�z�w㔄-~�����i���~v;��ú����C�ml�S��F��2q�f�b����HScy���z��]���Ϊ��r��jnO�P�|�YD9�$!$�>>.�םb�C�V}�Z����"��+"%Ek+�B,q��^�^^�qj��n��G��bT����Մ#�C�����G`��s��(od�C&Q#��~��~��� T�k��jb�&H��:��#"�kv5x8���J3ā��fmӔ�J��ZJ�T��~	)G��b�w������������o֣߮�z�w7�e+�~���8�5`�|��\��
����j�h�0��B]�����}z�w�L hZ91�yLI�C����c��b��g����[�u5�[�������<Y��� ד�1�
��LDD4l�<x���}�4`c�l����-N>�����I���'�踴��-s<},��?��r�L~�X��]�]�U�T�8�v�;o�J�*�Ƭ��x����l��e���=�������.7��"�ւZ��j�i�[" .c}��-<f��[&ER�W�H4]W(�.���:�r�����3XT-4�tlE�.�M	��n��ncن�5O��޺իF� ��iZ�Ĺ������ݿ�Ƀ�(��͝�ۿ��#>$|1�^nF]*�k`�ƋXR���y��b�j̔���[�z�|��Q�Yx��;-^P����݇�'�^�Q�����]pR�?��߷n��i��W�������=�r����ǜ���A�{$��Y�6�p�-'U)�\����|��Nt�b2���[���Z[K������
�¢�}i�wJ�W�t��N�a�� ��H�d�Ι����ˋM�L��]8�T��֞��w�V���_κ`Fƻi�)�Z��+C̕��ۀ0��d��!��-.~�p�Q/�gmv�nG��V�IB���&�,��HYA:�uٻ��O���?��ʏ�md��\&H�ƜN)���6j��u���mo�0,���E">ߣ�"-��AG�1�F�fcnF��K������z� u�4-^-�AR��Cy�N��^o [11�q���b?�S=4�<`��e�����_�3t�:W*wn�'���g�R˰ B�Ѣ�/�%?	����B����7�}tG]\�>;<�_�|������:5�y�H_;�. ���"eGX!x6���ȕ*"�u%�	����@Ha\��8��]:3U@w�G��o�z�|+���9֥"�u$	�]~�ʝ�V��w�!�67#7}J�:1�A�L��"W_
��=ٔ�7�{�\�9�'`?��!4���z��t��?_Ҷ���iQqP	@�ٙ�C	�=�fzI��.��B��<�L��[��R���T`�w���(���xRcVU��f\z�z���T�����n��\?]c�S+�sH)�ܰ����Tb�)W_��g����q.A��W.��0.�]qI�E�b懲�u(F��ȗ�CM7��wPr}u����e��G V�)5�}8�����!U ��LLL R�f?q~���=s]?V"��,q��QE�$�O�ax�K�=<҈Jau�� `��p��טG�G�v��z�;Y'k�?C
HjŎl�D�IE3nŋg�6;����=��SH3h-�A�Mդ��%BSU>Ħj�?�0i(���#٫���z�%L����3^
zƿx�IU�I����1�Rv�oA+�)�CZAs�zA�n��6��Ӹk-71s��QiJ9̂z��knV��;T��c��qmU�(�KJJ
+l>G�@g�|����{ﹰDs�+��{\a�o��� �#�@;�T6�\-3��>,n1b�����i�; ��JM� �á#):��e�ML~:y�g���i��
�5f��^��)w6E ��:6/D:u��uȻмoc9)aq7a~N�XY����)�WS�9N���5�2bc#�Ԇ��5A�)?�kG���m�t�e;�θ����d�!��(���s�:���'F1��:x����zo�]6�8�3"MGW��#`3��F]������7�$/������eƤ�e Es�����edd�Û���g�G�G�����''lϦ�"�oo t���!8�"K��b�H�y��T��IPP��P�I�w�.��	��h��ѱ�/�Ņ�+��=;ğ �,x~�C�@5���䤗R����8Pz�S��[���E.�RѴ�������s����ɂ�[U^]����gV�=�!������^o�˟#>'v �{�4��))(>��(G-	⭪z�ܰ�v����n��	7�9Jw7�f���o�9V~'W-��F���*�<uy����!-�+-��c���Gm��+)$���Y�l�V�w��v}���gc]�yA������{{�u>�ƈ��<��:*ѫ�#�J[�������"��DЖ'j��e�+��v�mjw��cɉP��	.4ꥸ��pVK�b<�U'b��S
�P��?;o�k'���OACy�� �Ӫ�o���"�lR~=�~hXj��N!i��a]�q��<t5W?hߏIp�gc�}����*eoo?��؜��Ԯ3��!����wHbk;g���2��5����Ejdd�X��F�c���+�-��Ⱪ"� ,v������� �g��tt��Ș_G7�Ck��qn!��)Q~z���Zn�g�9�ɖ���"s��&�*�?47�Z���{v��9,��X�*�WJV��PR�Vq4�E94�9՜�6�{5&��n_�3��~�LO}Z��O\:���{�g�`�C����P�����6��ه|al3�?�^������I������3�;�)�(()_k^C�4�
��*_��OL<���%·r��=�"	D���#Vټ5O��ʘW�ZW�X	`fUU�P�&4K���i�%�E��S�0��s�P�0��:|�L�KK1�9�L,,��by&Tj1.ė��"�d�/�dx)�/�5`�O�/��w�/F
�C�q�_�|��]�u��]H��DT�;xQ`P��T�%��֭4-��Pg�|�0R�2�#:�%��Ӵ�!���I��@�P�,�<9� ������*�O`����b_'�E�b�v�׳��A���k��px��Wcb��d�#��lWUF�6���������>���t�aZ���@A*#�3�}7t��j@)�)��'i�XIz>S3y������1|9�F������� �Jfx��|	D�����*_�>:���h!�j�ܜ������H_�]��;	hq#?o���j��U�N��ʙ���^~�����m�}���E��^����m�
��*�q|���'�����!�&�4����Ҩ�K@��D��ԄԶ�V��.a.��А�4�&]YY��� �A�����z�/	y�K	=�w�B`\8o8*ιIS�TŠ��h9��I�b`r

���!ó@0��rCS��n�9�[ނ���[��B����wO{DV�f��q�]�5DZ�mO��������?KY�	y}��#�r�p���z�mH �����ԤW��VGˀm��8U�s43颰{�K�<���%Yu2%�6+�)�}�FKt��d4|-S����y�����o����^TZt'�$	�R�R��~����^���INj�,W��I:�k��������J��9www�t��[\�1��I�w���\޴�����
AK�5���΀G%�K��|�]j���'c�܉�׫9�4��1~�2�?�91'/n]�|��ɍ͓�c�"��~�iB�Z*|pMsꚟOFbgf���ř��Hl����ǜ@�zhF�|��O�����~I��]�g��x�|`p��]|d$�ڦ*��2��ݫ��@a&�Z��y�;��a��KF�j===�H�9��"��T���'dn[;A��G��Sw=iVx�""$.ŧ��G�6�q�{� �ԩ����JB��7�*ӳ��z@*|i���7�O���p�E-M\
�[��p����������U�5����_ye��VH��[X{�J����oət����\��\̠J��~���4��Ԥz���t\���Z�T�5Q��`E�\9�I�B�+��)��Pq���
��	�B�y��k����&8���'��_��߿�A�W07��eb��/7��e��R��1�DR^F�Z��Kr����/����i?��5�ξR?�"���P52��?�-���p�����!K�9����|��cH�6�
G��pr�'i��Q-�����s���݄uP��=���������J�*�O����55A1�0�����-Z�(�*pЂ�F�}>�b/7בmaa!^�}�s[�P�R󽳲���1�.UO��m��Gf<pB99I��x�4Q���� ���̀�u9�h'��Q�^��_�NiX"3:�����R겙)�޹R�l,w��/]^4��u��(��Y��i&>�ٱ���T��+�
�=���n���_���u��-��ݣ<"r�:������DԤ��qR��G��ח�f���ۖ��A�"��$b��������C�Q��{�0��r�aQ�����.�^�������M���%�[�hh�ɠH;��UMMןS_�"	#ׄ�.(4���75��Y�7(�צ-gfa�n�w_�}F���
��o����Jv/.���BU?�tZ�`��SDCM�p	�J��#�?��wB�w���L
�<|IuKU�re�枸��8�Gd�ڽ	xR�,�BY&4����Gh���7|��'���z����Y��C;'� �	h�+ ���J�=,���>=vL
���I�h����Es|����axw^�Ź�KEh ��&��""�X���(Ɋ��hi+,L��x>�5+��15�:�H��4���̴eZ�(�K%Իܡ���v{qw ��(���%����xH8}Rx~��b�w$[=���cڹ��8��x���u��e:-29�	�O�D�`.��Gr�F�<���C����v	�a>�ԏ8�ډ[�����m�0�\,q��)w?��Y=}J�P��:ڧ׵��q���Ʊɘ�Ɣe�aj�Dj��-���v�����^���t��%c����2˲-SSc���R�V�R�/q�{{1:#&FR���.���Ѥ�{ۦꝲ#,D��3w�Ծ��§�/��aM��^�鬟K�
�`h!��b��O�́���+�3���C˪9[��s8if��j�f�[�I�^�$��F���NN�ߪ�{`�o������ʱq q�J���{�eDR6.&�Q9J��M`[n0.[Xx\���_>�wH��M�&D�_��7�,��^GF~Ө_PzX;����S���eR"5�st$ ��\[Zbj���/�Ё�v��B+�C�KJ�e���mk�n�˻�������Qq\�_-�k⚰�?&���5i�|.Vd�5c]�=^�P����)�J��?��Kّ��?�r\�d�2��!���κqG��v������w@N����F�©�?��d�Ƭ�N��X���N�Q��a��}x��a=�b����3�G8� $�Z��{���,��o�+�d�jM41]U_���6E8B���X(h���
!�����;��jtu-2��d۷�\.(��Pc6\32r[�]3�H���b]hi�!M\�����&�����y��e8'�W���[�j���Q�6]��Vdƃ�a,�4-�����E�t����Z1�>mr9��Z`|�W��Z=���6��a�ݽ�Vʹ�v�c
^JfXS�Q��G�jk'����'���������k�	!�m�z�G����|�����K4G���@@�-�gfޤ��-�<�Icg��.u�پ:H7KqSJ����	l�ņSS? ��'��y�Ȗ1�ħ�
M���Q�,��AZ�w*Ãc�!.������1W::�	��4�[�ir���5�u�NsH�҆��e�)��߳󭕪ܚN��Q�w&r�=�)���Ż�S.��g3�RvR��7�W����UMlC��R�a	_�޹ YcN��<�:�>>��
����Y�|�I����c��{���C��/��r��l��){�n�������JJ�s@���=�i,���!����wh�WU1pr�yvK�b�l͞(�b4c�9�m,A)񇠤�Sb���=:�����L��_�aۆ���!mxl��Q�,�ٟo�ko7дC�)u��q�uSoD_�\��A�����L�Z��K�G��Ӥ�3��͞8i�{mp�3��!���.����i�FC�߭���GЛ����	SP-̾NL��`�Y[�����S�%γ�i,�P�BLX�Ga�E,�g��<a�;Q��Kz7j�n
����v&�5��>���'r�Jڏ4d�G��;+���������;��Y�0�ͅ�l��.e�� �S4�_��ABs����=�C�$G��j�R��c]��mn��"Ɖ��?ؒ�1k�s���dT�҇��AXFW�w\jU�� �=ʼ.�B�!���)v�3O�wS�R	���4u���!���~�H���F�;�/�-�fҁz:�l�$��eirg�_ɺ�0�黹��E"�1�++�"o�^6)6���q�2�Ihw��K�Z6�o
\��Ov__��Gk>�oA��TP�����q|�"�t9��֖��i^���d�d �
�9?CNFF�ɂ����yf�5�Y2���v�-����
��Qp��%��]���=%K���<$P��"��mP'�}� o[�2'כ�Q<lJ��@�k+�c#U��Q����}����S[��.�9�韭G�B����dZ���{]E{ ƭc]M���2�1����Ɯ){+��$�p��Υ�]sK�g�>M�|��b7�r�Z{6�����,��ޕj�+k0{&�HT�%nS��[dbh�����{5�ܾ]H�|� Hc�		�΀�G
G  R�@�x�3	��o<P��Ⱥ[$�,�A�km�"�8�=�����u
�F��+�f>O�f��_�Τ+Z�E���qY����Z,�mjty�**��2�Xo��o �$i��V�q��4���ͅC����i�#v��@d������M���sjc<��m�TP M�r�2���W}~s�ב>�..l�^�H���nj�$$Q�GT(��,���Q���'�޽[}.��B���r@y�MP�������֡q)�Ck��ԋ߿>�x�s�/�@^������;|����Z�e�~���%���f���tk��i.�z�#�y��g�ܿ��{N�e��*�Y2p$�Q'uom?�lè�h9��l�yDV�v��?-P�W0�o�y�=�g�k�YY��a\�Ω�{T'a��k۷�f��k��������p;�����;��;��7B0�C?ڣy�f^�"\@6P%���<s�)��h�Jp0Ć-��ؙK�l|JI1�[q�QW�x;z����>����a0R���-�~G:��gci�©]h�������� �X82uX���%tt��ϥ�o��7�6�g+nR	0�N��MV���NM�rr�f���2uH���~��w|�4���,h}_l���q��qZU����Cp��U����:~'���yOu��'�qq����y���BxJ�J�
?�XwB�?���]O*֏���ww�"|��3�V$��c��a�Jk1�A�����E������9�G]�]GǇ�jh�g�������$G_~1.�~��y�~�R&SD��m����ƀS's�6�jZ#�a��^�"7�h���a�P=�D�ӛ��??D�϶+�SL�{���d�F��<�o�ڱT��ToI��@3u
sͫ+�N䮑�f��,�Mcޝ��u��C�|��\Q���D����x���� b�f:�RO摢���3/�����ǎ���� Y5uO�Cި�g���c�����j����WUz�ȿ���|�����=z�(� �=[n��i�{�9x���߆\k��-H���r&�*S�ۏ&YL�<Q ��g�@2��`n@��:��fk[�:�xo�[�� �2�@D	�v��DY5�3 � �[b���h\4⏿"�H�Oh�
��V�S��(��σ@u.�8R�E6W�#��lE���Z�<�ԕ6^L�&��[9�zPS]���ƺ�\��)�ᑾ�7�߿ �{>���s��(!5�BjiϠ8�iVAABq��"x.9����n�a�[^î�Ы���\����N�����_"�O�C��$�F����%�myNz�70���J�a���������m<`�'KꖜL�{���r'�fwq�K��=�SIA
�~�5��u%>~4�7;ED�=#qhA�l�G���2Vf�����yP�ŉT~�ٛ��ba�"/¸|~�x�27���������i*)�6ݻpx�_Dd��ߎ;�WZS�H�LEI
 �@u_������*��2z�J��������	zu������Y&��C����L����E,�^��Ϧc���h/t6kd��ODD�r���(�f.�?~֠iĐSM��Q���hypȽ���,i%V��-���E��B�O������?z��J42.���j���i�x��@]>��h[^�r�����Z�q�1���18��0�ԮZfA&��Q���1)eX���*��G��d�UWjN��1'�yv�RW�ć`q���iI�CK�m�|+�X���
4 !vf8-�����m$j��)�f��-Ⱦ>T��}���Q)��[B8_J��4�qy��{�[6@�p8�l�{}���@�uzZZ[cVۚ'��%��֘��̿�����k����CH8ۋ��Z����73o� ]���6��Hj)����Xeq����~N���q�K�<��QFbAE�{�����M.��O>���W���혤����9�A�-x���A�O��$�#X��=�V��;zs8����h������g_�:�)��J��E�yU��<+��e���"_3ss)WJh�M�"����y�!3�%��aSo�
�.�`�{}ccg�T�*]��ڄ%�#;੟H�bG���nK���:1�|�o�3�*�Y�#�|�	���j*�55Qj��徛�A3�2v�Z�q���J�<$�,��Z��ӳĜ�$�:�K��ۇ�Kfeo��W�Pu��1��7K\���d�9��߹���ڗM����������J�:��O���N\�d|����Yk����UP�z^!�F�lsII�L�97�N���֏Q�u�.2&;��ɒ���}�N�8yc!�\��O]���%d��q8{ߏ��K0� ��Ͷ6��&�>�����W76�_�/vw+|�x�Μ��A�DW_�H�ΨN!iG�z�9
51����Qg.LZ���������˱tM�G��J�[8~j��N�*S�}�<��≵�!�؆�*F��u���x��	D�2�B#�������^2��]���h����?7ܤ�-I�8/�{D<�4�������^��F��%p��x͈{;����[|��	?M��T�����v+��������=����P�L���oxXl}*�E-·��Ts7��0(�)?y���t��rr~�c���&��3�]\�i�aw�}*/O���7N&��_�� ��X��jl��3U������d�v�a�g��������c��rܷ���%��h����bB�I}�>�0y��r��!s�/��WnG>G����|��x�G�?y�h��Z�}uHH/���������~7��{�M���kb+ѻD�ND�-D����G��-�[�&�FD�D�[��}�s�8�e<c<�^�Zs^�k��ֺM��$W�PM[���������[g4 ������kt�6�9�����cOψ�h�h�\��@'�)tR�X�if�7X2,N�+p�c��� Y^C��Wޓ��i�^)H�[Ě��	x���ѡ��(9��(�7�74pm�\���n�R�$�~������Iz�|���_�����X:
!qJ�J��,֏��2V����Pm̘k۸!f�Y���̾��!��I�L W�Ұ�S��b��I�Ќ���dM��{�:=������`�k�X�Ew,';�Qx��
��@��W�KH`��D#�d;��#L��C�Q��s;�󬽋��gZ�z�3n�8�3I�;�1;�mW>?��R�^��$�"i��pK���t��QSW����J�����q"�6+*<Z'l��`e���0���q���\��ҙ�T���G&�(ǒ[RUђ(�Ճ&ߔX��U�� -��iN�\ނ���S��b�੼`��SD�c�*"G��R�c�T�h�ݦד�ԒI&~����nlz�y���G�t���h�xң���*ݘǔb���tGg]�������#����o�v��7ˡsT�e�sM+ӌ�����ҧa��{w�'�N�bï�I6���i1��c���/�F��N~=���Kx8�?A�T �����l�������ߗ�`�+�~����;���[y�+���g��"ECz2��/��������)1�SY䐺�o~��O�}��פ�xd�z�������=̽9~����A����:��ݝ���L.o�9i�O�vk�u.�8�xB��1�R��8@���ˌ[M�J?W%:�6@7�MM��*/��:�5�7�-Gj��9({s;�'����݄;֙������M��4�i�i+�hiU���-���X�'IQ3j�HQ�i�c���:�[c/���7� Ij�c���L+0�ؐ.�0v��T3��]x������s�Qӓ����^+�Sh��s6gf�Dn�N���,�]xe�Dal<�rtûYLra�� ���K�}��`x��<�����gP��F�jλ�m�{��AKX���P�{Ѧ�
��GV0i.m���Ğm4��6��f5 s��Zl���][�O����8����ո����� 
7�;:�:��s�tv�y��of��uv�*�Sz7.�#�:C�,�u.�<oSsQE��� ����LK6GD,K�ᐓ��:�;��R6g����\����5�z�.�/�~^9mv}ƙ��ӥ�T�@����t���Cf�A�â�����6*[���mEYs󏉷oΆ����}�l6���K��5�]k�O]b�?{����oZ�q�2p�	������T��h���'�j�v^�O��2xJd���@����47�U<~2i~�C���F�lU��J��Q{�VI�u~�FSk��t�t�uG�=)�����d��X�O3H:�݄�/Da�
���� R�D5��8Gt�H�Я���\9����-��L�L����;��}!��  sQ�oJ��=up���%��2�����w� ���T�؊ê�v;��9��~��������2���=����h�`���)Ѐ��k�vt\|<Q9ɫ�;/X�xn��xkr7�G��w�I3yJ�N	K�n�
N(L��q4OM���Sl���Č��[D��� �CN�!~fi��֚4ɞ����A�AΛ�Ɗ2���c��K<�
�XJ("��v�g�t�i�f�7c4y��$U�{�/fc�S��#T�W� �g�=֋m�10pG2��_ں���NM�$���%���D�n�w4�8������QJ��ȵ�c���B��|4PȷX�|�& ԡ� #���3�9u�����?Db��_��~&� �r���I*Y�ʊ��9W#���E��n���S�Rn'��N�k�f�����P��v������$_�W�D/���0�8[�x���c5�59�Td��Ԇ��anT�v����?���ha��s�zn,z��D��x��S(ӋFP����jUlf�|�###�����>Ûvu���y�v��ؚi�-�h*?���*fi>7�V��m8����a���;�[�%bP�Ҹ��W__�R �8���p����$�}#������*�4UD�L��`Y� �B�s��M�"����[�q�KȰ��As��bX��N�EG����K�Y(p?�����۲�ɂR)�, ;"���T|D�]�?Bp�V��U�EI	7�����?�@������/��ݓ��񕑕%̶x��񫑒vY))�� m���yx�vɓ��z��쑹�t���M )�]���/fFFK��R��I�����F|��E���~s�aċP�b��~EZjꗓ��
�����=���]�)g�o�ɉ	n	F/|�r� z���o+[gm���1M�cR�׼���w�&����F�}c��!���{��+,b���e��hN�ui�B!G����F�Cz�<�C�J@��D�2��>(����h����$'�Dm@�paa�=Y�Jc�	r�O	―~����1p��C��b0KVỈw��y^��������m�[�����Q�S�o��_]�Q`5�I��r6�:�ƗL���M��3�CJ�W$������?�r��1�G�<%��lu�q榕������sˮ&!��s� ���h ��ö�N0)_�$e}5h�G��dN���X;n>.p���]����41���׵��CJ�vE���///O���q�& ��Z4�a�n0����~�@@�����G;�=]�;�>i�B� �s�������N��_NL�Ȱ��P|�*G�o���*-�x'CF^&�-������f�b����/�bwd�wvh�<2��-��rۿ�Zߊ83H0���<�9�`��0���І�~=��wvt�֗N�s�$��Ls;l1�7|������#�T{X��5�ʓ��i6�D�H���5	�M��ޅ�����`��KX�jq�u@�+���P�O6$%(i:��n	8|����ǜ+f�v�u׆�䤘����nm�n���z�#���~����
��+n����䎊�''��ι�{y�F���9�&�]X�v�W
�0 ?b�(�
���`A�W#Uo3*�ڪ:�DSK4�J{&�sx������wu���k$��ro��h��w��z���	H��:�ߗz,�� �$6��H<�>ʴ����r��!&�Ud�%���Q0�oo��آZPa���C�1�`r򉘌��-�p�q���l���ߗE~o�|�<�Ё4ޣݗRCSs�I$���o�|�3��V�XV�wK�4�j(e���u���H&��Y�n��}7퐊�.�R�#�}c�v^!:�8}����8�&�e4Ի�o�m�U��B��-T�"Uoc��(�LIM}�N�]a��[*���fff���)
p�nˑ��I*
R�s#��$LR/
K�_��,�� ����� �)�c�QC#N�"
,��"�S]s�3����Xݒ�nnx̴_�'_D-K�����ˌ��2?�6*�?k�h,$*:W���߽0`�C�mF����G�9�]�pg��A���۫������j�G�s��B��Nea��r��%��M��D>޷
t�FmH�c�ٱ�{ˌ� ���T�v���У����cct �������L[s����s�Ƅ��yU�{&�]|]
�]�����@�K8��1\�oW�`.��������lL�b�W��g�M�
��hL>c#G�r��{'�JJ��h���7u=�o�\��x�,���/XD����=�#��˳&���M7*ߥXMx�HC�"�g�T��ERcF����|���w���T���U��夘e*���R��a��C��]ϦnB�	'�y�4�_Ic���K�x�4b�/95�'w�-ڀmLΑ����&1X�j`�#>���ޜ~�ez�K}��%�B�b��ȵ��(��^�(�_�'�ݹS��������B��`T:@{	�g��Z�0R�im�C��sg
��c������` ���@����#O���m�(.(����|�nEz��*�6f�/�v�~��~���������M�Q�����KV�;+*�x20�?�&0��Iʗ=X�n�j�罯��,���Ƌ��1՘R)�ć��>��ݳR"溔��(���R�O4>��2�Kd��~c��a#�fUX͊�?'�ޡ9܁daN��r2a��4���C�� �{ﮩ}.���v�9~G���?�;"�+-�S�C�Qp��,��C����o��k(2��ܸ��}�]x������cMr�?��l�G�?VZl0��ueD]S��\��e�փ�P���W�O;/5Wd#����7..��IH��eE����>�ԕ��nN7��+x>�|�{|o����h�ܵ���w�ܡֳtY٧k��s8;{�W��H��԰"�r�{��+1�B<D"Fi�?�*�:z{���m�}�-|0բ��ՑZW�\�%�m\&�ø
D*�4��kN����G��i�=�f-�:5�$ҳS�S���y/�B�9���c) |�bꂕw��/߿���8�:
��XQ�\V��MHȓ{`�������S�����ݫ����C+)���&t���u/���M�UKo�Ͽ�����(��~l�ٮz7�n�����ѳ�f;&{�+Ū���9�(�okk�5�1���VEߋ�^���z7�Y�8[���3��140j�G4d	P��^��w��XG������S5�����EҨ�1�$_cF�d����?Ժ6���{�Ux7|å��^�5`����X����[�ty�4��݄���_Ye����J�.?���,z��h m%����%1qq2�t;��¢9�]��55���"��b�?~�4�6$�b�^�����rQ�~_~#3)A?�r�Vf��2	/t�֗���M�놡�YX�4z�X��RT�	HcTrXD�o����p>�t'zIN�wǗ����`�PlZ��@)$�3ٹw� *���O�	�nl����������\m��^����rj}dXD���Ѷ �x{pfs�$�[$i���ݱm��O�Ē��ɔ�����Q�m���'�,��Ճ�����x	ʣ�?JP�y�|wЀ��yڽ5({��q0(��r�ǀ��H�hH�PkC��1�=+���ߋ����[8[ϱ�ttH��#E)�0�G|��= �,W���y����=���}���~Q������*�r�֒$��Zq8�Q�H�\L��e�l���8�"$�5�ހ�������f"�����:�o�1',�I|������n���O�%�_+�3�Q����;G�������
!A��d�>��74"O=<���y���ku�'p%�/{JDQ�_NS��8�7_��h�=1y�@�q�w�Z�� �Y>�g�s9��%`�Y���<mYW��P�/Y����T���ҽT�5��
��~�G	A��8��߅_=�4q���]�ϧor���i0�[LU)x1�{��S33���jf��^�6��مȈ�uG���C�/+#K�z5�Տ��K��v�Q����-���������vՕ�R���GU`��ݗ����>�vc1Ak�)o�'�58�I��ͤt]�c{܇��!��4�.H%r'���G�@2����[��o�����۳��
��Y�Y�$��kbt��R��{q� $SU���m���mւ�rr�o�%%p�o���^Xu��4�����z!��[��-��-:%��2���:��=�+�{�h_���B�3��%m� "66�~�\=3���s$�Cb�O7��l�SA�~�׳[����oI�Q�JF?^�Y�����"�6M�\���L��省���y����j��j�d)! ���O}��j�沆������cuEʉ���"�5��|�[�Tnk i?���k��^��o�ς���[&�vg[q��Hh��#�k���MiR4#C�i�-2�EW���	��@w�<�J�h����\%��s�$L[����[y�BO4���u�ws���3���U���@j=�����S�Q�/�223#���&z�y���XH1/I)(�q�»B���#��������ZL+�C�|�)4`f���')�R'���XG>�ծ'p8X��֎|���_z�M�H��}� ��뇕�=�i�T�Y�8V=%�(��g��ZEt�C����ͤa�:�S�G`a\V���pK1/4/O>��8u�W�;ZW�{Pt6�F��}0~7�¦mgxuF��k����+���I�8�NNq��Oc�����eC����n�z��?{��x �\%��z�
�J��ٔ�	�]�*�����`�i�,�dƧ���ؒ��f�ݮ��b���|�#�"�B�1�0���S|D��:Q+&�p�K��J�v�}����Nʫ���/�6�.��pz�ϝL V���{��cw�fׯm�۲ӼO�W�qk�uqm�C#�휭����P����`��-鬟�������+<��8
�����JJf�-U�0���<Pd �&F�}��mr�����D	�~��f8n9������1�V'�n�W�i��UZ�!6��K<s �d(v󎌈�>��YX���u7�P��^6�@�^�>$�B��b�H \�����CCP�!u��E��,�kk��YV;�|�:(TT�	�:��íYaM���'zt�--����q�zh��SB��'�ij�U�?;�׷�+�
��Dh �xJ�-����	r�4��+I�3*�A5|��!��5aDR�H�����~r K2������9����Y���k���XŐӁF �f9|�č��Rvl�e�0/hB�����ID����a�ũ���	Z���S��Sx�V�-62���2�� '�=�4y؏��H�T��_�3�p.�B����4t�z�V���.3��O�]�����Z�I�Ν�¦�4�w��D�B�w$4��'(��j�"�5=�K7�^��$��9���ǾvW�w��ty��E�(U��JGĬx7;1�B����5K��؁����G�`�g��@.�ly"�yJCc�\�yfFoa���|�nD��/�.�F.GQ�&+~�P�:�X��|���j�Wpp���Ы.2$\{1��(9L/U��3.����W��O�+X#��B�*D��S������x&�ge-��n�<5��ǋ�>Zƴ4��Y��L��0��i3�)P���5D�^B��@Ϣ=�Gf�l,�|�.�VbB"*��^�vͅ]~S��?���2��@�f�оѿ{$�e�߇�BC?��k�|�y��[������^�4����Z�0�W�&-Q~_K�U�K���Gcﯛ��M� ��D�4��qr�7�\�^��O���@(��H��쬼D��}�+�$�srq���h)Ҝ�;S�^�,r*�8ON�Ґ���"���{�ѵ�7߬�A%��-#�������\{k����Ɋa� ��`�3ӌ��8��~ro[Ú���bZݣ�����6�>�FYޝ�>�RT{j����Wȁ��!�'� r?��v%�$r���L��F��*�m�z!Q�����7���������(�)��V#.J+oo��B���ӧ#�Q��W�%�ۺ�?�>�����ke�F\||�_���֐�ŚlAK���Hd�Z!oi,"kPX�k�O�������F�
��n�@b���=���J�SĪ�ȭ�����D8���g��(F
9��[�v0}�&�����mё����G?��*Ddk4��(e���3�Hd�f�w�9<�m�PX� U>�;a��Y��ΐL�@6z�H/A���$��K��B�Y/'��W�b�=��R��mR���M����V��Q�ּ�?����0��;��ڧ���~�7�aig�d\_�OC��W��ŗ����n	��Gc���X�����(5~�D�b~&X$65��FWN;�阱|j������QP��f��vr6�/�{�Y e�2g�}Nh���c��G1������z��m���u��4��«��e��z;7N|~������ U�mF��4���Q読��j�A���3J~��t�u� ����(���o/":��#N���
E�T	dNxP����WRP�GO_���MW���{m��X
p��U�O���tq���ɡ}�7�/X�J1A�#�������s�ef��I7�F�u�&þ�c2�sw��������:5���:���O>�(%���Cc�SdF�������Y�D���1ǺR@}#�����JJ����@���d���[M�^(�Sfo?��ini��O�͝\D@EPh;��]��[�_J�Y���\��'O҆��N��q�a���D������u�ua�K�� #�Ao��| ����l�	x�]�W䙶02����Ä�z�-i�F>%6��"�y>r�3�v���(;t��?k~|#�V�5��H��L��8u\_6pR�^9ZU��	؛�,�J��sQ��� [���>Lѩ�&,6����&ѵ�����u�ۦI��l�P}�	Ѱ�M����*eY�nxߪ4�kV�ٚ	B�	 ez���@%��$:����D7��t�nnH+�܈:u�5?j�ĸb���N� �ؓ�?h&!Ē+�7e���B�ofvU�!)� ���f�'q��v�y����PoZ����E��޷� ������ö`�Rt.�q��a����?��8�����|t��|g�g�f^���3Ms�$H�<����D	Q~�=ܼ�C���
m֍�y�e��4��@�)��=��-),�ظ���b�@�B:�cR��w��G!#+��������4O;IX�u2h�_��%�ܖr����=��OMJ��7�y�ɋ�J���Ò��v��6����4ޞ�FA�<s�*;þ/����>���k�R@��p2����'wN�lLC��])Z�`�F4�?wd�^�90� u����m��>�#{�4E#k����&��֗����ﰰ �_�pU)��77#֦�E3e���ð���ŉ	r4�_�z	Ҵ����pd�M��5o����M@��ܱ��(ƨ��H�_T䢬���~�/�/�Ș�2ܔ]k�9���J��-kW���Û�T��rE��>o��J�q��� ���L�UkAj�xziY��I�q�q��vG#��lm��%hy��s5�d�}ҭ����o l����%&Z��0�E���xfvV��*lA�#��Q��`:�	y�e�h��U>�����V mTP�$w�E��-�rj@�Z�(�O�;�Id���֯8d*�ӱ�[TK�waU�_|C��G�]�����1�0)F�J�;��&�c��]�ȑ}��Mr��J2*��d��c����h��"�,2fc\�P���'��<����#����R���&+\��桻dm��kS)�J�����O�s��@��JV�o��>�D/8�������ml���{s����^�p��eD��9�W�u?u��f�tÛ�<�?p�<��y�81����*7�k���rȠ���x���f�3���]�kH���,�r��XJt	��	����������A�e���ɴ�B���Psv!�N�	�DOg=��g�̏�����䒃T�J�f��������x��g��U]��E(��o0�D<q���GF(�F"���2||�Q�r�O� J�D�g���$%{�j9��0�l�c�\Ůէ	`Aً�O9a�YK�.�*7!�KD#�����&��e�3h�إ��r".̾[��EQaa7�w����	6
��K[�At��e�����i�=?Xɚt��᝚�W���ec��ϣ������A/��HJJ�Tļ�޸��"d��=��߁;PO?�I��P��,js-��I��AX�Է�s�.��KJ����oƿ��wz����	��%i̾�� C_��hr%(�w��/��4�EE��@A��&�:𷸟����P�k_�t�2�I6�&�۲#���9$+{6!#�;W�󕡭�<T�'X�hX����H5	�$�dL�}�8�F�����q�k�|�:��S��j�h�_hQ�gӻ���@��~${t��������\ah+�`�U�������;��5O	1�q����k�?�D~i�V�}_|K���߇e�|i���XevKmaG�܆�vב���<��GG�}}�I�R6&i���ڶ���:�y`����@�A�@g)2��lo��2W��qUm�X�o2�b�h��.ہ�R��>G���
���#�~��}R$K6�am@sc>�*Ж�OM��7��(�I&7T����X]-=2�	KQ���쥆n�GZ�q$v��$4�1ęu��R^��G�c ���sB3�{Cպ�n1	�X��N�}�%��L.�q>��b����N0�����lY��ɨ����e�^G|����c��E�n_(��aUb_�"�R=	����fc�O�f��34�FmHc[]ň���QKMyz:>.9�=���8�>|Q�P�7��U{�-}gb�{��nM[񊹻�K|{<Y���#�����oT�q�MO3�S؂�J��$`�����]19>R�c��`�L}����,�`�'�/�#+��G����^4>mfDf�5�.g���Œ"h]E�l�OE����f�5aqP$,�j �6úc����S�Y:6)������<I�o�;9:����4�!�WC8�f���?/i�ˤwG�Y��Tq�/`0�s�=_)߳����i煱2��oi�s�@���G<e�	|Y����}�r��`��MWW���z	�ck^n*+SSR�|�
T���Ǎ'/4x��^����O�t~�|V�q���ɞ�q+9�*�a����Gl�������!��=�fW����@�c)y9n�N�u/�0@� �G7�|��m������QǺ�k�Ƽ���B)� ���Lѫ��Xc_�g�0��fY��|)�&��w���3;v�p�*�p�^m!�,��J�]o:�����Xw�l/�Ј��� �y�>�N�ƕuk�%�S8MAs��{�Yf�WNBП��������KSb��^���M��MO�Ɂ��ŝ}�?�����H5G���$+:ÿ��P6���Dr�2z��ѐBw0���A(a�\ ��V��c]*���/��:	�b:%��t$�s�x둝����\�;�U��G���߁��y�������!�'7�\��fh#Q[��ve��j�!ܦc�h�ʲG��D��	�����)]I»\��������`��ә��nړY߾ 0�96i����I�R���tE ҥ�� 4T�a[�+XR� �(IѲ��㣵����8����"�e��C-��5���e3l�k�Muj4�����cy97tcek�I4O.3ytOէO�w(	�$$>]y��91IIa������P��tшA�c##jNb�+c	�ˀV]���|��^�S"�� y�`=S�z�w�_�٩��</u�B�)�K�2K=��'n0���:�:��.8��"�΃���f:�j@n���?P�L��H�����C[[�w�<24��'�D��2��xY׮&�xD"ɝ�%�;67~A�̠%�=��y�8���I��Iu764tLֻ�B}��Ы�A3���@�,��pȊ��Y��DƣǏ�
Y��m��댾_��Yɦ��r�^g!��T����265�Ao[���4�iD.�t�O�(P������C�RN��#�~�Z����4�$�P�o�V"���m�"`rg÷bw��1��!�-u:Z͵��#�/#1��{f������I/0���5�qm|u�K&��_�� ���?�E�����A�.�Zk��ң�#�`�)�YC�6����5�>4����x����,66��"�B*�Ĥ��+"��Oq����t����t�%���7� "	a�MEZ���!���T�5)$���=��10��z���Nߥ�����tm�֪����p�Yォ(_����^v�ڄh��ީ�:�EІw���pQ�������*>�|�߶ߍ��FT���5X<���H�`���J�k����?:~ed<��Y�%��?0�3ߤ��rlL�0�yt���������] �?j�|[�w&6I�,Щ�g�O�dH���0�)O�)>��0�����g��8p5DRC������3�:x�h�/p����aqnBC?� �ߊ�/z��~ YJ��J�����:��u�#"���<�.K�(��cZMI�Lc�ZN\[AT嵭����
,C��<=��c�{��xn&9o.7u�2BY���\4�����?_`#�ɑH�cBa�^QwZ��3[r?:_��*�1�<��f�7g�}�k`YRn�����{lB�1�m�.�w�L��l�h��9�V�@���
[�a����lƸ�����G؛��楒�]\2���4�4H���-%��_�񃢑���"riO�bJ}޻9��S`�<�ώӞyy�$����A	�i��=%v�v(�S����]f�ꊡ�2�޳gϢX%���t����*�\\����p5-X���s���^`P�,}T��fZ�)�x��������qz�x�5pS��|��1��������� %C�	: ^�v9������=��l2��--�2����칛�y����C��Q~\}���ǚ�9<����t���������q����h�>������1|��
���^� *x�T���D+�M��^ sO����������(���j��k��{JM��@] �d������ma���XX�;�;������A�]��r ,�oơ�(��T�?��`7�+6������1A'Z	�M�G&��2!��{û�K�^M��u�v7%�+�gk�����]�ul�z=��Mz�R�v�<Ffzu5�w���>̴�N[��D*�c}=����%yk *gs
��\_w�^#�����Au�io7fNN��K2Y$��"���PM��k� נK���N�+�	�-��M>dުC�tDP&��餫�¨=B��ˣD�Ք��'���>��ݓP��P�]�]��Cm��kfC$Wm��c���(�q�z�o"�ڍ�<������l��Au� �aSkJ�Xaaủ�cyc+#ǁ�;[�e��h0Y:���Ι��d�7����"ꊇ��)�[�R<��3��ܙ��\�:����o�r6�A���n�����}�t<��'���
�hܮ��������g+P��x�5/ҚL����,�s��cwH7/�Ytd��0T`oH�b�|^�4O�\�N%�J��<���G{�\Z�6sMU��6n+����N"VPK�l{v���ɶN*�_1^.��(+J&)�kɪ����;�������n�qA9�p��]E�Ũ����⏬��}4�R����wa!!����5��@�h��E��z�A�E�3wnj4���L�Q�b�?��ገP#��D�g���w?v���y+BR������uT���Ń�X%_,��������3�v��?����h�N���Ŷ��1���p7/���NP�B���5�#�WQN��D��ߜ���2�B��y-�����'zT&h{ěۤ�r�N�-k4����y�[� � 1~�/�7ʾPc㪴}��"H��R��A^Us��.G"�^ ��=�:#�	��uV�Þ�2�T~�t��簳,�0�d��uLE�F�F�[���wI�(�(�����r��� �F�u��he:k��8�O25/!KN3�{�n���>2K�g���|ӿS-������1�^��6wת^�M��>�O�^k��,=��i��Ͼ��}?�H�@�~����GxW�����2�hr#{�1�)���^I�<Ylm���fXN!&��"�����Τx�=u�%.�9�k�Q����Qd���C���F�r�����Ų��>Ǌ�[�e2�����D��]s�,I��W~��Hw��7�����)$@�0�)�TF�����[
!�}���F�N	���R����tO���waŶ��"I�:Pu6�w���p���>��l8+��M�*�+=+9�i~-����;��Bf^2�a�%������V���iNS�9�i��ޞ����Z�x�"�IKQ�e��M�͆���1�ԮEnb�yЩU3x����HZ�ظ�,�n�d�FE��E�v�V��IC��T ����l���O}��7���Z�N�x��W��8�k{v!�<_8����wP)�C;��BT�P�Z-���ocǵ�ܓ3NJ�=��7�p��D��V~�,	���w,Z�����{0/�O낱|��������<{6G��	&��(f�������6�C�ze��H�%�FR"< ������A[��b���U��7���j�y�����ꌨ���n�z�!E;~�/)�e�������|��y���,��ȭ��$~k��w���h������zM�H�^�H\yH�gU�UX8J�i�:�lH�do�r����/�F�.��s�_�wͿ��7��:�v�c��i�4�O�#��~�?���](%~:���#t�w��;��]܄�K���#/�4.ѿ��Fq#U�[W8�����5Qq�}��M/'�1t�l����g�wN�#����vv�3�"Vӓ���/+F7㙤�I��x�����K�[9�����,>B������3�3m��f��;����W��:{� OV��k�z�O��Z�j���� 0QK�I�#�+&��όX2����70x��YnҸ�J0Yz���қ�a4�C[�.�;*��'�A"de8(2 �($�nOk h�'���t�P:�����₠/FO�M��s���)��6����eNsN���H�+����t �Un�{���4��[�u�o � <�����Կr�/ٰ"%#��ޏk�`Mo��ӀO�Bwq�,�����"�s�-ػ��赜�MA�J&�d	I`8�X��ӗ�1��5�p6}�0t�`�ÎO�7R�#}�(����K�(Ⱦ��
ߴut$���'�,�FWXD���e{��}�v ��ᆔ�L�@�����B\l\�����֡����q}}}u��hccc�'����˽}}Y<I�s;��p*���8��,�%R�D-�;� ��i>�5��@��Nwx:��J��772�����B�xS[�����$�3��_H�t�&p�y?��Rґ��qo��~m4�y��#}̨@�S��PB�]dn�q6���)��� ���x�iF���<#�C���2�_��W�'���2�����W�t�ᓌ��LNN��>���b��[��YjF��-�V���զ��t��k��i�s�*�6�r���Śbz@oN��
8�T@k&��d�j��XN8GwB.�>-���umb
;
�,�:bSJ}�֡=�;�+��0�Ww�T%�*ec���}�!���Df���[���/�3R��9���W�vu�:����ۋ@�N#Z�fڂ�4<�q֔����|��*�QP`5	���Ҿl&H�ΐѕ�J��Z��'x��]'��(0��Ug)�A�=�n%����D_!+������0-U���N�E��,̥��L{s�?�9����tm89e�Z��5!%�,!�<�dl��b�X������u��^ǳV��w����X��c�'j5X쫙�����?^;C��䣷�W�x�o-����(_JA�f�����a�`Rؘ����ޖa�־�!�X��:�`���R�*�jEB��5�I�6"��n�x���7g�,CB��&��*��X��##���+82��MI����`F�'���nQK�,G�z8q���D��7t�-�v����űc���}�(�7n��R�#���o`�>imj?�����y�d��T�̵�~��y�J��g%z��^��J S�C^�9Z�~$��"��2�1w`te,��Q�Va�3�a�x�3X%��}r2iU#{��&��>$�C�cza�����ǁ��7��
jV��S�X)	�lY���;�K��
ᔕ����s���p~I��X��mk�vP��20@�������P3u�?���.nQ ��I��Hcy&��	:;"2���փX��ӧ�u���r,-��r�\��cS Y9�"����1��J��7�'7��������Ve]۶q*jB�@�|��*ҋ�r#����%h���\2���� 2Z�ɵDi׿@'��Q��¹�lYkW]3�c�����'w�Ѩ5/�Ҿ���G>U��;�J<�^��RcKӗM&��Д�Ԃv��>�/kJ��eΤD{M9�&�~,/!�T����/��`4q�p]��R��o��J���gn:�:D�(�=����C���&Ly�Id�����^��O��$�f�hL��}k��=W�,)\�	lT �db�%Qw�{\�|�=�s"�4����Q=?z3��Dz ��GC�6���K9k�6d���wH�c>��$ߒ>s@�OMA	�^�h䫮&#Ŗ�����~/i5
������W8G���pI5�����<E�i-"ݶ6Ҡ��E�wˮDV�Û�ßX�p?��K�4���]�5��-F~�mF��G#5<�ڂ��b�#)���-s� ��Y���o:���5�J��iSG�b	��D�u�Hd�`�#c�bz��޴*����Y掩)�E�:��A�pF	O����L���==�P�!�����$@R�L���TdUӟ��L�f�H�ݞ�ꩍt�^��(C�p�;�W�`
�Q ��3�C�U@���[��tK��'�n���&j��sGDH�ކ]�v����p��N�$�;�Ǚ�\_7��N��&40�S�R�Ew��-�`�^8�|�~�Att�H�����r���ǖ�-��-5����iz�e7����JY�r0=?{�#	�EU|�=����H��wz�MC�m�a����!��v��3ц'�v�M$�R#�<I��M�	߬>^v+wqt���������/�|��XX�.JS�e���@ݱ ����hAV̻T�P�l��.q:,|TY�����ܕE�N����)R���{�=��5�W%�n?�)QZ�����}��m�'�NQVv����ݦ�蕍XE��\	���<��k;m��4� ��]YbɄ�盽B��l1a���J�R�E����dx�[�i���%B��V�)��G���ל�.�g~�e9�xIH_��}��d�__�"v�Fu�#�X8��q��w\LU�����G��1Ҙd�\��F_@p%Y��x���k(��Qy�8kr��	�)��7S[݉7�]aʟ$2���P�5���Pu��T���?""�ұ�U�8٣8�3#9��(�H������22BV6�J��3�w����?~�[�ԍӹ���|<��u]�Wγ�ַ�<ob'�vF+� �m�<�k���R��@ʝ�:����"\Cګs�7r�X���*C.6�fN�� y��l}�:�IO�S�2o����R��F!��ռ��Q@F⊐�u9#��F���hV�h.�K
0Y����V�)�V5�_����%��O��3t͏t��q<ڪY=��c�#��-��gX1���V��w��P��2�����+Ȼ�z�	�>벢��z�����[��I�3��{@{څF��\�(�I���y����VYuh�����8��l����J�Zg+^��_X�1��_= �
2~�D��b�A|�̢�[�յv�$)�ӬXOㆉx<w��e��)�4+��e������W���uiV���[&u���Ra�=,{(���'jl�Qe���kn� �������%ý�%�t�ЙtޘC�ﰹ�z�,#ic�73�u*��e�-Йtv�!ǝ�q]8I��L�F��v�ߑ��y��C�E�����6�P����4�Y��W����)",��L��t�Y?��[!�$����y�s�8��Wj�]���6�њ���RKU6zѫ.e�)}�M���ڕs��X��/�;}� V������m�߿�KN�=緍Cb/�fЍ�D�_I}x��K��J�i�y���tŘ�dt����)�S�*f�G�-܄���P�^+�u�o ��;��X�$������#W�-�$�����͹�\���;.���ƺV��٬����z�/����"��4*����$լ[n�X��h����Ak��F�?KV�!�q'1���P�+��*C�"��r�6�����2Z�� {�cc��s!V�OB?h�1��I/�#��}d3�/g�`3��N�-��;ԏ�N.��E��a �$k�t���R>���Y��1�2}X�W��z�&A���ѯ������tҴsmOr�fi+V�^�B"r���ik�ZHɩ]*���;#�~�GS`�swY-;mHd���L��d���n5�Z��=[[(벛y�>,,�X%]��q����[y����irE���ٽc���9��hJ¿ou��b�Ƴ�m�c�
��z.V$��~�D���Q�(�F+��y\
H�X3����{0��p�Ha�snW���h7���	G��Ɍ�0hJ!
j{��_}D���f�<��f
�V�s�E�<��u/^�3��o����:u�}�����U��ޑߏ��t-�+�=�'�ҿ������d;-����n�9:�yR�뗗��Dk�+�ѧ�+$#���D$�j�Я)7���dYu��nq����W�A�VF�-+���cP/���9;\�S%j���|���&�Y�?�X�O3a���'ߗ�I�057o����6e����}�n�JnM�� ZG�	T�/�Ɍx�F�3�4�fOڀq�(n���#�5<��$�F�k��~��+iLV�W�����V\;�)K{:;-����z� ���`��QF��u��3 ������ɝ�o�$����t���d�'hTX��nI���δ��� ���]�����GT���O7���M���5�|3����; ��<)�S��{���u�2��nթ�l	�����s��|��&��T��;����j���L����ҫ/�2���	�ͭ&R �����+#��x�e����ڢK0͊�b����T��h�K+PI��S�4�׀|�)���"�m/1�H�`��%�>�_�㭮hg�I��klW��I�ۅ`��@�S�ݢC8��N�o���m���L�?�������{!�Ҁ�z����\\:	�q��f%��ȶr���]CP�.���!�0	��&$\6�k� �7up$J�׉��Y�����'�`.�����gS��%�'��2��?�D��N�Y?���H���?;?������m/��G�)��X�ʱϏn��]�b�|)�}��~��E��v٤����c���+��F%#����i����ۮ�!�I<�h���5N\vְ�>D�P�z_���B8%�eM�;�����r2Q=6�0��}	+8x��QGl�`u���NB�͗�	>&˘��A~ͱ��Ԟ���y�X��e�]i�jo�G�[*��-π�a�������4tZ̪��R�-^�����̩y��G���M�B���ʂ�Z}aa�l�w����e�n����'��J�C���H$�TAg^�]�~��5@w���H������w�sN�/�L��"ږ��iپ��z�7����3��^i���H�2�.��aD�t��#�ҟ"��k�4}�E㕡��7PI�
5f�H�G���!�W�/��Hר`g,�������hX�=*������V�hc)�F��_�grgU-����&k�1�{�	$iؽ��3�0i/W/`���r�C�4���A���&� �0���V��3ir۬|�@����Is\o��T���3�6�$�'��rzl�X��8u|��߰��NE}�
�n���2wK�Jt@�+�3\���쯨��IL��w���N�c�O�G����G��Ľ!W����cͭ����+JFn���X�~�W\0����EQZN�20��j`#E�?h��o-�-��DSL�|�J����F,�	����;V�m!���b��}\��fp���ͺ�)�pd�ud�+�c�g/M�e�
�I�Ubo����M��}ۄ��\X(�(���X��g]��]~	����ͳ��KM�iΣ�o��Etު?g�x6��p���E��W�g+7:�;��><3���S!�t�~�p6#bFjj�M����
�Uе[�m��j�>~�حH��߱w�@�6S9}V�c��҇~P��8��e?�2_P��4�[2�y��aB��ƭ���m�D�7H�lJڹ�>}���6H�kƍ�\�X�t��оTފ��ă��6Nt��J���X��M��7I��$���E�T�+����k�%7������~Z�\\���>`�V�P� g�j}��X� ��Q9˒ ujW�y�;�W��B�*�@���`���_Ǯy��2}�h{bD '̵G{l�:Lsp�2EHo���{6Gk�]�d⓻�29�ႋ�{骏>tdg�F,d����:�wչI�z�ϋ��u
��u���uNQ#�SyB1V��!��c���8�j	Ų͍�[�2˒vrw0A�mq����{�^�ƃ��]��.7P:�`{Ȁ��/�my�|
d��߫Y�,l�-���2����!�V���'�.�L�2~���
==υ������ �L<놖�7�ێ�6�$tx����c*A8���!dݒy�)P��#��pI�RAc$�Ї	�Y������&��e�]����LT���<�C܉�R�9�ߘy���^F�'�G �#�ق\|Bm�9�:�ӟ�S7��Ҿ_`�TX�ǡ�~�gc�pE�s�
\Fi�P#�uA�$@y��W��JF`O|�~,�>�Z�����9����2c\��X�r�t�������; �UV	}���H�+�g����z-�����B��I���^1v��ؽ(�=���j&+v��9+�ܫ�[:���$��<�s>f�����?I�߁��vx��7Dk�.��7��}�uI�rל����`�nʛJŒ*_:� y��͂����`��ۼǇ�{z3���Iz�$�yX�ڀV2�sv�	:��=΄���(�M�Mm��B�R�kAb?q�ċ�����3<4#��5�!M�KI��N���.N�����H�	9A���0H�T1�=aX�����v�魼A�?�5�qwQ噤�II�W�x�P���e2�>����XA!2�yW6�/����s�d޽�BZD��*�i�H�S1�1/p�/�
��+����m��;!�V-���b�p�N��*׳���N������P��C�^���O�5��,�->�A���N�x�F�����] �|�τu��K�i��^X�:�e�Tl��,�z����"o/�y3�r�L���.%<r����r����&KM� ��n��S�M̶�ir.v��qmT[h�>�<	���QLi����i���EFYי�0m��ؒ�nJ�(�Z�*_��1 8�*	�&L�X�i[�W��бe�`�>{r���Mi��R�� �K
�*V3崜�1g1�B�{�5��1Z������Ug//��G? r�M�����yjʚܹ�0U�QT�&S�E|y�='���D���?�c��MZ�)��x���q���c�ǼL�;*�n��mn��${԰7�24�XYJ�?%�r�T��2	3�":,�����땒�E�@?��Γ��Qg'^�;V1��z���ݟx��q�T�ʐj�����|Z/��2� ����������P�"yHl2iJ�و�h�:����|�D�@����E���I0��cP�`��ڀ���]��`�q��ɒ�ڞFC�`΁�U��W����m.�ۡ���/iVv�~=i���S�F�03P�83�*�֩���,(�B񬻒�)��Kߍf
&����+z�Rf��fQ��޸���+��Z8����KV?��g˭�f��^ '��ʍ��u�jMѢUb��X�K"������l��:2Q-�StYBNꚺ���A���
J������bx(�����嵲B���9��馐�]�=�^���W���� ��X�%ɒ�U1���.�/�x��!��N��`���Y��E��|�_�Ы�Y���G ���+'A��ȳ+,�*Q{����a{J�ǚ�ux����a��vv+#
���?*q0x>F�i8Z�N=�\���r��`���E�k�+2����%Lt��W�̈́g]��L����.�?Ҋ�4��s�[����hl����[T �O�����1���w�����a�`�����Z��	��\� y���T�g��G~S��ض������/����6(V��w���.�E}�g#��n2�4� Ӆ\�5T�j���;�J�Uk��;9=�J��O%[����_�#d�6��[<'G�j�L����4��+P���z.�`y��"r�9�ED�j�Ɂ�f��Zӷ���=�����0���_\���M��|]�r��2� n�B-]z�U����������#�%�xr�ܘ��whd�OJW]Fy�}&�j�g���R����0{���Ot���9��2���6j�v�_�y��Eͫ��\0�s,�暦�8㳄<؞�]��^`M�2�{����6y��e�nH�]�������ݵ�w�yi�6w�F�@찕]���/w�����,b]��GG��'
�
�yՌFkv�~@� _��>�*���O�ʝьqެ�����^=��`��Wߚ*�v��w;L�l��.�2OA	�9��͈xl�#cc�I�۱�x��>"�<����9G��Vo��O���a5���ӃĴz"��u�ܕ��mDG�k��Q����30YJ����/�}q�5O�x�U�S�R�u�����.H��ѿP�Ԍ��hu�4쯞e��0�Pף�����L���q��h�M�޾4읏lȝ;u�ե��Ti���K�����۔�+?]��!}v�S�rNIXe}�eS{�_�������nwF���<��͋�������e���P�{i�D�{�e_�P�����c=q��;A��9p����z/A2�\����rz�Pc��mRc�|r�ax�Y�"l��w}��Ŧ�m����s��8���v.%�O�F�.��'���E�d���2�v�������K�rZ .�Z&}h9Mw&�������!颹 R
Z�¤�М��Z��(^ �C�/
�g�N���-���f�]Ÿ�uv�=��ec�������˿����Ț%kP��W/���юsT��n�ۀ���fP�����n��J�H�q�u��G~h$��:r� s�����~����3$�Łb-����A�����̿	���׈*w���M��װs;mZo�%j�Y�ԑ�:V�	��J
D�dO?-Y�����jiC"�3cw�|�6��O�/,CY�-X����?����h�������"Ra�����
��"m�%�^��߼q3Yږ�g_	���-�ue�^�TW��dӔ��������8&Id�bA��_�U·����h̃7��H�����=�2�����ꠡ#�uoh2�O��e��0�q	5N��՛آbڬ���9@�h*��}�(*�����O�g=��I)��&M��p��FZ㕉!,c� �X�q�(<��D�~�������nE�t!��fǭ�y�1��q/�,����]?~��bۘ'̿N�]�.����ej�r˰��|	EG�x�؅,=�M�,���\��){&�K��[�;I|.�4�W�H���I	��MM�q"
�8cv92��A�ߒ�v���|5{�'�o�ԩ��x�$��%%v�����!��g`66>�~ν��´�e�b��6�-)��X�1�)![�o���y�=$Ĩ��?���J�d���u^0�����7��)��9ɺ� 8��:/�
WW��r��p�{�MQ�����h�dL�t>�'�����
<P�}��$�ߤ[$�xՂ�E�M��� ��Y���I�.�-3K���Ei�`�-Dy<��RBvnmw�M��E�&���m�(c�z<�w]Uno������>�.뛢M�J�H�v��,��.K8��h컸8P��P1jRV��+��^Mc�˲'A�f2v'�sN��$Ф�?D!>�&�o)ǯ�脗�s\�a�������ܛ���(�|�~&�~�sl-f�=}~J��'������4�4��"��o�=���*�ƨ3��>)�*�f3�汌g��G"���`_i�t�[)��Ő2`�O	���e�A�������A�������Cƅ��s,*IW�x�,��YX���Z�e�새�s�2����@��VAW�e�b[U�A�%gkiI�>��7��:}���^Ún$�*�Ә��7~Pajj�<wh9�o��ɹ�����Qby<Ww}`��0/ҷC�z�;M����(9)�����W4+nXB�쫦ᳫ���#�+��.���➝&�y�A��'�k*������zپ�v{?�����U����jS��ݽ�/�W��7.�Lr�1�����w�G��e����_-
X$fda/�d6g�ͮ`������oy*��hp�u�v�;��n�L�%ʾL��zy��q	>�:�~O�����9�
g��/���a-o�������nb�2����su��"�`!uַ�'Iy2>6�-{"��P����^�N9<wLjh4�M��s�U�"�_��V:G*au�� �*�D\P<O�0cՌ�x_�dо⧭(U�b�w~[�s
���X%�z �齱��H���H�_ׅñ��M!t�yt�ꎽ4�3Bgw�eJ�I+E��,8�p!{�l{�{:���d����@�Nq�s��GG�����u��~�C�=�m�˲�!���L�ǐ>�;��B�NK��ٗ4]c�-$]��א5��,&���ˈ�O�����ޖ�}A[_����%�WW��1c�|��`��W��&T��[ҽ߻=�����}�J')s�<E������K�-�Ejj嚼�Jc�lw�J�߿�����u����&^����5���g�0w�GS�U�;�x��<\�2��
:�����Cc�����f�����Ph^�?c���=/Ӈ�E�A5dZ	<3we��]��t)�!5��r|�[�� 
�_t���.^Ä�V2����j�^+u����O���~Q��I�V�j�g�7|)�;<,���?jNr�b5�^���$����9���d��BU�o��ҋ��dC*<�z)�{�g��H�i ���֍[��
�H�1��U�]܈���l ��CP�6O�-M�[���]�����!�,�c�����A&]CX�vh��_mD�'�f3?�A!��"��T�nN?��V���N�K���He]ψR	������2����Pͨ�$�i	ı�Boy�Q��~`�pA��s�p&|Ȉ"�gHm�O����B٭
�����`ĘZ0 ��VGR��\��>��"�߳�H���g���{��=Lf��'�J���-�����<�@�����2�Ր��뙇}�n�Ή�=��̓�8՜C"�����
�	[	[�{>���"�w�-2���5l��J��|�Ps�g��@���*�֩ss����Ϙ���U��+8N}�{^U%Q�yq>H���xM�r��&��rB ��l���=��5���(N��72�o�3��ٙ�#R~�)w��
���������ζaQ���k�s�E�"��D��`�_��"��(�M����U.,���'� ̀b�������{y�6��i�'���aMz��d$}�FRWv��(U�s��2�	�2=�� O;k~N��.v/HG�Ũ�hN��5S�
�Y@t�AV7� ���lU�;�!�k������<-��E)�� �iƘ���y6�͟o�H���	�nQx�&�wҒ���Rɿ�ɇ]~Z�a%�Fd�k�
sO��<�������=.�kl�;yK=۠��L��}9'��X*�8�T[�:���Ǩv�'^5ə�:�P��D�ǈ�o˖����ʸ����zJz���kͩ�˴�}ח�n����`�>_KIpZ[��9#"��J�F��ee�txϬ���*}#B/�[��L�SjI������L��������-��;���f&$
<�L<����������@X��BR�Ա{��64+��w~B�c���ԓnla�]���1�-�`g�Q�D�)tsJ6R�x3�%f9<�&��6�'�V4���� P�J��>��'r_��)�K�^�w�V����Cܠ��*#�ޔ������A�٧���Ʋ�1�y.����<�3>��Ԉ@U�Ǫ^e�wcZt!�^)���̆s3�����(�|WT�L�~0��$�'�P��13',kTy3��͡UKqe��՜��X����}ʱMp�qsCe�R���s���7���.}6�$s����y�t���(�Ɛ��P*��N�����gF+��Mޛ��ۑ�d#�%����h���2%�4����I�2�>d	����7"�	trk$���ኧy�"�����*9�3��u��H`�6R�MG�c^���܁pE��+W��P1VV[�E�a���}�
��Am�&_Y$�5�2��iE[Nj� *D�/}Cބ�7Jc,N���<�����M2����>�R�Vm�C���]��~�0{\C��x�����s��bR��L�}�G]~�
Oe���jjH{y��x�^� U������N�}�<
n���p�����
e��{qG��\ǩ��3f��#D��"����72C@m��Q]� =^:>�)�L�d��"z9��@|I�b��Ǡ�rH�e�"w��!�l;ZT��[c�ڷ�<Gv�4m�@����DY���i�ЬtG��]���΀��џ#k�,��Bl�r�J@�eWg��G���I�Xq�-^����w��&�����w�P��e� �w�	/+�z߇}Z��J驫�-p���g��U<}�Ue�_s�='(4%F���=�4�����ӄ�3��s�,�3��n����7�B`�D$�n�%�\���L�(�1wV
�_@�~]�#2P7?���O�-�6|��ֿ������p�[�uUU�?]]9	@Y?[9a45guv�"X�/C-'<wT�B�Aa={j�IOs����Pןb EF��j.X����}�I�X�5.���\�GQ����R��v�x��8���Z`4-cQc�ճll��ڨu��x �
9W41'[<����f���U@I�`S�IQ&���Ԓ��&��=���]��|d"�T�Xm��W��Q^�p~�����E/�^�=����9;�����y���2�Z��;���)p0��Q�nK�g���yga�7�6~�ԫN�}-999pj��#r�����q�d��G����#�۷�}�� ��p���O��jLN-3�,b����9j��jz+�v��1oe&M�`�o�e�'��*�N�]O���[��p��%ٙ��3��^���	�R�zn����BH='��~�@���~��ĩ��'�����t��e���^��D�K=d�S��>���,�5�aH�M����NE��`_4�e��L�P�4�Ȗ��k��&G_��Nņ�oH��\�=�&�I���Eڄ}�ѷፃ����8d"�C����{��e�V�Rt��ON�xi{�D*��P7�
1���9�� 3���K�P��ܝ穰 �
Y-?���3x�Ѻ�����7�IT@=�O��;�;�A*�KxÙ�}\�js���9�r�[���L�3���G����2}��E��������?Ɣ���k|��%�-�O�ZU�bp�8���k�I�yq�� =�-�����k����t�rX���-�yJ�2��l�C!H� ʕ���6�Tt
[���=�S9�S��i��>���T����o�e,߇�ډfkqe�BD���3��@)K8T(=\�a�>���a���c=��u�̞�{�_��`���H�2��o�ϵ��dr!_h(�7\%����_��r6�EMW��F�'��9�';�Y_Њ��ٶ:f4�t�֠T_#���t+�f�{�������/5&����,B������j�Ơ2of��d�Bj�,�fn�7�n��1�\��{k�~B�NNŮ�([R�4�s�Kgo5,ԯ�}��-Ɓ��#4�/�7��E)�fvvz���
�T�A��;Uа�]�_���W��\��^Byyy�ؑ��Y��S$��q�������zF�����+ԕ��rP�X�j�k���`~��<�I��_��\��iK,e�����0LXa�]�[$�D��\��h����}ؾ�Ƹ0�)!w?��6�%u~���F��?����W,�����j1�\^�q<�vp�aJ�iAaN��ѪYUR����`�ʻ���5]��!�s4	6o��g�"P��AB�tN h��h�4�FQ���0�|0�3�p��ƣ�0{�~_������U�i��R}(�ޏ1�n9��&q�ı�����K]X�sR�C^��!1�WLb���A	����F��S�Y{0Qi{��Jg	:Z�U��oy��ԉ�ޑ(b�"�%��������>��k�4���l��#c�d��r�V���.���y+����]}�_h�n�KE'�A=H}���<l���%�S�y�ա�&�K�"�J7�kn��y�ȥPŌ�t���o��_6��h���Y S�3��@��`�0�U���Q,�E ���O���x��g�Sl��l""%ޯZ���4������CP��L_w���BZ�.�Z����<ꡟ��[#!�W3�Ս�u X�dx�����a�{��H3��N�PIm��,:�N�X� /�o�_�ξ��hw�Q_"X�-odz�ש���0 �ga�a��<�t�,�\J��Zo��񵪈��-�eNk�$����ZbB��f��K�����d��1�w��C�u��_@Ҩ�	���)T�lEc�d$g��%c���<�m	Wx��.�����O5���U7�|xb'��<��y���0ʤ��#E�z	��װ4���rS'��s�4�Wݧ"�\��D&z��#�V���E�$߇�%��ME}�A���x�� �Ș�vXa��7��p�?*�� �z��X7���e��r�8�[��Ed�Pqb	����I'y��+*�K�N}N�5HOn2�<��|��}��0����C�$&Y����,l(Q��y*f�Ն�P��̟v���WҖO�� R�}���.:�l�%�ܶP��������]4z�|UIEu��?����ΝHYh�C��P��O\&�;V')xv��%�f{��m���M�t�H���,Ȭ�J�%�o'X���#��ny<�%\f�ƌ��q` �[;ڐ^��b�7
������YV`�]�@1pl���޸��m�Zj�e�P���>u��ct��JR�ƣ30��>H��-�2w����h�k7Ϩ�r_,�}��@9��[Af4
�7�D��������7������E�t%EO�T��Ͻ[�a�8��dOGݥB��<��?�f�/�&$͒ݷB!f�����+~Z���*S���?yE�3����W-
ص(�1��Pz�����_ !x�����{[��p�]T������iV�-m#��]j�Ӌg7��T�y.�g���'��!y��E|��N���� ��jE���k��ę`Q����q�,��M��v3���w�_�]��C����}z�{��]�d(w�܃�݃����V�~�ﰈ��u^й�u��0$r�}���o���[:%�`u�~�������Y4�S�
b�m�����8kp����x�����^l�6��^{
\��=j�¯��L��/���rw�>fP��㒺����"xb����գS�آT�KV���=U�ˮ��U�5�3��T����(Ӓ^�t�ъ�(�ɲ���%�4�_?�mZ0�$������$�O5���U�]E�����eM�6����Y*x=T�b�ra\u�v���.K�������*`%M3URP�~��b��������&rW�V�����e8a��T�斷D+�I�/�2x��un���$��v�ZF�^��r]����2WTǲ�@����7��zq}���H�01�,�~EIII�r�j��&���ƲI���yF�Pi�~Ը�,�cy��GK.�fQ�[�n9���B��+�J��C�/�|P�خ�O �+3�ތ'��8��)C�,�� %���϶�54:��1!`��m7%�fZ��i^	}������oV�]A�9J�l�EbF���jp��$I�����G] 39���suc̿`�B_ƻ|�rKO�������0 �N��C�4b�k��3;;;;��q����՘��+�^y䵐>ʩ��XU)ݮ��_�� '�7���D�\���1 ��#�V~`)��iLJ0���m4�X3!�8K
��G�xF139���"�h� a�V��:�ڕ�m�*s�֚?�V��ݾ�?>2�@���I|�:*5|m�mT�����.Z<��k羄�<>���I��\�N&��au��(#ߊ�S��d��n�ܕ-������
��7��u�w���`<���F[i�|e�U�{��H���;|����N�x�=�&{��2�
�L����DUs�~�Pz(���=�K�_u�����o�t��I����CUF����J3�I�N@c���\]�y*ɦ*\��}d_�^��{ �-k��SkwG��C�^ޒVt�Ut�ؤ�6�*�sm���]hèW�Y�ӏZ�����`h�)�����׆g���Ӕ�4N�au�ȕ������p��ka�"ǔ��q��㖐mb��<i�78��:�E_F�Ph�Db~[?�;�N�U����ӧ#P�	�߿�џtL"*]�	�V٩�o"
�[;�m@�������"�� 5鼓���h��<l�Rt��<�}��UWP)@�7�m%x��ѕ���R0V������7¦�j!3�J��M�����G��=��@o�#�@�](�M'ݐ��tB|�Rp�Pts��q�{���r�r�xi�����@M���n�q;�۱z�}j6�����N�����o^������Z�3�M��˓[�Pް�X���*�2�q�y���511�L':�z���N�z�)�ژ��A�Lh̯�X����!חMK�!h�f2��'o�Ki���U78�wZ��!�9���x�
���I�R�O��S&#��a���5�Վ��n��^�Z���&��"�i���*��8�E�_qqqPs���`=��7V����/�� ���B��Ï���{�bf����6V!!eP��Y����jz#��Hy��p��V4���1�Sb���8Qʅon{D�ϯ�a�K��G�Uz���g���Ѐ_�i��J/w-��f2�6OT�:��Mh$����^/�5աzOQ��/t��9������Vw�q���S�D��2�7�P�����O���S*X�	�K��$罬U�h�F��u���L�a(E0o�ʦ�h��ŏ�ϼ_,���U6������Q�� ��Dn\�K�nha��]�H|M���2�tY{����!h����kY:�ae�q�'�B�����:]3�^�.���i�W@}5>��#��������[�E���㽾Y�v��9�~TQu��ZP@�|��Ʃ>�U��
o%����500�8�ĉ���[��V^-�)�*j9�X�)b99J{r�W 4��M����A���
���,G��xF#K�\?�l�^�'��EX����ʄwB}A�@�y1-=���D�,�Ím���w�Ըuf��^ ��0��ݟ���!l�6��Ч��H�x��n���,�L���_O�s-S�[(��At	�ƫ���X�&{j5l��J��t�TI���>=��j7�v`*���l�[0f�G.�%9�l-J��K�����>M�&��AM������?%EQ�`R��� f��4@��c��N��+�'퓯V�akEkK�J�����F��"v~�)� 
���n��㾻!��n-���5r/7��z ���6o�a���8��q�|�ҏ��`��P|o�y�7N��mJ�?{UÖ��^��e��|��#P����
k��#X���˕k��M� v5��S��(0�I�M�z��%i���S��D2�W������-�����Y���N��ʂ�(ɚhM���S���U��N�:rE��r�O�����ȾIy-Ol�LJ����s�Oc�\7�^s�_P��A�W5&OM��r�ܠ�T�z9���g�w��hV~�Ȧ
�9���r��)"�oX\�r
O$s�Ûۘ�NfF�%*QWG)JQm&�t�CoI���!Z)�f���6K}��Է�G&ZL�w}�8㓒 JI�ɓ@��n���/(�O�r1R�s5�76�|��n��x��]d�����G��A�k�P�S�������
c�� N��H�A�{�34��_Zoj%����N[�Ua4+5CD7O�d+��9
�� BO�r�����l����g��?�P��s��o�	g��y���j�M=}m�^)fLk�F��r�!�r4]2��u�[��և�y���j�L�}�����v�EL���l7� �
��ff�>��59�c]�P�Ivc�
b�l��/�Uf�x_J�T���l��J_���9��v�>v�gJ�v�L������$Ұ����"=��r�v�$l�����g"}X�؝��g����1�������K@�Խ�$��eM�gM���Z �&���I���B+��L\m3TC���y�z;8�P#��_�-��Th�Kզ��^
�GQ3A~,����:��9�jA��ż����}[��,a��e������O��M	�9!p���|7V�r����J.����r�����U��S�r��Y����x:�t�sfQ�b��#��h2�������H��54��o��*��4d�= }�u��
[��{NZ�_��(ȘZ����m�<[���׶џ�
�-.ag��;�Q�1��G�d-�1F��(�_�l��X�Qv�%���;h�����Fd��4+*0��B^*��mՏ�T���3T�ZP��R<uN�K ��,)}�iR�0�i����J��[�y���5�����;�/���	��_����ݝ��(<<}�}���F�+G�;�c����� u���|������y+��X���r9��Nh�j�g`8�MnCrpxd�D8��j ��=�XI���3�����^ܗ�ĕT�g�tm �pj\w�YL��!hȦ��[�{Iy����*��(g�|	.!?�z8��;��؉c��$��?�������A�//�I�v���rs����.O�$�l����4cw��2��8qjL?�2��L�ݹ�ǍLl����|�'��$���e"<[�Q��Z|-/+-�%�1�(��m�$�kY�k����OEh�ym��0�B���R����N=�뉶�.��uƅi���p�9'�?��}oM��>q�fR������~|�EG8�r�ߦ�cY��t����Ih�}&��jP]��2��^_.��j>��K��6�+8~���q�(��uEf�a`)5r�<��QW�Cڒ �cTqq�� �FS��/vޓ�m��p�z� ����P#Ҫ[7"��w?�Xx��u�JA���h�t�)#6�
H���3�K��u�R����a�m�����D�U��ՙ�p �7>8��\��tK{J/a��4���_E�dP��=4rZ�Zt�1}����q��>� �!��!O�?#�o��O�V���0�G��e��l�yÂ��f�^�m���RFފ��ips)usD:h�+��T?�L��T\ou��ON���l��h�� }x�P݊��a|[���Fܬ�ɼ���J��y�����y&Dʖ}�2aS(釀-��M)�����xJ���ֹM�H���?Gh�7�c��O��"-�G��e�����=<�t!�p|LT|]A��۽�C�j�o��,�A��D��ā�-���@��>�э�'�V�(��=��#���R��W��m�K�x�j���~��l_�
�N깺s�睠]�`��l��>͢KG�+�_��m����.Ĩ�����{����)=mj�a��OB&����`&�;f֝��� o�NQ3B�c�|���[ ���	�����pO8�x���=;�$u������N� k����4�m�n/G�,��e��Up��Y�T��S�[_L�~���Sj���6�$�z�P����Dl0ەw����V�� ���h��Q"A��LPj?�4��?�4�F���3��c<�#�ſȀf� Vە%�"(~���2���nd[^f�P_�&�u)�jxA�],)W%�đ�d~���nM���NN��WM�=}���0�Dr
#oiݻ��C�Wj�\)��?�������6I�&�k��d��D���Ԅ����j6c��}�����o���!j��/�.1:�{�'X��1�<��3jC���ݔ��uErN=��r�[�ˡ�����Ę�5*Q�k@������O���*GBd3y��˲�>�΄��q��cPe*�]���0�-Ķ�P��[^���t��{f����^���m߭�KJ�d�.�+e���h]p0�5�({꣈V�ʓx�r�X�"Ů���K����hn�ո�vi+�vL�X�.K����'�d)��:�ޫ0�������?9dS��ɮ�tdD�讄�d���SVG����EQ�l99Ƒ��BV��d�C���]o���{<�'�^�k<���N��2�g~ӯh�qiNx��R�g$��>��$��37�#XMuIa�M}�Y�^mB���Yy�~K�ːӔ��?� x��,Z���{�XjA3u��ro���{���F�T��(�<�m��}���i+?���:����n���k�v���B�����0���o�,��B��`�=-�;v��ș�e��m^���-�Њ߶�z���jAȟ1���c�OoN��� �i�q3_e�0q��L���ֲ:��%���������},@�z���%|�gpp�kx8k�+A�4Aڠ1Y'Nݼ�����=%<'*T(44t�m��Z�s�q&��	v�ƺ��p7JN��9 k�Ue%{(��� �t�Q=R�6������q�F���� ەo�ׯ��jjj�_}&�8��օ͗A���33-w9��'vT�~5U�q+mK�':��G;h��J��=��m��)^++ny^��M�����KZO0��s-n�ЃNyq�"K���_g��F
VPWW��q� ��03Lޓ��u�EԚ�u.W�Z
j��OS�Z�0�jLLX=nk}=8��u����2��������wɑ'^�|��e����=�%txE'�<�%�5���S5�����Ur���nCӱ�A~▽VXQ5q�0��sm'"x��˃�z�+����H��X�nl<���}a�޳ۥ��y��l|Rj��Kv���k�ќ�S��a~N��-}��:\37�X�#�)?=n�ٮ��p�F��+}�J��7&�i�􅋕Y�Ž�ѐzd�z%� 6��U��Ǧ��iȧ?�7���I���Sտ�C�9jUA˼{��j�%�Ec`_?u����@�7��"�h�!����'� ��$rL����#ZI�^����JW�N�a��4>8��W��A��'i���NL0ϖ����b�j97�e�b�L�����|о���(]"��S���p~��ku�]%%Ogg��С��̱�Dm��Pm7���{��W<�OM1��Jc^��$���ʲ�'��g����s�R�!����!�&�G��j^I��O���b*��ia��ӳ�f�%v_Yʟ��Y�Y�q��u��ͼ�b��]O�ۭ.s�6�555��v�h��\/��EEY
�m�`}G��'Y����72��yE��8m����=&��x� o.pM����P��ɦ��Bp:o���(]����w?@II��zr�I��tD���/)��+�}���}*�49Z���]���(��w������lV�`�A#%ޯx�����UE��N����Ӑv�=c��J���H��+�����D�Qć�⯛����C�I���J�x�z���>�V=X�#cxK��XS�
��3��RN��`���NE�U>�F�9�l�)֎%���Byu��*PVl��ȕϚ�z�h�c������'%����	�F�`?3���e�p�c���5�ϲ�z�x��2Tߨ(�>��������+?���k��S�E?Qǈ�V81���!9��z��v����z����ыd�2)j넄��L�g��h��
5��i"�o*d]b�N�!G�Dd_��x�	Ý�;����$m׭�	{�VZ^~�2F�� �|`&�yM�N�Q.4�^%_�F�7x�x\��/}��_Y��W��b.�[n��R���]��(��瘖�h�~/�w��g�=Ŏ����?��������,��OM��H���f�)���m�Ճ�|���Cᒔ�]�����6=+.Zb�G:�F��_#��. �C����x�f��9i��9]H1	��?�������1��=�> �PȞ�*IЗ	\H��{�cm+I���	)��'骺��UUn>�~qXwyk������������Fp�]�	i�r�Y��-�Я��x͟�������t�dW��qT�� �ɷ[�J+** ��~TĒ��K��7��D��Ԡ`kk�ãzb���`SsklD�[�34n��l���O���O=��l>��q����g+mi�d�jƏ
�>��u#�~���'�˴���@�ͪRc�=Z���������_�ml��,wz�E�`'C�&o�A��p3�f!�h����?`4^����'���iR�Q$ԭ����&v�+^ԫI�颉�Q�0r����>炶�	y����a��΃lD�)� �2�&�o1��2Ÿc�ֿښ}��(Q ,3��ۛi-�# G���)����Q�V���M��Y��Rl��v�==�Ū�K�A{=���0�*-t:���,U\.�H���a߉�J���"&/�Y�u8ꘙ`2%�?;��F۵�X(�,��t���QV\L�� ��W3h;��í��W��`�w�$�u����@Z^~S��9Y6��Ca������+L���f_�L�W�c{V���ܳ��&��

�֏����&�ߓ�X�������'�/����T�ѻ�G��f[��.'�/6 a����M���i��Vud�}a�;��&ݣ��зdt��|3��	�am,�%�P�=4����vS�o���ʰ��j���85a�@_��֦�&��m�ǩ����X��[iVb^�Q��
���hN@r\i��d�5�_�S������C3�����i}]+56�B��z/�k�]фl����OV�:��\5a���ړ��l��0��0�B�0�_JyM�@�qz%=�JF����vpx1��E��s�F�qvmD&P(7$��R�	h==K��~S�Ԫ�m�f� ���J�9,�����_���S���vW�R��׫5�$e�t���񲲱au2���?X���$�<_����h7^O96�42RN�iS� �D��3D�K#n�f��0�[����ֱ����wA����y��>�'����#0��$�������r<q*�>�2�GX�M�/n�>0O=-gQ�}�ڵk���Wն	@�$��Ss��2^��f�[bp�*5�F6vr.���e��<�u�H֒	���f����e��Q����TK�09�<7�^x���ԯ�ȫ���	�_����6~�Hz+���A`;6":�7��8��e�����YZ���[֨y�r�~��o/a��U(�O�y��7�ۏr#oHE��Q��6喅97A���k�N�@<��i���8b�_�����F���>" S�K�G����/��<�8s�!$�Ԉ��#2�~���;��ȾT(��i���+�#�0�T�2;q+`�����ܜh��r|��4�?؀%b��$tv�$&�͘���uԛ���ܸ}�v��[b��|&,
���Q�|��sk�7����2�?�йq����ʕ��6"a8fO���E��.���F(6���j(;�f�$n���aᎵ]yU�b�L}�-��,�Аkn����"��+�.��*��u���3�U��?�ؚ�32p�[��r���b>��R&�<Y�P��G��[�O#r��J7�^�3�pJ�/Mоw��%EE�����͟{~�2͟���6X�+��)��nl�Xm��E����j��K�h�dLFj%j�4��������13ށ�`��`����"%����҇;&�Px�_��V�?x-����W�� =rn����NQ�A�}	���aGBr97ʁئ�A_Y��iKȐTza����Ċ{�l k�*nO)�����a8nLHz��-�]^�vw�F�tPj�r��۰I> Zzꑍ����!lp�V9��*�؍� ) ��z頋�N=>�U�8]t�od�sq`�ݲ��7u�����;_k^	l�,��˃�tuoFV; q@��p7Z�����l>��>���0^�U1 }v�W[�s"Ƿo����w�`�����f���l��ӣ��1��	nA;V�nx�R5x7�������ܬ2ʽ �5�Ǽj��dۻ�a+�U/�C���Wf�Kʦ��I��N�e�=Ы�֏�.��>'}�Nl�A q����θ��&�B�w_�	W�"ޡ,&���|� �bs���gI�߸0P��R���&V&�c__@Ӡ�+9p���0��+�?N��S�������2C�ih�ӑ#l�7�n����c@������� 2��v1��Er�S"��%�
h"3��5��y纴��L(�O�ssHC�w���2�?�;dWZ��ðy�d`���%4D/��#�3(�)�%��M(]@U��]/����X�xAB[�kVV?�5�Q���b����
�
ac���4��I��Nzaha暎A��IX˱��}b�6�z��qn�0��<7��4.��H��0�}D=��R��7�
�^ �U,�=�m�m���������K���OT�Q[�k{�5�qP^Y���-u�[.�F������[in��Y6q�zdfhtD�����SH�_g�7�,�gJI�/^�|5&�`�����Lk{���_�0�2i��eI�vl���tU�GIc~�`O�Y�����p6@E�C�����C�S�]p����(`v�H���jLM���N�iY":��s���3a��i��_=�*�7\\��Ҷ���,��#������I�9Ɩw��l�VSgN���?�z�87D9�#]#�g3�e�+��B5���^l����n�_��X��f&���ي�o"N�e��0�����8$��}��y�Y�d��=,��e���vb̍�0�S^K`eR�\�~o���F��9�g�B�#�pz��<񔀂"P���~j19-�P74�n$�^�\�s�����--iZV�AbY-�4~3b7.z(s���ׁ:���+�R3`'X�ĚFG_������/;��4��ɖV��Y�6��ne�V%8��C���[W��ސ�X��T�&gg�� M��TVT|ו#P�"�N�ƕs>�%��Y L+)YH-���T�i��X�\��ȥqeA.b��n��E&nE�1�K�[�Xoؤy�X��jKQx1��NSS+(��ƹ��v��S}��n����RPRB/��J���t^��x�����Ye��Ҕ=}�^��ުl�(��NVfwK���@�z$.T(Џ�a���>(���uh1'�2_tm��P?������/<3��}�Fh@}ϕ�������Ձ=��:;��OҊ���I�
3g�1UW����8K�89����]���L\����|Lo}8(&�}c Ia��*.����n��u�R����vjMxhh:�QA�u�����{�P!&��5�vևրQ=|������xs �� 5��k�}O����Tu����S����ӫ��t	� w�t�t�[5��{3�ޚjSc�P��E�2��΍)��f�Wi�!�ӏS�l�cx����_�ul��O����?[ݍڞ�db���T�G�G���Ɪ��w��vWߍ��H�s{e�s�$drf�z`��u^I���j�;��bb���������7��45e�Z;#(���K�f�����{�c��#�/��ޮ�P���%��ƲR���V�(�����y3֜��s��H�Ϯ�n�d�92�_�~��s�'Q��G�[g��ԋio��{j����˳��:1�̙�-��d�v)���f�-�WJ
����:iђ`����tǽ�ິ�Sd��U�����2H��M���1P��Ir�SiZ���r��r���ai��#�j{%���Q�t���Co�H<}Z��6<��vW���,*�>x��2!�������C�+���;�m�˹���6�B�߮q�m�j^+'�g[����/�z��@N,M3�QO�Ac��>/"4�p\��p���"���~0�c�W��cg~�LVĆn��\�^��Z��9���ڍ�g�Oas|
����Yp<�A�9>Å�&�{�c�gN��h�~p3�����+=�a���̓;����a4����z�7Htwt!{����{�]n��F������kc��Z��c^ ��\ �1lm��C��\�	��k�=��`i��~*�T��5�Lpx�F��V��5J�p��\��\8��=8�}DP��(XN"}�:��6������Lq�e���r)Z�z�}�=u!΁���J�|~��ծ�����F_d���w�P�2kl@�v�YE�N�E�Lp:�ʸ��6�x�?5׻]���U�+�~[��&�X|�i��JoyL�p����{�O\�(��XD����1���?��uߘ���.���%���KHye��}]��xYi�(����NǶ�R/�nd�|@3� 3�z�M����J�Z��9���H�0- )��S��4���O+9P<Ի��À:gA�O>v�����������L6+~j������'w!�c��W��C�7������\�N��0ڍl"�#O�f�CY����a���d����~T�q�vy^]�m*����Nݵ�"�jS�T�LM�lO�SeUϬ�/>M��ٺ�.��׵�m�������u�YW`���!��f�BBDGL��0�^���)'���k
��<!ٞ����D|E���u�&�|�%f)h#���[=��,���!%�e�`�{�Km��0��u�3g1�25f�1>���h�ދɛ��y�Wd���%ج;6�q/�:y�	�N������֝�(�c��{Fx]��x��N�lI�<���,�YZX!��n޻����U���cS��M������{*P����N	����v���(�a�W?t��9�Q��,���W�������9�GZ�m�KD�M���!�t�lRg�݆��<%Eˊ禧
��wK��/T�v��i���z�*�n/u�,�����;�Ζ���>�hi2B�_
�J�[���Қ���?\)�s�,�u��![>t�ݘ�.�1P�E7��Q���A4�לk��7B���<H�%w���A�-Iy��H L.��:�\�M,�l��)b�;nm�jH�wePÎb �Z�Y��@����ҳkՍ��������:o�]�M��e.��Y��	�B��5
7���'�m$9?��~]^&<?ϢQQ�J����Klu��8ۭ�xD�.A?�c�{�@��WF$7���m��Ŀ=��g�������rU0fĔ׵��*����8r����yv�gU���u�'����V	�a��\.�do�����<�V�|!$&�U&\��qA�W�^���忱x���!�����΋��a_U������v�'�\<1sJ}8|-'��Q��ߐ�2�))lA����v�_'E#kj�SQ�/�Gb?�x�4s�w�
R�eqrph�%��s�j��g�_Oˡ��+����7�x���Q����#���URY����C����{��ث1�X�-! :�n���SU�V����u^�Q�,LCj��M6�G[B�j������ݏ��h�x4������n��R.]�q4f��׍��3�,���fM7%rX�J��s%&�;��]��H��+)a�]�a�Ar��ʏd�zZ�f0;LEM���=�c����� +�Ia[��d�O�����<�4�&r�ˆ��x��Z{���$W��
��Vv��B��ͻ/9c�ٻ�����#�'i�8ɫ~�����JOǙj��E�'�����řN��N�`�>��ؑJ�b:�[��;0�Uֆ�84S!T��u�XVTR����k},*p+��S��s����n��Q[q��\+'Rj��@���>����g,�J�%�
�Ŝ35�t=M���,�e"M@Z��;�+hik$�l����l|։{|�}��`�o�joK�Ӯ>�wX9K����QN�$B���ѓ�a������[A?��b���2)���:�C^�%��	ti��W)�m4�J111^��GX￧J�Ȳv��>�T��AWW� 6J655a���|������z�nd�M?�R\�	�����?t�N��Y,..�y�pa�
�����5'�����3��� >o�)uzĞ����E��~���;�βݗ��Č܋�q��LfG*�>�	�����w������&-��%�,��P�?p����ń�W��K몧"Y��g{y��Ps8쐙KLa�7CCM�@ch�+�o��-lSB�u��F��m���w��YEf��K����I��?��\��k��_���۞&���/��������;n]��D��Ǽ��3��ǂ%�<��&@W@�U۱v�kR� 뎮�������#�H�� ��aq�Px��X,��' ��͏fCa���G��B�3��~�e��&�����.�w�p�W�a�XE��}'B��'�p΅��F�W<�ǣ��u�	��Ӵ,E�T�IK�|隋��չo6����GHK�r4�P_Nq��RMC��~`���}�����sU���fl�:��7���ފ#�+��N�
tH���C��|�B�GOlWW�ng�
> ����Ü���>�j��#�HDw)��k�FK���1�|å_1����iPc$%r��Ng��+�r�<��F">Kv&�E�$BS���jv<���N�	`A��-�kE�Va��b�[2�u��Qx��/�ѩmv����I?]���ƤB�,b/�\�bJ<r^Q�(������.��Gi����4������t�0�2]ӵ[�����6��n��������s��?3��!-�i�G�Q�3�D�۬|�7����0���Mi�[�Iy<�,�S$�O�F���	�9���LWV�d�-��[ ��GOZ`��w�4)�y�\7EHk%m�2;�=�ug}RZs䯳}+�程�
��C�7H�jl�J����X�'�Ѻ4'�LN�(�ܯC��/,77~��E#5D�~2����.�b��!�t�f��F	TUlJ�*��Sb�ώ���f�m�i�A�КNX�U�9���'�Ze�}�/e�BM�u�[�d�dj.wG�MԾ2��>/V�J8�K�������CZ�^[��*\$�#���3�ϩ\j��_)N���ש������WYe�8����k��Z�����NZ��V�������	I��6��v�L�]�C�v���S#��7���8�`x{[�;n� ��>�� 73c⦟�g'��Θ����X���S uY:\�&���iݫ����J���!��[���S����џ�_�u�����Ɗ��`Z���D8��	���1�[���ڽ�ne��0ioY(����.+�t��Sct��[���}ԅ�V��qa�X��{Vw��oUX�8�bX|�r�e.����y���n?M8|������V[��=�d,�ޯ+@��?1�,�s4M�A/��9s�4#���WEA!ܾU�A�r|����:����/�	{dʽ	�8���:��)�*�*��g�SS$�{@�c2=h���h�|���VR�B�0?���ز���wa����7>��<�.�6';"����a�\�m�n���OL:b6�0���lJ���5�����ޞqįD��6K�/l&D��)����:��0��~G�4���|t��m�w�g�.�B�;h�  96M�S4���cy�1��L���a��GG��CI8t�����FM�r:@9����wV�p����'�لL3�B��lӂ�5��I�Y^|���� �Č)�f�u�ߟ�̬�;���%+���)����9}�wy����0�`�9�9��F:�K5��zIfKb<Xq��H�٘���Y���q$�m�+�e�?9�Z̟�9�PB;k&��r<�CĆ��Ѝ��[�&�2��.�Z���;��`;�sO���7]~ͬ=�[X9Zמ9޺�(���)(`b�ګ�~�KryUPקE��!���1��I	��I����d�#�v�H�ॴ���"\��q�� *~=xS�:tb>�ku7�M���D�u��?c��[������>��A�1mZ�X~�-��5�Wt��8Q0�����ҷ��'�����?�H$)5_k�on(3��:�Ǩ�!��b�jo�-�3��u|~vl���mf��X�6���o�f��d��S�Ҟ9������l�Gi��oi� ����an�+j@Q���iH��zV]~�EN��B�Oݺ����cz�H�@��I�O,,K+x�{��"��ne	�����6�*8�+^ـ�S+9��$�ZgA�3�����J�.VR�v��9�.�R_R���R�A�uj��D��>F�TW7?���q%��o8e�1��}�G}e%:� <B���y�L`n������~�Q$�Uۇ�w�P@�Ը:ܩ�����(����J����aFc�!9Po[S�p���Bܖ�4ŕ{�1!/�+L�����Ջ�:q���V�T��&��&��g��U���ׄ����������g�u#S��*�@7)[�݀�~f�ObE��(��h��y;}4П��+��o�3s)6GA��������̄)�6�o�5ٞMVJ�\���(��)C-�:�U0T�����C��ּ{I⽫�_��4�jeE4�]��լT����?Q��	�����,�A,��K��v��1�$w�mEb��I,N'������ �K�"�{n�(7)�6�˃�z�LW�� ���&�_�đI)�o�M^?���O�%y���G���7���H׻)y�EIl�^���DM$Em�"��F��-2�n.��C{��&
>�~�b+od�*n-����;"H}���ov����g�Y�o&�y6�����q^��]F�U���w����V�1-A]�����S�+��y�xQ$�o@P jȼ����Q%���u�s�?]K?�t���Wc���w��[en7+��I�_�����R�V^!�쥙~/��4��&�t�:��j����IT��FEEř�t�}��QԷ�R���"{A�j=���-.IJ������1�Xh���Ť�E�1��ts8��5B`Y��g��k�x��6����y�����a��ȿPUP~G���n, ����y�� �"���8����qY��4]��P�����1�P6+��;��wZ+�O0�����"�z������;�F	���Z~E��!4�2�� ���*���T���FB%{a���ȣ���=DE�V��K�W_�k��_�mhOt�n���Uٴ���:��%��q%����@A�UnУ�
J�LX��K(�p# ���S�b�����Yϓ,���f�R��֊�W�n��:�/ũ�dBW~����	��Xz����.C���g��=p�(1Ff�f^�ҷо�/3k�AB�md ��2�E�Qи:�1��)��f����P�����\B=<�t��D�y�m��D�ʐMh���~�]�"�#���X�_�ޙ�E��N�ܮ��8��K�,.�`�%y)�25��|��e2GM�H�mB�c�=���Ր��(�f?M�<�s=���\���aQ�[����4�����Tf2&��<f)�7U���bl��4Ѝ�����f%�s㦦AȺ�P��_�M��d�߻����fe�C �y�y�%3�阇E�ܹ��;^ vOW�n�ΝD�MŠ�y��ʈ���� ���;fD=ۺ��W�OL����6x��X����ĝ�]�=���s��R�9K�/t���B�����:5|��:,_'=���Wt�ǭo;m�CN*~�	��3��F��T<�$�gӦ�Zs�ܫƙ�r٭4������t�F�jc�#Il?�t��@�2	�O��������\8ﴮ��焯��Z |��B�$-���1*�hE�A��W#8t3��3*�BV��9�ʰ���R?W���u�I����.~�3E/t�z��m�sj����!��Ԩyq�;h�'z�� *���a�����!��~Խ�67p؋�K��������.g�{�i���;�_ɱl�
^�e�ZS�4}%���dO=2� ��~LV���V~����5
�*V��4����=�&Dl�Ww8� <Q��$NͯP]���n�>��+`�>Jz�0/;�c�Fi�=ˉ�|�:hS�k8�R퓝jU0��l�J7��j���{�x�z��� 4ݜ�z���J9�s���*�����~�.V��������!)��A�1�O)t����Y���E���L�g4c��`�g�!��Ѣ��gZ�+-��6�d2�ئP&�W���ș�R̬R�@�r7؆9eĺ�	�M&����8 t�nj�
�0K	~ڦS�ș�ӧV�� �֟�ӾMIk��}���Y(�^��G�����Kn�X6~U �o�`�V�0�R�P;�k�A�<"h-��ͫm"ٴnJ���J\/����"T"�^�&���SV���M�z��Ȳ�&љJ&�Ն� g��B80���׶Wt1�G�g�^іm�AH����ٖ�u,T`�:7J�̖8&P�K�6~��*�;{c��NP`YSǯ*}�es�	Š��Y�cA�$����9��=*��J�����O`����~Z?=�j	�-έ���F���� +�J����mm�Y��
z�gP�8��KD�p����K�di :��)�_@�3��t���g��G��_K�S��R�]S��{<��&K9��ݐE��N����4p;��xb�21��Rڐ�6�W�U���ՠ��#�3R��0\���G��-q�B�1�[&�����*İ8 ��6(�|�a������1� �N,Z��ǹ�Z�-�S��=! _�w��q���V%��O�9�
��}�p�u������&��yqhP'�N�|c'f�4�D��������#G'�_k��D��cP���; ��ԑ��0�ʕ����rm/�Y(��oefV@=�zC�.p:To�Sf'�$��{�T�P橺���V�6�D�����xF�����H �Ǚ�4j@���ȫ�l0�����PasLI\
�`eflv����<k����_
r�0�艀44�˄k�>.Ëߟ�?��dҝ� %�j�i	���NZ����w��u��/w*��a�����g�݃��>��������/�0K�~�Y�Qk�^:�n�_\3G���XS ?�$Ǘ�2�Җ����ʹ��DGr�������?r�ey-:w��Ma���q�[�_[���ɑ�^~W�,�ѻH�1;�}`@s�m���p�� �-m�t(��\?��;�에�7���Q���f>�	\w.��t}��J�=-�E�L�����a _�:��������c ��u�����$'�N[t���<���E���Ō���=��ro7F�,0Q}�|���A�������~��v�w�a'bC�g�G���cxi	�y��s� �8�w�� b�	�?6}Jz�*H������T���lD��=@�PF6�ȩ	lQ��C�K�j��-����p;�u���H�b�gL�&(=��G�����0��D�: ��q�@�����=��#��GI�8�_q�Ys.�7���RE��h���:���_¡�q�SS�3�;п��}�Z:7`3�����(cr�[�@�f��/�����v��G�s}�����h����r`�(&Q��ɱ�a��0�@ >~����Y[k�]��%��.��%���',�-��/������A\�'�_����A�bͯ��J	J��<}_x�ȸ؉11T�i	6��dӼ
+����
|/*��{���/�aϷ�tT�s��%uQ��CKe`��W�G��|~�}��L���=�ؕ�N����׻o�|@�@���J�i޷�v9�7�ԅ@O�tr;
T�>|N�LE|�x���_��C�,�v��M�gdPHR�&�r	��.�{��ز����y�N�+=�N��8���_�S�ܰIwݿ o]�N�+cb�_�3v�Kڧ~�/�1{�`��Y�Nr���.ՇE�eڱЍ"��a}7���B����LX����.RP+_H�f�������N��2 �.�3��a�Q^ϛ�ĩ;���㥷���O�lTr
���rf�y�:I�ΘcȄK�
�S~�����> ;@m�	(��bJQo����w:�S��U�f"7����M���=��nS�X{�Ӆ��>�"��/��<��Z�;�q�����(�wcP�,���Q�An���I�*�l �P	����J0��=|�$��d�h���ǾZs��UA$}�ц��-y�p��(U�;/z�!��@��G�ʵ��2���r!��p����;����;�*&�Lu��2���U_�z�7��A�v-��L؛�6׀~}�*�3��AJ��,Ԋ�s*��c�AuN�f�����۸P՚
jc�j�3/�ʄ���I)�`�u�t�����"f/���2�D���8 N�������j`�r���Z�t���F��g�Kb�m fRϵiJ�!̎���~�p�7|-�M��b��L.�Fj���^�6uI��Zf�[�ָX���@�^Z���<}�U�Z�˪M�@#)8݆�8k���,��Y�|GNO1V`�]M�2�Db�ૺ`}�>hx��>k�Ʊt�-IC�Gq�N�$Г�Tgi'��a���� c�I/T���/���x��6��� �٩����m�BR�>�(3	��5���$�^6���w��D�ۑ'�0�����
�pERPyL�(�D�65���/C�$�j�
0���J)����߂�E־}y�R�,�KJiٿN�d�g���y��s�-!�����^}���r��`�[�1�e/���-��7VX��0v�{u9o��?z�?���8ٵYa�ͨf���p����ӆ�l~�(gmI�<��>��;
��+P�i���a44�,���U����Z�62Pu<1�|�i��-�;�/��R�@w���4�w��9^9�M���B�2�s��
�e 7Q��Q�U)w��� pF�`�����]�Z����� &4�ŗi�l��+K�F~�{y��C�-v��y̅iMx_�k+��BF�u�<�q�w.��o�=�@�U��갾Q�W�Q�8�2��7�g}���$�.R����U�����@$O��Z=mt^u�V��/o���+x�l"լ�wI3_�[�Wԣ�/���+_5}�D��C�$����▿��Of�(�u`#n�O��9��W���g4�)��2N���{*������X�J:�����(�d;�J����'^;z�K�1�~�� �Č��	��r2�' 4�c�$q(����#�^n���%�Bhjن�>�ϸW#��"i��c��������5J�kJ�5�(y�6-�f݃�W�cb���&��G��J�m�Gu�)����V߻:�=���v�%��#��6�KhK	� �C�u��85��u���{	_���ɨ���H�^�&]W�/�-=ŧҤ[l�f�:�i�N-f��GA~q�u����7�]i��I�*�K��M~q�^#5�t�������	�y5z �@� ���t)(�c�ێ���j�J�P�����oB[d#8LׯH�⻼�8{�I���yl��2˒��%E&�o�oK��t��ޮ~X�_z�8�|�d�6�Í��PW��1\��h�۵�漦���\�)����w�_�c�"���B�va:�� �2�W���';	�~͟����
5RE�dJ�����ZK+��`41EC�%ߺ��k_���^��1�D����!�G5�͑'`hs炠3�y�+l8۱��������[�/[v<�!k��Y���T9K�k���'Ǆ�x��J�d�8I$�NU�QA؇Jd��6�:6�����(�l���}��n�W�l�JVOݫS�n�Q8L�K�&ĔA{����|A��
�>k6�VLNq���*����x�#���b@9���*����i2������<}�mF�ة����U�'I��#+{�L�P4}�+�������268�)3��:(�-!U��^]RcC1�F��lƒu�$��N��A]�������D���W������S���BMw�/1��I�I�'h$�|:鏁�����G�[������@�O��~δ �Ҫ!g� �4�Q���~F��/��E�\�'�W�),���J�2�u|�Q�j<�����͜9:L7�)U��	����5��/��}�ⰾN���UL,u#�'n�g��g�[x�o�ˇg�m:�OPq��Ԗj�DY�����ӡ���� :�����q��
�r���0���[NP`�������"~J.w���)>�~�XpHeZI%Q>�F�%����~N��f�hx��S	��a��[��|0ܦ��0�|���c�1*B�?�XJS��,�/FJ��Q.bp��$�8=���h��i�oD�σ�$U�.  �W���b�� ��FZ��O�9�=
�sʸt{A�'	fy����O�����a;�&bX�{�-��~�#({e8̃J�!�r�P6;�@���aiQƜ�FxT�����v �dw N�}a�3�6���^����
���%���tM�8�6��b$  �I�V�9 �F%X@��E3�%������]�DY��J+T������S��_Q��1l]L�e���;�
Eנ���kDFj��d�/Ϡ��@��Ρ!!�n>_���	�r��5]�H��\�b�|�̢(�0X�S�s���F$�`2����{Jk�ʁ[6��V�zH�y�=��QP�!
� ɻ*��gb�-����-}�?�DGX�oc��
��F��P�W�o�h7�m	�e,�b�k��Ą�h<%�������ʶ�<Q`���Z"/�Տg�0^�{���a�s%���l�������Q�P�"�ߛ�R�
�լm��"y9A=�@xb��
�;ٶ��#�y��,?�r���lBS��f��9J;��.�k�埰_�yf��\��4�g=s%���
,�D�ԻJ���d��m�1N��k����k������;��~"��6��l��iD�}!�qE�����S��5�����V���ب�A��%���e񺯊�YK>��N����D�����B��(�14X���Y�i6����F��s%{.3ᚏ��������0�f�+0�~���:�9����D��\�#�R�?w,�j��l�P�/l����|� cA'ЦG�{U��X�Z!&=�^���\�,�WH�Ls;9��w�Dn��sC\��LH���Bw��T��5��H�4�J���r�+x*ܬ#dl�,�S�k!���_a��O��5�S�"}���vL�	r��ï�R�������P�ǳ���"�E�{��i0�A��=��`����U�59KT+�H� ��0Uf.��#3	�����]��F���P8���/��{����%���fC�ei�}ɾ�]c�¨�-%*#�d#!	E�6#K��}_~����^��ԕ�>���k��y�i,l�E��p�h�:�Qe5��4�Ԋ?ߞ�mw*�t����mM���DYfg_���d����O�u.�J���'r������bA�A�js���� �Ӏh5�SC+���ʟ���8���Φƫi>H�@1ʽ"Q|����k,,�`�$�� *�ߒ]i�ʿ�~J���S�м3 �YF�+'�����`RE����>���H�f��B� p�;��Bo�vwQ��K-x���92w6�Q �,P��u���K��A����i�)!��C�3!�:��+��nԠ���n��ݷ�?9�-!��;43m�s�V�.V�AJ�;�"����]������'��� ���n�*��#�S�M�@��Op�Kp@�ټg���nnZ�w���/���3xV,x�fyl�-��R�����L�$P.�*s;�{s�(�s_@o�b�����&\����}ޠj	{Z׿�ê�.`��w7��{l.��ć�,C��O��c"}80�aնH�@_���xm�A���|o;$Q���r�R����'�
��N���sq8I~p�P6I��,@D����7;)�^���r��u��y��Yz����Yi�awO=D�P0}\/G稙AV��VS[����n��J���]�*KMBI��9��LJ8]���<��31��CN��N<
�+@���Dۄ�|��+��m��7+���W$s��W�5WQ^�ʹ���A��7\���Hh���f�d��^V�qm��^~ {}����T�+jmQ�<��'����� W;^�	Oɾ�u���jw�m���1�p�!�+��#���Ns��'��;z�s���������%���K'��{zz S��P�K���"�7�i��q�ҽn�8%�7A:��M�j��!�:�;��*��e!SU�	\��o�9f���)���u�c��R�#3�oF� �8������@G���-�ꑀ(M.f����3$UB%!Y�C��|Dn�	f��j˭���왯�6��a��7L�DlAy^ڿr%�\.����|?���Jc��M<%^�m�^�ؼ
 �4)�a݂�FN}N����a��f�9h+=�ҕ�(��R��|>�*S����ࣰ�\�O�{W� j!� D��������]���SBJ���,?G�܄���'�ɒ�ơ+��ӫ�n2��������"獀�����ujN��>�ۍ�X�4�.To�м��r&�M��їV��*tQ���@�e$k�2��Ea�j
P�q��y_����X�{-f0��c�����x	��ᖼ�eEM�BJg��!���֗i�� �~�$�R;���=����'?���
�>�����|�j�Z��.Q�D��R}Z�͖'?��>�,e��&
�+˛v���)n]�]-�����D$'z���y?<_x��C�X��]HyEj�2�,�`6�7��mM�����d��
�e�4���ܦG�o
�=x��r�	��TN������#��@=�r]L�>/���X��隇���,�QdzUϸ��e��@ ���������u!��h]�0���"��	J�zru�^:)J����|�f4�g���ɺ��W��,`�⽻Pc��NA=1��ح�����'g�O�@r�T��?���F�?�~�@�b�=�T�6DKL~�Y������5��� �F�ų'�e���ϟ!F�=�T���P�:���{"��|̃i>j�Rb��m�}Qjʗͫ�P �
�J ��v0��2r���;��r[bZ�@�e��ua�.�ToQ���D�l�Őc0t����jPҋ���&�d���!�H9he/��`f�s��>�8�/�,��?m�FhO��D	��v�����dʔyv�/�X��La��k���_K$�RV��x�IYEW_u���.[Z���Q�3^R�$��]=�=�҃`?���̾��3G���P�;/��f�(fiN�?SW�%N �j�����^�d_�5F�1�Rs G���S����9>����,���y<S�QKՋ��yM�FMsy�;'��#]3�7;{�u]�:��3_H��'%�k�\�t9�����RF {Ӹ#P. �xx�n��Y�e�
�~�,F:"LQJtCG���������ј��D!i�ٞ���:�&�܉.}!�w�>�>���.cn���ׁK����_O�l��o7���X*���8��%���mW��,� s�.��<�n\r%Jϯ�"�hJBQY�l�B
���t���)8V���f���ḻ���{���C{UlMG�M�i���}G�y�)��0�a1U�Y+�ޠ1�б�RA�fd��i8�G��1䘃��7w��i9j�dQ6��aє۟��N;v��?���Fy7�	���Ʒ���E�;v�z�����;n������x�K����--d��	,~��,�g���/�%TO�&9��oe��G�I�i7n.�p�wd��AJq!3���S�6tU�M���hzb����azQ� �7'$���r��qE��џ�����},�e���[�t?# ���W^QS�s:yV)������l��S�Y&��^�Z�7�hXIY�X��u�"��J�P_
n����#�x���'��sTr+������8HE�9�|�5b��$@8/er1c��(��|�qIk���ZW���J�$O�h懓�8iYI��+,m���o�/N�@$u{)��X(�p�b]Z�CG�cs�m��J.[Bx�?��"ק@1����KԈv(���XQ�P�^�W��ϻ��5(��B�Y����i$���E0�����g�*<�EVY�Wϳ�sS�_��3::zT�^#�ǦɅb�;�QjX��%���Qa�D���G���cJ�TF�^���d:�I��P�>�u��̈��U�@��p�෼G�ۅ�P����x��z?�9�2-���T����G�
���b��ʖ��B�k���v����}�@|<Aj|��	��N�s�r+�1z'a���"���m�m���"Z}�&;R ^�� ���B��Š"�s<[�tb��^�B� �>^)=�C䝛� s��p�2Rͫ�i�BT]���xux<HP50�ve�q�%mM[�W�^�Sٽ���h��E	Q�Ά_�ۛ�쫺��L�$�Oz�a��]�y�OInM���L��:{�*7��Ř�㣡0@�����R� a�8�:����])����"YV�f�Q:)0�!����OC;�dG�\J:+U�q�����(�[e���ӣv�!RS[�~��l�K��/$�u�����$$^��(�$�vx����♸�>L��:;��5��p���>����Dw{�I�  aW�e\q��xa+�O�?DKЖ[��l�������-����3�u4��)%��ב-[>�Ŀ��լ���x@6YmM^�fg����ϥ�����_K��d�ypZ�Dqril����j�Q�B��ӊ_��/�typ �2���Ж:�a�:�'0�N}��D�$����c�=�����b����D�6m�Mhj���Y(Q���p�)P }±�7�u�ӗ�5�5�*���X��a�x��h�ۯ�_���%C�Pt����`�"�:E�Ly�跂��"S^�s����͗�	�X�#9H�w(E���ZJ"r�"�F��:�pV=���n
"ݬjN��w���T#��6�8��ٰ��G�K!j��17]�9:�Z�
4��׮��Te�9��������wfbS���J��Xi��'�&n������֗�B�?�ٵ��J�N�'��� pv�j>��̸"��Y
gu��<�R�Ͳ6L('��a��%Y���T9���p�ҦH�O�e=�R�aQq�v�"Za�
���3�m嶘�A��k\��0eO�]b�NÔ���:vh?�e+Υ��i���|M>Ӈ��c��Ē��t�����>�,��q��ocϡ0��[������_��R������,�uf�pַ��|:A0��CA>����Vx�maz�	��x�MD�*H�p>�/����}V�٦X��\�VU����(FcVr�l2nK��@`?n�з6�r�4.d���%�j:�%tR�*ƥ~V�S��D+9�}���g0����{Z�6`�
u��BI<������EÛ��hnR2n�����8�&/C�b�H�(�Q�-����oiM�%T�ky=ۮq��(v@.^Ӥ�:}y �V��.?1���� 9���y�<'X������>���Ÿ��W%��h+�oj��2���ZC�N1[��2���¬� Lልo�U~�c7�h&�o�����B���L,��ن��ٺ���EZ�r�&�;$_��o�2�x�"����y�#�'�mRu�֎懎�@1�𙔺i�On�\�0{���LE/MݯHЍWc�K��
BZ�p���ᏼL���gwt�7��`
��;i��fώ�k��O�jbY
����-Yv�1$Yܐb2�
$H�4~��!O\^7������<ֽ�F�3am�K� D����>�;�ZPm���3�kotE�})>mQ�4nycn$�Q�vU(wh����VAg���?�1OJc
�A�=H;@�u��X�������=��SE�q�Iiۓ;���!�r�*��Ƴ�GM�����ulp�	 	_�4�(R6��(��ǎd@�����mb�U.|5�
mO��󖦚��J"ذ8F 2��z 1�b/b�ŧ���O?z�$$�Us�&{��}�B���ޭ�i\-�5a��s���)D�a���8��!��z��-K�<��-�W��#/�G\#oTbY�����F@��ý�w�8](��7�J0K�ݪ�w��3'{�)ϻ�`�K~��z�Qw��/�� �R4a�駜K{��5r��vM! Z+�p�������ӈM��*=�4�����&�O���:����?��{�������3��<V�Y	�����]Pi�����4�U�Ƈ�LZVtitF�XQ�d�x�`�
��)��<��z�	M�]E��� ��K�"�yA͠s�z����:�b̰���I�i��w�,�dU��j��F�Ϊ��`n7o��^��5�qO� I{��j�i<�F|��@�j{���o�Z_��d�H�Ķ�Y��������k\x�w����K��d�>+���.��vHz]�:�vO�B�H�2����S=*	�T0��3-u�v'����7n�qwY����$ z�ޫg�һ�ݨ)P�;���W�n ir��<u��kT�+��d!�b?<o�`ꗱ�T�p��{���|������E���oL��k��9�-o�hStyeA���LtƦ�P�j}��!/ͺ$-q_��c�IH�C`��i������	�)���iY�f%�����zfQ�F|Y��\FE`�[*��"�E�.�èB�g�2��b���'���cG���`��QBp��mH��>U��2Xp��ǯN�P��n#k��y �d[�3-�iJ:��"Y�4���˂a������g��=����*R����yr]���*Yy`�<`�`7{�� /Hy\�a�Ɵj�Ú�}ָ:Pt)��,�=��L�
?����z,y��gf�~�D5��oofy+1�3�yMӡ���%�Xn�z��ʚ��ˮbh���b�O3h��%^�Sq��	a ��=7(�x&6A�lT5���ٽI��ZBV���H�jͣ�Y�>��AQ \y�P�]���3S�������]��w�R�e�J��A����V?�:�5�rZ����|e�[lk[���q��iGܘ��'��;���2"���P��1����3ĳ@�>��k�,�\��pEk��ф�x q�4NKL��q�/�0)Ց��"�)������/�$�Y�ƴ^=A��z��U���z�}~�q]̡U��d�Y?�)��Hߺ���y({�8��n揤:�tB�_�(�L4$��<�O}�E��{mﯰ��`�y�vv��_Sϖ�`��1>[Z X����\�H�|,��k�'��y���!�6Jv�;�j�l�s-�7KI�XFv�
�u����h9���X�>�+Ϳ'@u�ɢ�UQ���Լ�[�H����#���J_
G�=�DH�]���i#,��k��q�h����gP��I�:��A�62<��&7���BI�Y���A�Vt�P#����bo6�	n�� 4��Q��B&��&������EK="2�W,�~N{����m�A�)R�����0��?�bM�@�|�2h0�o��\�ȑ�A6@oO�`����^��}�����u���w3�x4-b07��Ӝ���e#'�T��gu �*����Zg�_���O~ڐg�j��<�x�q�Ao�����y�j?0���Y�z+�{)8��,��x>(L ��@f>� �:qI./��q�a{�l�>D�:��O#T�P�df�nC�r�]��gI@�&NMv�@�F"q�F ��7~z�i�ɟ`P� �v�n�w;T���)�N�y����#-G��E`�o�+�` ̟�>{4����>�H9l]�A�C�l�&0���Wn�a��'�+�^��iG����F_�g'3����p0�v���j{�f���Q��I�P�i��*HxՒ��hc*����~b+��Q��P~�T���W�&��H`v�4VR7kuҨ`
��{����_gP����&�s��E�}>O=yȲH�4,=�@Q��O�f���������oщ��*#3a�{n�=�sh!;�x��_�C�"*�Ť,�w(Z�T�;�	�2�����oB��#,J��h57��֋�$?:=�F���y0��/T����l�D���"J���67�Hu�[�@�7Q���7��+i(��;r������W�;\4Ү?����CJ��)����jL^+#�v[C�Pfl2��5Pi>,/>�_���B ���R~۾B�p壻��iӸ��5����PR+kQS�n��/Fn�B����1}:��ӈ u/9�K}��?�L*�IB���Uw��Go$��^���̽#�0�ϒ���_l%�#A�g����E�:XaЀ�}��������k�g�r�Kg�VG��5|m�2x!��5��OR�=md:��{���%~�dkH��	�#��[���r�_�ڄD?����l�( 5p.$?�*9ѻ��Ч��Z�����>��veϋb�\v]0[����V��Í�5���=�20�bI13����=B��v�$ߡz������X��ca>���
�Pd?�N�3�u]�s���H�xZSo!��=g�vstz��E�����`�Am��@z3{GE���%h�FM���w�3��+�$<���{�:B���_���@ӡ����U#鏲�3�V�Ԕ�����2�&�r�&7����ѐ���3D}�}!*K[���Kʧ��#�m{6���7��3O�Z��kr��gO{���Q��, 
��y:�7P��Pc�+����45~p����mp�dme�5%[Ce�E�d �gbRa\U}D��bTN�j����R������8|������w�8�j�<[-ǹc7BYO��\�����A>��Z������k�f�\� �I2X���y��.w|�)<��S�������
��!0�E�������R�_��|�W'��� H�2��po�(��x]#/UFʩ��V�̹�"���^�+ Qn���>��{����R�)%�7�֯+X�#��Z0T�U��Y�}�S�"D��a��^$�k�E4�v��~g�у�bS��1���RL�Y��g�ٻ삉wv�0���<m����4�/K�9���J��R�8��94)����Ũ�cu{��~�ә��3���;s��\�%�^L�� ��bWP5��u�Fz
�ǒ�j`�d5U{�F�����O�zg����&�`�9�p�e���j�d�Z���1�cfӟ��p�o�2�>���)i�_�x���X� � ���$uzc\�)!9/F;�jEgqa��@3|�&x9Tvn��f�w�i���	�l����Ҟ�0�Oj���y�M��q���@����I�m~w���Ց'X=Ýf����Z����7�=,��tMѤ�C 9��5%�c���un�)�Fw��}>�����܆��w>���	�8Rd����d��Chq�<~Á@%�<<t��DX<�HI�#���5�>��$.��<ñx�[��龍l�Co:%���*���$ HF���?��Yޕ��K�����x��:L.����ЄL&��7�:�Of%�fM��2rT��@n��)���0
�Tm�����sj�����[#���26�����e�l��q�.G�e�Bȳb$��'
��Nу��n1i���ֺj.���X��$�� ��nsk6L�2��_� 8_h� ���:Y)v@��s��x�JX+ʳo111�v�^�@%�*5���3���p�c��_c���\W��5 qu��s~���'5�e�"��8Π�[�$9��/v�ߠ�ђpw$��H,Ҩ?�Q����ɺ+�>s} ƍ*��E���0ﱈVo�P5Hg���s�:��A�]�:���+f�gg�E�6/G���_��m9!EE�#��/"is^�{�sѶU��e��E��*G7��)`�@EձI�I&M9�(7OF2F�]̣������X�>���c�˾.<Q�[�L),�?d2{�isc��!������*�16�]k�P���̠�cpaq�hƟ6�jb�T���T �fy����f�Pԥ'?�~`nu����%�4��#&>������ЋP�u��X�M*qN�!q>���`��)�ښM��gE���Jg�m�ͫ%i'��p}����:knV��bO��Em%[��4n�+a����>=���H�nKG7�ڪL�h�C�5��o1���b�n�ׂ��TU�=��������(��
��%+�i+&��7��h�a�H�0k潻J{=='�[E7ި
�[X\W���.ǯ|�Ak
�Ǚ��4��������*@ӷ�$%G�$�b�ڜR�t��{�ڄ'
���!�W-@�O��S{���~Ku)D}�-;k�*�m�����Ru3BU�t�c��i���>��U�RCk���h6�w�;|[<�L˾a~sYJ$��P���6��բ�`}x�fS�V�y�Fk�`7+N�g������BN)r�p*� a�{D�����o@�]�172��#�5����z��#yy0U�C��vZ�c�,��*�є�l�ە���n�&�F^�_Zpc�G5�����^	���Y���ɫ�r����FX�)уg��b�ŅL�&r� ������D��H��
�O�H|�e5����WY��T�N�4�ą[a;����?������yE�1��H�Fצ�r���M KA��i˄Ռ\ڕ�Q6j���YR�Y�19��K���hf�b�NYm�Q��/-�����<�C:�iJ\�[H��FB��/�˓��4�����Z����bIQ����eY�Y嬀��<�Kk2 <`*���W�4����l��}~L�K�_Ɠ
]�v���of�#����C�P;5ۂ������u6�!>�?�(ٔ��>w����M��+b����V.�HJۮ��@5q����]�	��qǸ!P��P���[w��� 
��Y�F/�ا�����Z�>��_w���oi#��<{G��&��1)���u��]B�m��	ּ7#A*�-X�U7���V�9u5��y(4v�ă�C��v�\�,Ԕ� �c�W%c���
�-���Љ�3O����Z�|���v��fo.�����>�M�x���&�[y��f��S�M��.�����ZQқ���#5ɹ�Q.����-[��� a��Q��5��#�#@_��O��,=d�j=��'��oƺ��Q/\j�O� �{"�D�2����/��׃-�����Vb�7�pV�fv"
�-�ܑ�[���ZS��jҷ</7wGñ��2�Z_ RbN����cK-��t,-*�) �ӻg��jMv}R���J^=�]�ɔ8Z�d�
����\��R*�Z"7U+B���If�U�f�{c�C�{����Q���@��;��
T2�l���*T��]��a���ތ������JᑬPB@v�z2f�¼̆�R�м��V�}L��q�5��ٺ�F����<,[���E�=��	n�"ˡ"�������( �K��G��C�幥��m����"�����9!��|1ȑYf#��Li���*��<6�V��H}�Hӻ6mj-�§��jBl9�Yԉ��k8ܡ��ы4Us<_v�%đI���R�����AG��-LAY��V��zŭ�3\����þ�m$��{�����z�e:#�+4v�~��[�m��!��;'9� zp�΃����#;�e��U���c��uP��g	�LC5Q�-��]��jp�Wvg�I�U�9u��ï��z+5k�ut����1uu�půs2��^����DX��aUڼ�ld�鬧WҨaE �G��x��������TQ��1F��{H"���4���+�o�P�������/!�'�o-�Q�
M�FT~�}�y��sU���8��(f��`�."a[�t[j��������T5w8+i�U��]{4��Y��ƾ_vi���? z�u���׶��_���M�ҋE0��x�oN�/��>�� 7:����� ���׈p=l�����΀*g[+��(μ�.���7�:�N�s��}�����V�A\�֓��jd�pgVV�����a����=JCs��Q�sf0��Q��#Ì�?~%���+���3;���}<�����tM�cy����A<$	_��xgu�z�^�*TPϲ�Ok��&�l���>ͷQH���Y?�d��v�}r3܍Bh�>
��+i�/&��	��Z�<��\�?w�X]t([�8��`����Qlf�)�f�3�B��#ic������n�on�(7g�*�G;?<�whqGJ$Ǫ�qY
���<����N��)G��{׼{~D'+W�΀��
��󀟆ktu5im%��Wb�]-�۬�֟?��/%֓����Ê	� ���7���i���2�u�[P����j%Q5&;�J5�HJ�-<�a�|����'5��cr-]Gz�B�X����hX��!�A�7�%��H�J֥���c'p
����Tpb���M_�[!h`5�O�f�MF�]t����|���]���ӳ��c�K���z�^�~w�I'��K���c����J��):������Xz�	�����6!�?�M��6t�w��-3��I!v~�v2�s!x�/�+2�����3�g��i���%��;���W��"/ !Ժ����3Z\W�E g�w;6��bJƖ���O0q��T�jo/�!������Hn�j�+���/�V��k$���f��y ����<Kq�Y��.�j"����t��L2���4+S��|=jo������D���?t��N]?�V tZ���n���Y�&<\�|��'j�����4YYh�(|�3� x$��P�����
1J�x����qJ�FN�fH���rt�@�\>di+�A=�G�Z�_�x�_�UM���/��QI�� �;,�UVn�Jc?�l0/{�r��Y8kx�mt�Z�6�)�>�z��+H��M��S���}=sŲ�,]>�m�kkk��`��VW��y�Q��1��6��H"���	W/��hn6��ΐͥ�
|�.��,|�\K��z?���b���8W�ҶPp��U�������RH��\2�b'�����Wj���*�Ԉ`��Sx��������f��(.k��yb.d��尮��6�q*�,�yK�_HM;��K�qo�sߵ#��@��R�M#��Q�?�uҨ�����ed�Z��C���p�aYA{�m9��B�F�Q}����o�hը����'�����>�	��1�٥�JC�cXQۚ0��ѻ���x��T\�H�� oX��N����S��?%��UT*�㭕#�q�����jꜬ>n5��mO����Y5L�v�@êjj?&V�|ˬ�[�������1U.��q0�O~�Sᡭ��z<n�����`"�����t���gЈ����Ua!|�x^��7i����8>�,����y�vA9P@�z�׬$�j*�
��D�H�����&�~�l�|V��@�~㿄�[�`��O<�(�d�߲�Dv]F��P
��B��7�zX�,������a1K`
_�����4�u���N���ԝc���K}�,r���~u���p��,�}�e ��o]85;�Ĕ�"�@�K��bK�ɡ�죸�e���N�|�J�3n��r�`R�صnmc�iW688t�kCOO=[�u�2��p�x�K�؇��|\62Yl�O���0����]�fjʯ��󦿘`hX�~��G�p5�i4�]=�:��
������:F�^?�fNn�t�pIG"ǹ�>,vo����a��?>�[����5�PJ��Ћ\}S�����	FE��cZ�s�[(b:-lG��]�艠#��/񷜁9tX`,��?���>�4�i%Y� h> 1ZY��B1Mݥ��R��v:�8SR��F��Y�~0���mۨ`@>Z�ٙ�s�<񭭩�?�J��m� ���gve{]���i��ͼ߻������q)V�5�A���#l�}s��"�W�`��s��,l�;�c ����]�kdK�k�ǎ�.!�;���\�hX�8�/��6^^
�eg瞮�2���S���c�E�s��JM�KAHX��߰αc�ﾵ�{۴�&�jc��b]�Kɤ��9k�R>�$�k#���+����#M LJ�����ƞ����V8tc���A͖�>t�h����#Y����k�xl����v�w�����Y����ް��s����;��R��'[��䥜�k��X���/��r�]�ģ������^���`)�	�VA��Yֲ��׳
�߭z}��}/�bh��W�,y����VS��k�eD�����o�7[/,	A��n3�NO�9��ïBWy����G����Ѧ0<s��(P��Hp3��X�\��`�L���A��J����`%%H��-����|���]��[�粨ۃ��vL�<�1Ʒ�L�6��?̵W,��I)H�\7���<_���0\üԥ��ɝ�k�S�E�.p_۹V�t�C�΍}��#WC;��']W/pN�5 ��#�Շ&��cgd���`�7n��4�����4���>�
��i����v�y�<�]E�y�^�x���B��~���GT>k�cV�06�~j�s���ŴlP>�Ý;[Ŋ,��"�C�g�.{�~\ы�(�%01ݥ�T7���������ū+s�g��p,b�rҠ�����_	QF�{�1���&n��6�I1¸b��������, �f0��S�_S�&�:�1�;VwP��^�@�ha��C�q	9���t�������F�&���},��u�C�n²�R�t��OPY�U�U���K��;v�?TM2����y�Pw}������-������,¹	v�rɫ��)�@����K���^��i3Z��A��v3ͭ��}�C�o���k���k���4X���뫮#'���1W�5�x6�� ��ܼ�����˓m�e�PF�����z��ʍ$��7��KJ>-#��=��i�K�5���ԡ� `n��K���k��B7�K�KK0���b}��T}\��7�6��-c���pw���e�� �?Z<����5Pn#~|����vM~݌��gS�`�Y�8��\Mn�=gZ�aչ�RZV�T�D�#������7�x�0�F��wv���N}N|\�t�י)�o�w�9��cc�I�_���c���_���x��8u��6������^�S�98�"D�nQm�E:\���{i��|��O�^g�~)J�S��r�K!�=���S��m�K�8?[�G�/��:�E��`>����>0�� ~��A���L˟��T�>:#lI��D��l��ͺ�1��諔#e7F~<>Gx�-#~�Rד'4�R�:4F���̓�Ca�;C�^�~E<�2m1�����h'�Ӯ�T�o<�Ɠ�[�D?0`SU��Y�n�Qz~?���4c+*ԡ���A�ǃ�h�Ɠ������}�q�hR0t/%�!�������i@ּ�>;��}��V7+	��ƚ������w<,�����Kg64�a�`R��Y{S�������wR�'+�[�'�`��et��*-̍�咱�����?��D^�(V���v��3H�z��2�T8Rs|��"�:���ˁ�kg?�D����?����{���O�X�#89�M��Ժ��WU�G���T8��� <�+�,X�'��ݮ�[�+r�K�A|�N�>y �U{χ�Z��_�2�h���k0��O���/<aDS�U���������Z�lJ��ol͏�m�U���V��Vmɳ;�����pA��m��P�/j@:_�'so��g���54��H�ռ�F���nJ��<wO_�/Vgˠ�a��.��J�[2�ZY�l-�h ��
���V�
�32���T��$��M�w�G�`�z   �ݭ���f�7��&�qz���r��/6���я:򃞃�hk��g����NNm;J時�Nt��Rn����Ϳ�*�"7���"�"N�0��s�,�LG��V���/-ۨ&�'~>�;����R�Q��H{bIN���� �mG�f���*[�R�5�Z���K��i��!z��b+e��;o��x������$$��0�)t^���4��_��+-[z�5��VS�wW��ʑ���x]�;��2�@L�D�?R�����*e|yrg\E)�x��)��DV����������bP�p1�����U0�N�����q�̕���ʷ���0��G���F"Q��^7�a0�^@t���%��[�ԽN�<s��	kߨ�j�J���dM�S�����d"9�����Y*n m������l���Gg/��mZ�f�6|����N�p)hƥ���z���+V��~s�t�	02��h����FX(gŗ[��Ġ�Z����Ɇ���F�(+�H������I���/��e;JԘ�V}T�q{���(��e�g~\BO�6����(:�n�k6��e���99��}��.���Ҥ�%��[1�jo8 s�	�����f�ry-t'=P�H0����H��9u�,��IH��F��tcN�?j����*�������S��-��'�����3x~~~���у�(�8��0���z��;p�k)����D%}y�����}\}���T��E���h��#:�A��r�����UN��[R�}�x{�=���,,~N�@
�S�iwZX"�?][��$�u���ꕘ���u{�y��{��|N���X����qm}��Y7+r�UQ��QjX8�՘��{���5;6�`\�B#�`��T9$]�O��Q�LB�ԩ�T]x01>�vR@����UyI��P��O���o�
.�k�P4�}�E�eW��̬���77����wO��UG���h-�oW��X%�L��!P����{�5�^w庻%{;=���|}MF��7WLJ���:cW�|X�8����w�糪���]r���;��6�Ѽl)"o���,.Vy��P�z� I�2Q�E|aJ��rh�jGW�A�&q��.ǈ%��T�P��.�|x�g=%������^ڒ����lQ� O��m���%P҄,����||�XG�w8����<��\[��۲4-f��<���@�>��c��Ѷ�C#*t��$�O�w�6��]��K�ђ�s~�fW;q)3��>�C�Y�����A-�Ǜ�S��>V����j�9���
#N����&�d�n_�7��6|�$��;��*ka<�/� �g�D���ڏb�\�/`u�v>�O�15�����k��;v%� �c���{d�d�9���c�_H��6Qp�\���p��kx>X���5G�k4Nm�P`�E�Tt8�^��O|���ީE-,:<gHB�'5��Q$I�I��6&��O{��ׁK;0��$�ޒ��!�;�(�^kZ����Ky�Z��N�jhOn���J\�G0�!O5�����y!��������E�ꀢwS���&�o�>̓�17�l�_�[�](�
�"_�ʢ>��cϊ�C��À!�	zy��8c{\�"Y�,���#"����o���}�֒��+t%��H��o�4(��?K~G
��-@�?��rG�Z����P4=�'��ܰ ��û���`��Kp&�2Z�T����X*��-v����=-��
���g�'������䨰lה�)]�MN�K�"��A[�{��.�|����4C����b���%JTY[[j�>��S-�Z[�>V�b�18�=w6QA	,`?:�f�֯pm���#�+�.�FO7�Y����T�V��O����r�l���Ӱ��2�$l��.Շng�]|�z\�W�2K��?1=�[�BK���������:�quq�c6���ʨ��IByyC�wq���z@�wp�/ZIi��N���:���.SUE��Q?w��5:��\�����;Hh8:܃�HPsE	�o����]���_]}���I(��*J%��5P�ꕾ�:kk��JsZL�l��y�4WS,N��66p	��
MO�y�L�� ˶x��~=:�5:ܴ��h�vw�
��u��W�X�T��V����u@�W)��/=k��N�����TR:虓�P�i9������|�/�ˠ}�7�Ι��U`�1�&�����b�h{B����Q論�_��=q5�����Gj���*V�;e��ȹ��Ζ��dkZQx�oҴg����M�>������+� k�v��њ0cK����*�x������ǆ��{wq��w��s��4�ͥN��pxe��w8�k?������@�{ۓ	g4˻`�s(Ԇ@sҘ�\����l�>`0Z1x��������b]i��۴^�'����it�jV��\�rs`��\�Bu���m�	mL��f*��=7���[5s��]۵����i��������.q��)�ˎz(<��`h���P��O�o�s��'Iʰ�����w�ؽ���x@�ۤ�O�>ͷ\���wc ��2ld��?��S�˖�1 �?��W|��j�|h�m��^>.NʊU��W�0�v�ua�p���X忨�A�U��^c%�[��&�߅z1���xJ��9Ƹ�y�����RCS̴���V �߷����2��k�� e�tW���MgU�~�!Ei%��E���A��[���A�[$�F����F����=���χ��쳯k���{�;߫,�2����H۝5��7Z��Y�VF7��^�k���+�B��x҆O�R���LWr����IG���;,�Ŝ(�?,�Ṉ��~ޖbtr�}��󇏱��=�
{�ҲC y�Y���a�Kt�[��@?O^>$��x��\��V�����7���=ϳ���*�W@|H��zz'Wm��4��P������܌��|�Pd:a~�]v��M�VI��$���^s�i�X"58��xzz� M�	�����=�v�=��n?~�����C���q��/=�K_O����hr�s��}�B������U���59攢򭖓7��mc�f�m4L^j�-����j�jJ�8o}=1� ��wv6�g��c��G��|�e]��SD1H��y��V�H/x�bDc��t]ʿ3i5��vC���&T�y�C��5N �)��QI
��C���DY����@�o3ޥi�$�/^���4����z1@��V2���jb���i���������i�/��ތִ��̧�s��ܾJ��#,
�I��n�9�����2 ]ѿ�Ж�߈����G.��x&�j������ROk���6ZVx�#�=� 7�:�&�*Z���)U���R��Lmd�]9ڢϑ��d�X?�z�e5��-����	��E�iY�z�����s��q�>ŬvY722G���k�+ú����:F�:�pd��p|����Aj;,���m�ڇ.g5�Jļ&K��0���v��H���V@5��T�J%B�"u������golile%'���ϥp�7��s���=��iY��8����#�p:���L"_�=C���s�^Q_�.�;~D�!�|LY���n��U�&�
�a�1��6��!]�ߙ/]'��hS�����������_Dy�5P`�j`����N�8X�UM�z"�{U�5�p�,8�.I�L��_���߿��q�Ve�EO�O�KT��&W��������x��'%�����K&���	�o��D��%k�>8v3@�pU�l��d�
L�LGߏsJ�k���<c��R���z�4����l����k�=O˟��.u��|�8|l_ڈӯ�bp����J����ݿ[�ؙ��ݥg��"+tm��k�m��A3��]l3��~.�����~~v�S,���~�8u�;\O�j��X?�	W�5$���o��S���~�V�����ݲ�m�2B���d.56iG�m�\e<�D/ � ?@v��
���K��g�E���R��i�}p���0}�7/�O�g�N�$���5�����Q���H��ʩ����_� |�]"NQ@�1�!y7�n�ka߀7�KN;��1-�G8Gd����!��罓���,�����\��X�br�#��!�N1�h��\�m��q'��&�A����g. ��LF2b%�%3_�F{�F��a�����v&� �V�tU���I��F�fy��6z�L���(���og��lZ��AC��0C��0�+�ZN�~�s�¬s=�_w��pR֕�d>S�t���nS�����}��`����4Q� vN�6\��.��"$VւcU	ls~�^��Ĩ�l�F����	�����C���y�s�?c��v�߯=����,+��s޴�<4~��N��B���iF������+S슊}���1�gנ�� e�UWg?���.r؎�-��������aݏ�$��wD�{z�+�:�+��d	���G����p�`�"ȼ���P���ʭ��䎳���AhX�o���kŻ:7�(��I�<H8��	�@;��w�`D�	y�i�Z�F2{ڤ�tv�O�Q��o��p3�Ou4c�w����1h��m%�k���������㜇�LbD�eC�����ȶ�b���XIp���������9Ek�߂Q%�����u�1V�}�����A�">Ԋ��]�l�G"�Ӡ� ~)�myo�9+P�~�!��Z�̴�n�X?~Nz�O��_�֥�S��ʡ�����+��7�|�ꑙ�rƌ�]�ٮ��}���߃�{qN��Jr��T�^Z�Bw^T�N/A}�L��:/��X{��0�q�;�����������
2���:����T�ɬ�J�\z�0E����w��\]�a1�E,�C�62���Svk����d/�7i!��B���ʎ�<k5.}�?t;6��<�m���SL��5 ����;�:�G&��W�G�j�G`#����|��U��{^��TB��0)���&k�����mz$�N�Z�I�0hm�����AE��5�8x{�@�֝},Ϡ�R@�Kr����^���������I��sJ,��NayAԝ��Bqz2	?�� ɯ�B���e�t�ڿm�34Oɢ�P)q�Ęg]�0����u�ߧF��9��Wn�i��?��и���>֗�\���v�ױ1�������[��wd��ԟ�_~���s^"�ܷ�:an����{߸��K%:4̜kxo>�f�*S��t�g���1�(��b>�鿚*C�0sٺ.dG�丠]H�С{{�QXh��v����i�y���*�6����MC~��=�/B����.3�o8����&�c��2L�ֿ�Dd�6�`�4!+���jk� ������mqp�XG���*��}i�d�Bɑ���ς�����_c�h���dwW�-���Ps����e�|���'���P'��jV�>�'�6�C9}[��4$�1�9p,Aԫ��{7"�-�]4�I�Ƽ�B-��@��+8-2�����l�|Rd*�H��֥�L@u�á�#3�Mgݖ���_��T�JĦ���¢:��l��4�i]6~Ѻ:�����˟k޽�ʣ�8K�%~�}��;��Ct�|����#�VY�VxT��Uf�e-3ֿ`{)��2�#n�؆X�WV��5�>|�\�-=�0bՀ�ҞAQ�A�9�7ϧ�(�2���d�I���J���L��ǈ�<���l+?�QQ5���5JV���RS�aJ��{���VZ���[};ˠ-�b:c镊&���z,�0���\��ǣ�є�sYh��֛�����_����c䨬������R�>���۝벗�?h3�F���[+SŞ����rh���	��a�)H���I)x/��L���2�"?�A-6n��m��A���T	�2����Q�	��vދ�@�}���l�B�+7�w::+g[�չ��{k��i ��+�DC}�f��V�-��۫Ӏ1�|*?*!��sa��FP���3��U&�����`��&%e�mGr��[�m[+w���2����!��G�>k�t!$١H�����J��k�q��>,�W{ONk<<:zlD2�_�ONz<���Q�Eg�l�JsO�[MÎL%b��	�߰����b}WE�6�y��_ف#�� c�k7�qm�=���I�\�tG�[�����\l�����ȱ���f�V�S����!gக�Q[���)uЪ.��2f��9_�#i�^ tJ:LQ�_�z~�z�'-�=���vQ�a�xRXR^���	����shR�)�'kJ�Zs��l[�[�V]�B�1益q��f��Y���c'�.B�qK�q�����@�~��!��DEE��}^}
R>3�yCX��j �V$�;62|[�}�1^�N/C�dVOZn�;Z���lT�I�R�~�?௩YA=� ֨;b�T�΋:��V;$��a���x�j�c���k���p ��<A^�S0zCO���ο h�:�@�Fq懚�H򞪗7Q(���S�������T^j�>����D;�̊���b��0��Jl�������]><���ׯuUK�D��Aĝxhp��ߪ! tԉ}�+߻Rj��j0&�Zl��;]!��5���m��^�L?2���}rv�:U��3�Ώ?�t9�!2�Z��(\����c�Y7�uJ|�)�$cha��)n[�I@}�"9x�����4�}J���Ҳw� i�DD|�󞙆a�'%!q�A��Q/�G�1�sko�.�ϋ�v�C_��O��]H�tSUQ���nd�Sz/gm�Ĵ^�sl5������.'��塢$,�N�K���\rg�3��^ȝS���Qm�&[�$s7����7��p�8����JKqj�����I��b��󬵋T�l׋�n��7�^��%Ϭ7%��ht�Rʕg{{�|��|bb���s&*>�.N�b}���#Y81F�D��3<�)+�K4k\�ݴd��cK��-��ap��@%���Gy�� ������m@5����Z����-Ό�"��~�Y��c7D���ZG�x�W;c���ks%�ԖhE������D��"oCV���#y�V���C�B����a@��C(�CD$1\�c'Aȶ%7yu�'Χx$n�6��f��OF757˫��
�6�U��w���n�cm�u�v����-�J>�ɶ��[���蟲���s���C��H{��;���)�K�7��f�ұ��@-\j���a������D���p�����[����
*��ʸ��@�+rr}��t�b��z���Z�X��Y:��>�q�k���_����ҫ�fC!�'�ɯ��LfZ#��1q("Ex��� �tw~�Ŕtc` �4�T���o:cd=�9�Ix-������7�Lx���o众"�Lx��gT.wVt���i�o4�^f�����2�fY>�5Qri����O)3"aI�����!2�K��4��O�!9',�`�ۘ�B;>~(����W�Z��X��g�:����N�+=��	_('����u�_�r�����*�q0��j�N�l���L[M¸�Xdx!�W��i��X����1�xZD�T�}ڔt�����Z�a��['�#"zt9a�1����wO����_��������<`hQ��*q!�	�P�uz���A�	���(��W2��˱�DJ�9Jbz�6A6�.��7A�|i/�SK��$�/VV!M=��ڦ8��[��聳8��/�s�4nwW��f��A�X�l�GVm���<G�UC�`��"�1J䎜`��^������E������s�%r��݃�c������}*A����y��ᱵW�匛���8�=���M��[4�bB��O�f�v�ȸ��X����=LB���;�"E�<���M��Q��2��3K��,"Da���ת�p��.�����1�f}���TC�>:�uu9��s����2}������սo�0�#BEO�A��_/�
e๸�ʗ��S�a�ɜ�O8�VGA������X~������_��e��yWKF���a^�j��i����>��d�݇2An�&��6&/U�����7b��$�x�(�B]v։�tE&�z܄a��є%�fk��8P����M�{{/�S��z2%����u�mݙZ��9>��������!^�/�tGh$�;���W(nK:����4��cf���Ϩhu�����Zs�w߼����We&�$u9�{�~?��?�y�;(RvͻQ&���Ġ*��B2���T� ׼~R����CjF��DRa�1�����<� �C����.�v>�eOF�l��9rˤZ����1�eETux;������m}��[�y"��e,�j\4��HR�Ϙ3UV˕������7����FF*��?��,Ty��eX�6�ݹ���r�x�-^h���EK]��	{g�4�Xa��@
��`����g9��HG��\�рئ����w��CO �c����&��?���جY�t=�W&�m�����)Lm��\���2��^��Cȓ��w���BB �#C�m_�NLA|Iu�YmXK��z��e��o�[E���$%��0J#[�=�ga���z]_�:�N��S�K!�B��a3���MI(����o���}�����3�G�d%2�S���.9�/�T~Y$�$a�3x��HVL���Ցjn|���������ֽC3��҇�t9�LTP�4���J9'�:\��] ^��p�U�\�h)u��,�����5�"Gw��Y�cs��,y�W���SD�(�BW'��|�v�uǋ/&�}W &}_3=I��3ܖ���؃6�fe���V�Lk��_�@�a��Y�Ư致ȉ��������kyE���^�S�3a��>lz|�5Ж���]�������^̓fc����Ek�'��� ��G["��@�C�|����_kr�&aP��Eo�ŷc�q�[��;i���>46�H���RsW�<aէ\H��4��R���5��ūF����˹����끶���N20�>���s�����KA
�0���7�f_�`�	�z�Y����O
�?w�6 ��q� �~��}F��� 7�k�����Ŕ���Zc�~Ԝ�f[_z��tjH@8�]uo����V5����m���́~��y�&������w7TbOL�*y]x�=�'��SVl�U���ܸG��Q�I�,Y!]F�e\T��m8	���S呈/��^9�9[�1'��)A�Q�qDs���~p{���b�, ���RiȠ���؈:�=�3'��U���'�y���'|nO��r��7��,	yZk����ڟ���1�$;P��������~������"��PB��c^R)�إ�J0G��̰�5��x~�=�Z��+P���?�t���������K1%��Y���f[ķ�Kp{\����o�����7�4��y�H��^[h��\[uINX�w'���kC�ܩ�8Y����;�f>\V�wg_�F���)-�J�+Æ����iR�Kݟrn�~u�2/�������rg�L�k2ѳ�v��4�]�����������v7i�f���=�+Q�F�ë`�38�N�͠�r�e_��nM��\\\��7b�U� v�w�8�<5��zx�{wC	���2'�-�Q����o|M�r�s:"{�����M�v~CCCe�y�s�L� 1?��2l|����i���L���������A��2�����2��4�k��/����a,�F�����̣/���)c���]��^>M�t��Mܶ8�*���v�&=#���_w� 8bg5C&dR��������z8<�k��� �(n�hwo/gL�����8�o ��z�#����b[YY�06�͵�ѻ.�cS��=rZ�SY?��^	��&k4�\�斾��������H[��YC�@8j��=������:
f��s���U$/T@���lU%$L��Ю�&�%w�S	���a}�~BO�S�Тk��b�5gв~n`�Jab:���V��lsNG���ѯ��y<i
G��t��@�I#�4JxTh��+v�gg�+�KI�(���QS�^ۃZ����@!I�b�h������f}��3�1#iD�����\�:��8\�pBZ:�,V�d�v�����ڑ�}����2���Җ���t�O7��w��鶻6L�8�A�A���;�],`�~ΐJ��Pt����������i����^v �)f�y��(� �;��F�UL�ٷ^3����}o���	�(V��4wtT6�8aV�.��,���v��������Z��\Z�{e'���L*p�K��T4��(��b�������ƖS�� ��B���W��A�YBrZ~��Ď<{���)Vl�{�~���a���D�"�+m�s��n�@;��%��%?}��x�čLZ���I����&!^�L����O�XΧ���D������M#�/�
�IC��3~$�P��|��� K"��m�3ڶe6�8��[FȒ.�Mn�~�vsw���;�s9��O#�U0A.�c\Rw�/�!i�#�7�=���i�pp���Z@Kd ��4��4��gzi!�bg��u�9୞>�f*�˳q���U����mq@��q��	��?�fe)8KxKgQ�3k���鼃#})��	��-`���m]v�̤�d&}h^wy烑�ߔ�Y�Pa&I�23�-����wjl�)u��L����D������c�f��m�О��,�=M��47}!������=�=/'�������M�ƅ�Z��D+}�r�e�gq��
G�٨5��:��a-ψ>-nd(R$�|xI����=�Y?k�1�\27[��8P��_�����h�}�(;nB*� !���N�lh[c��O�U�q�I\-N^�V m#�DU�>�UD8۟�q��0�w�8���2J�����
�$�/���<�7s�6����N
�jJ�WNl-ez*.��y?l=��F�i�=�7Gtv���<�tWc�ت��--z���,yF)C�2�Ӂ����͊�@�$1?����A-`x!oѲ����8	��/jf�)�w�g���p!֞����ڡ>d��� 	*=
�}�!w��0x���:�_����+G��lEx��~M����egaꐉ��p<h������+�	ny%�n�0��w����l��Չ�[��q�
%ыϓ��+��J+I7�E�"�e9n��h*�o���>���e��f�����3��*F&��7�X��0mƴ"C%OD�"&	�'(Q�`�,�mN�ۭE�ׂ��ܹT� k=��ç��&^�`c�ڋ�Z�r�K�H�h��Z�1�RY���eR�!�3��k��v��j1˅�R����%/��)����6��Y�b�=��K���W�y��؜���$@n�;��iŇß��KoL�_��ˊ�?����7ܚ)HIKS�Ho>�BWS�^����쿇/N�'�<:}i�5W�~w�������]E �x��$+o⺝�F�Qpr͙��(�=��T��&�`������P#���uĞ=��d�1�����No������v�[��ZUX�~h�������k�� Ik����f��<�Т��9�k�����Z���t-	�dgA*��㬮4[z�� Ő�f.��k'g<���,�V}:$��B:yp&oǧ�V������VZ�h�8y=~��/qSաW����k��H-97��2vSʪ����{�v����CCٕ&	����SN ����k�,���l��WF?����1�N��Y���e��a�b"�)��O�Ɨo���������)���;	LH�1�+��A������BЎ}��b'�v]�>B�u�),�xI���l����㻻�oT�W'��э��yx�����f�J�h/}*�ׁ�����ɥ=�P�%�4��@LH��	��F�S2k�-o#1a�@1md���� q��OY�vF�_B
'@:�W"7�+���a����W��]O�ܞYܿ����z�ក�'>��;���!#�d�ћ(v`��X����%��!�Q-=������S�B7F���b_P	�`������&�x)T�����Q�QU�6��/�7�\^֎#��Z���h�\�=�1'q����.�<}A��s���;{D@U��:��əv��o����a<��i���S1]˯��H �X����+���KƊ�qc�I�Je�u��Z37=#�x���k�P����R�z�Ȥ%�Q�f����yᡛR���!G#��T4w��tD�?�������.o����/Þ�}�x�ě�&��{]E�a�Xt[fr:�Dq��eUf���.�����C"r݃��V���u�Qn��鴄�.����.�AZ���q�9� �i z�Oj����$�.YI'e�ǋ��ӝ_-�ɗ��}��	�l�Pd�}"/8�u|a�в�dZ���r<q'���n-S�z�'�����e۝k�~�ʹ][�������뉬�a;/��ƍΠ�PI;w��>ǭ��12c�q��J�^9,I��y�c;hׁF��OLW�����L�\���)sa��-��E
���]��7@�JY�ښ۰� <�1y�c�K�0�H <��h���t�7B��7U��n�Ϩ�@����i��0��g��N�>F��~�8��O=����I΁XnY ��.��\>κ�\�M�I�.��CM�e$8���g�=�"�7[bo�U���� �\�@k9��%�Ñ+�[6�&�{3Ҝ)�@�֎���`�����;}30���{x�sܨ��ҠQt�jta��&����cO:±'3���%���@O�s􆧐�p0��Oj���yX��F>��&c��'������E�0n!p,��+�qx����ȫ�D��\׭q����ߒ��-���ȱ�tp3:Q��o�!N���Z�Q�o�Z��Zp.Կ&�S�J��*�A����e��b����H^�r��Q3�8.S��A	Kb��?��y<��{�\W�D򒢓�h���g�' {�v+���=�ITa�����Q��&::А�뜂�2����O�+���z�Y'��Ǎ��G%�P̿�&�����2�u>�����{_��fs�'�ڮ�^�KT���?�ta��ׄBe��MD��%sJ�2���߶�ʖ��7�	ATJqqBC}�b�
{�BI_k��،�W�%�F���D���IO4na��7��9�Ҟ5�t�Q+.����"�W	!}#�gz0]A�X~䧉�`2���� �泀b�]E��qg�E�;��3K����P�l�%1G�n|u��)Y�>���B�-����{P�8��������Z{�n�VV��.�dJ1T�'�8(=�i�|Ϸ�cN48��CG�H�!*
�z,�u��L�u=!�����*�b��'��ɑ�]�.�&����*3�(�i�A%s{t�����uW�P�;�_��$
�HeM|��J2�TQ �?���ԕ�}��!��?�~�6�Ϸ5��x"���ɬ��!�if.Ш���I�����
?	˹�u�����`��t�Χ�Oy�c$uI�F76�@�oM����%Z���}��U�$44xҚ�(�Ç���zߝ��÷��`��LY^��ȳW��=|K���V�L�jFvw)������?.������+�������s�g��Xh��4�7�ōr9�� q���p�d�* Vh��kZ������Ϧ�y�P��76�ttj^�� U�6��a4�x~h��A�3)'��X�<	/c3�q���3�t둇�u��Mb�5\����X�6?�$*($47�+�9k����=w��6v��գduBB*����s_����7�G\�ZO�����z^7;�(�um]��7N�ַȔ�j�I�~w��!���~k<\��LR�j��F�O������'X�[`<U�1�8<G2�Ϩ�F���J	��
�]�5*	p�WKOW�R)���gԉu���6�hi��T�˕�����Ɇ�@oP@S���8�f&��8�Y
n�d������
}p�b����|̪~\��^0���$Y���cϕ0�����c�#M�Ӥ�E����`��Czq��������žag�����	|�g��s0�^�v�l�7����p$^���
�,9#<nJ��}i�a"}���0��ރOpٖ�L:�2T���	����h3��U��$kG\B�a \�{ X%�G6��mz�s�(@p<�|�X�; #�_z�����������i���H��ԭ-��<M��0.7�����FwLt���tt�e���JwkJ���m8���<�e��iK�����P����r=RB܎=�Ƃ�-C�ĻR
�C##,SNm}�'�[H�����/���%�xӸ�3e
-R�\V�:.�D�3*\U��B7aG�I/��\�h�8�0گ ^��aN�v�4(��qA\T�S�=�V�i�( P\��:�{_m>J����_��������Q��o皽n�y����o/�a�..S��KA
ϗ�I-0r�h �����~=Ka߿ĜB ��#�~�ׇ�.x�-�N�� �^�9�Ns�+&9��>�)/ %����.US���Z�xFt'Z{�/�Ʒ�)Q~\��z��XX{pl[?c���\Xw��dw$�~5�Tщ$�:F�w׻-����`��	À����qF~/���W).�P�c{������H	7���M,���!����f��]���P*�+/�����\8@/��m||�RR�c��vw��j0�((��<:��^ȴ�l���k����\Au�Ѣ�B�l~��A�e��]�ǐ(�ӏ\t�v��	�x���6k��$g(�VNZ��Q�v�X��s���<���1GϪ q\V\@�,�>���Q <�[!�����Jhn�`�B.z��h�D�d����: iI���~�/͍߅�X�v���6��;	t���M>)�տ�8�Q�)fG�8�ȝ���	7L��L����Y֥:L�$�f�jTd��ΪC�@2ɘr^A5>J	��5�&��|x�c�K=x�%h�ˎ��kGK����>��m����V�+}E'��[�{��.^�� �Z�?���)�����s�|pĹ�/�:�om������l|�BăD��t�N�勍�(�g�'����J2��0�F}�2��+�[��T�BȪ.�s�����0e���� y��~�4��%��i{/[EP��� %���6mq�.iDmGF>��0%^�2,gn�#������8E�`��ꚃ���Йw�4�̒m���T4�ޕ��++�BY������9����	�`�p�<�{���N�́�/��D��^�_ܑ7�s����Cʷ�ť�;�p]#I
��9��a����Ŀ��l�#D�Q�9�4K����&�Ƕ�r<�r�S��?!��{�{+?g�v���Q���E�~��Y�����R�"S@��('I�f��ﭽt3Y	�p1�C8dV���ez�6��o�E֎�<���0%��-z�*�[�N�]�d��^�.��f����u� ���r�����U�ڧ=�3!����zb��Ei:������U�L/,tV�z#� M��LA�-�]D/|Z��A���>�-�#3a���kw�CL�f[s5X��o��y�*K� }�͍��a�]'�����%�/޼�"CS�Y\��h���+���Γ�o�\]��\��wS5x@ 0圯�Lu�&�=�}+M��{p�X�%�p}C�vF�e�_Z�柗5Lӂ�7���U?Bڰ��� ���mIr��~J�������m(-��
��L�PZx)#�k�Ee�������nc�e޴��o|U Ot�/���'��N&lqNLL�Q����:uW��hc4��������i$�~�=\��v]~;��?tʃ'
�VA�@�����V�܆�l*��V:m�����$�]\����6�ŋW���>IR2�n�!]�^ihJZZ�Ėzhy��BJJ���)g�_~t�@O�Aoqz5�79H�H�n\@c��Ln;��[h�Q��B��N���6���A|����-�FX���d�g�^�����ǹ���@%F�B�O������i��N����;����WCC��	��f��2M<�|M:��)*gOo/�5��������^��{zF<��im�V+T\�	2��:�/�<��2����x���LgOV��aj��i���j��1/~�[xw���M��#�yFF*��}���i���y����X���~P硇� ϣΗ_����nȗ���Q9ݐ�����P*C���=#Ԝᖺ�b(��:� ti�rMٮ�y!�����w�ru�GA�%��݄�c �F��ͻ�º��� 
k��X~QE�}�˰'�I�\��¡�i*�J
�U5c?á�5*?�� T=KN�J����}N1O����ϟ�?,�ߟ����
^__�F����*-]-���5�M���z��jЈy��DsU�����+�������"L����6C;IC����m����5�PpGDX���(I�ۺ��%H6�3�,933��by�|������#t}�H�%�*K�y���`F�D� h�hTH�:�G�K4��ꭄi���5�4?�* �T�Lh^��0��[�ҥR��t��S�?6>zB �9Q�T?e��>@�GXn߬���G���ԫ�LpK䪘r
ss�BkcLz�^��c�E�W�U�W}��*�r��J�W*O���V�}_sxU���󦠚����	Um��@lg�)Q�i\֍�g�T�w�ݍ�/
�ۚ��G�ݬ��bG����j�A�h�W����#����~[n����d��#gf�S]�QrI f��M�ɧc�Q(��13�4���s&�M��0�پ������y��C�C������S�m��@(ɼm��Ӊ�rR������E�����h}�+�z�T��m����[H{��;���P������N?��_-�l�4!�e��t��>��q��U��ZGM���(qQ�V�H�`�_#)��!.M������x�[=|G��5�����uP? p���m�����v*}��a�L��"��w�>�� �C}�ɿ������DaKۥ�=r��t�W0���-{q��=^������kwᣟ�����������L��4�Ob/�6i����ml�Y|[}}aC(-A�Q�>3�9�&��OK��9�Xl^DNK�5�E����1;��k]&U堏_�ؽLt9�7�~��/uMp ��[�C%ȭd��]]���6Q9�~�����:'ЯAиD9��9S���� r�+yg��K�"����R��` ٛ�Y��`Λ�����o^�������3�s����V�>����|&�-�b[J��w�3�˗4���oj<�eDD���V��
���L0�T��'>=?�(%�YU55�2��YYY���$�9��b�rt��5�뺫ղ�(��C�ss��*ɼ�3��h�lC���[3N�e��m1Z�XR�����,m�Ķ�6�A��������8��˛�ƥ�>��$�`l�BB�8�⍥5�I��G9�Q6m�;]��Ћ'h��B���0�������ojg��K���y��n�0]V #�x�����<�j��l��A �=y�3�ѭ�Շ���ɷv�ߖ��hs���٤�����㪟�jl`���u���*;�=z�@���C���:g���FJ`����ŵ���8J����i1ql��-�פ���ؽP�?��m|��##�wԑ�	���������8^݊N�E�94���e1�58�7�G���o�y7j>IL��b��8���x'��g��!8Kz�[�����x4[�e|J� � 
fDO�D1Zp���^ ^��<���Я�?H�bv�1~_o���s�l�XiN�C8\h �\��!�k��hz�TL��v�㚆��X���1�ml�||��C��K+E�zi�*�	���t�>|�M�Љ�ؒ��b#�b[��qȸ�ԃ	R��#Y;?]�Ϭ���9���[�|S8�&_W>��S��o�wOހ��L�����ו��i뮦�l����DE�3��_V>K��Ƈ��e����%({su������t����(�r�2�����o�Zl��cFk��e�Fe2�Q����ݡ/���ޙ��6|�yi_��X�@J��6np� �1�!��0���w��J'�7?����FU�<�������;�����7oG�f&��'Q�n,�����܉��-�3�l#�,vv����32l���h�b�p��ٓʆZ54��e;��N�c���* t���YX��SD0@2w�U��"� �G�h�1 ]������\¸[��w����1�,���/�)�%�d��c��z
Y�J��͇�yK0���2v뭦h��
Z��la�%ȧ2����d�����@�lQ�ޕ}�Ճ��c�6�o?��\��]p$���\;�0��sj%f��gQ�䵵�]NM�ii+f���92��pdOw�Og&E��"BB±%n�.��Υ��Ƶ��~22z3�0���RԠk�@tSX�־�>1'E���/4j�e�I��D�)��w� �ƛ􍩫O�"_��1�ی�V"±��!ׯ�����z��£b|!�&�[�⯰P�o�'�v	�7Ϟ|o�̩��<?��v8����o�WA��c����&���a^���g��̦@��*�`�=R�~�Ƞ"��nC�������*|F^Z��D�B%�ϧ3�6��a��Sų�aq��PPRb�hw��]�������q/�Ȅ4���ޢ{�㰼*J ��77�/��+K��EKH�`��ԣ���>���_͇,����⢐\�$���̬:^P�|=�r�
���\�w:(<]Ōn����@���y��b7�;����L��2��t���䲶���-	��:���У���2������O�J^����ؘ��*�̳ܥ'�`=�r֓�M{U�ӟ$͐8�s�4�&��}��f�<�����	~���S�nA����qK, �g������ $�"�b.���3r�6��5�"Sh)�Q���x���&/�a�!͐�o�R�Mr����K��Z� 픬N���c���K�Ӆ�q���xC���g<"����̥�ޒ�[��S�9�s��,S�D�1>�2	}o¡� .�%G��{~9�r�n�3�hl���U�D�V�������E�$�-QC��H i�
?�4��4�Ӡ+K]�(ח�ڪ�'�崯Y�ig+��h��`���^�E�=sbUus�ȣ�:i�a�0�xv�ܞ$g�ɵ���fa��";{�:.Z{��9��4�Rє��Qe���%$�&\�;���~��^�s�o���8��&������Y���lL9�/y2�����!��
o�
n�����[��/�p�|���V��r}�ґ�Hʾ��hn�u���Wc׾��1�%}+9Z:r����⚠f����tvP�2yc� �k�'i��;f\�P�MZ�h��}��n�({o�A����vTK|�7]v���u�uB��u`���k}*ьP06AHLo`i� m�m�7��C�� ��3�2��Նy�^CfT�z���ң���wtFn��[��&���D,��4�'atfI1��u�QQ?a�_Z�I]$�n�%%$DBBZr		X�DJ@�KZbAJ�;�[Z���<�{�(�ߙ����\3�]W�E_�f��|���ȶD�\ ����n��]�n��Q�v��I���R���!��d������^8��cWQ��ǚ�2sxA����3�E�v��H�m�9+h
E�1i8m"�9v��		؞�Ab��;X��ڕ�CH���3�y�C� ӪB�c|<O����1���ߚ�c̴p�w�}Yo�JC�`j˙�c����1����y��L&�QaJϚ�p/��1���e�z���=}0��3'v�e��m/����R��ba��%��]���&��A��G%7��BE)\ ���ippmK��ԩW��#���ݨ�/w�w%(��}��$&z�Cu�d�{c�!E(�OZ�QK�(!&��a���c�<�oW9�$RTUk_6��̆�kTr�k)K^E+�?�9)����DT?E�*���vo|����R\�E�h̶wm�OZ� �D�Ҙ�;�r�D�!zC�	N��&�mrqޤq����[IK���Ӆv�|�&��As���p�
j�`��9��Հ�7��t�h��[���G�\R�9KMrJ?0찭(�0?���.��;�M ����;<��r&<��)����x�s��G�cy����{��N"�W�=�>CNL$O2c\"���Ӭw-�I:M�W�~�������H7��c���y=1�P���ƾ�g_��gT���d�>O�W�I�߱�O	X�9�� f���>��� �Uv�Pٚq���xWUc#��*���oݞ/_�v��������֯��J@�5�s���<��7o�r��EAFI AAHXX��tK��/�{��c�����'����N�>g{I��1e-�9��JKD]*C��<ٷw�Ҩ]?�|v�]&4��/�q)��%��F���D�Ndg_��Q�B(�͸v湔c��l�V �.,0�n�%�p��ؤO>SP�ǲ2�.��!��+e�� i(5777���ulfi9�~~P�}'����2L���M${�g����(��T.w�����
A�
�Y�v�_�N9���ۀ��۪�~m�"���Q�YO�S��8���k�q8��m<�zG�D�t{�2J&4��D����{���N�6�@ ds�}�B�ψ�♒��1!E{�>���P& ��)�2����Q���Ȯ�%+���4��r�6-�%�1��y?ŉ�2_�޲����h]�)/�X����8�n��(�7�	�wj��5�YJgfga���2�^߳�x@���R	�=��P^U�&�P��H	.]T��k�f����Ƨ`���'Kt�1�`�_�r�m^2d��ߋjW���Pr��w���o��nR�J��.�Z�0���l�F'�;i��Q�K�(�Z*��D���|,$j9􀗊�a�:WF��H�>&��QfJ�#I��H��F��咲�LN�	�4uC��K���%�3y���=c/���pv�5��Jv����@*0�����+�^�l����r�6�N�I���")Ca��/�&��l�p�;Gi�P�W�ء��ѧWZE��5�-l����V�?	�d�7:*�:��n�Z,}L'
`��~AшuRr�YQ�yΕ�$�4����aGk�x�Yb�<�6FsQ���L$��2US0��a���3�Ӕ]��;�|J���ҵ�11�6��ٞ�uU�:/?/���hD#t!��P鿻�[[v�Ҡ'z,��o��t�$V�u��j<�i5�hm�Í��}�ȧ��1�a�]�����C�E��S�����wp��ơ��.H��[yK�Bm_��@mc���mFA�G�ԣ���S��4.X��9��;\��/(e���k�|�~����$����m?�&������K++˷p߮�G����	X���߁����K'����^�Z�'���������%����&��h-�.��~��3�fŶ������E	�y��Ml�`YDI��0�"�I���=�c4��C ��Y��YrE�h�F����w���衪�ji�K
=HՈ���U���.Ԅ��E���Ⱥ-� �e���R�/[		:�~��b�A�h�}��y�Qe���e�Q�`�ޠA	jgJA� �6�3kM����p­��4E'R�&���������bP-OtD��z�̩q�V�\��17Q>�ΐ�_֔�]m�<򩴁�e����+�P��'>������A�U-c�goZ� L������ww}p�d`!�[f,}��G�"Zj���da=�e�K.�/VɅ
]��o545K��ZF��"�e��R��Jn��&|Z�$QkV2)�*�q
D m����DA�".����HH�Q_��5~���QC�u1�q�Ä�9�禦�Kt���U�P����v�gtyyZ�T�ޟ��百~�j�Pw�Au�9����R�`b�������S��L.��B4q[%!����[C�ެ�DV������a�� ������V��a�gZ�ӛ��wH�y{�����Eӷ���q�'Hě��C�-_�k���1z�T�3W
��!XwzS�eC��'Wwp�A�B���Ώ�ص,�媃��zlO>2I����U��W����H"��@Y�Pv�G.xsx� �&�e��qe����C��V��b��4�v2U��$6��fX�ǲ���G�j��S�}2FrF�������|�&��f�4�����]��$�{n���B$��b()�xDד�G�_&�5`�x�� MD0?�D�Pc]r������-�����±7�<���[Z3� �u����{=�����1�S3�,�E�N�"N"u��h�q�Jѡ�\8:x/�F�1>N~�2�T��Di��������d�O(8𿎅���!Q2����{;mÀ��'���-a��ꊞ̒��48�yg1�ț�B�G�}(Ѯ bMJ����Ev�Y�ŢuA$#��/����]����&eT�1x�ٷ�C��u���ͩ~2��sϹB<�윃�߄��������"�i����~�<<mX5�p���p1�N������St�!/��J�ҡ�y�B�ĵN������q��ׯ��ЛƀY(�gs%9茹���}���(�rI	[B�E��||��hA,V;��x����Ϧ�zy��I���5� �-��\Ӷ�A�_!��"d����<�HT+��I?%$�@����L7�@9�v�H-�8F�7+�0�
HJ�q"�Ǣ#r#���[�K�r��wα��[u���xR~��Y|�
��/��4^9;+�~�f+�U���ϒ���MX>�5������D��)�B�whg־gӿ��j����!�Z4���PoD  �.�%�.������㵷�P��9燤���倮��T����8������+�� �.���nynn����6x��*Lr��4���q�C��=��Ȕ�G�/$�+����pp��Eޣ�a�N�ϩ��ٸ*����~̐��"��=�it-�� [b�n�ǙP��es�3��A�[1���y�� ��n*�|I���\zx�=�7��sŊȧ�q�k�M/G�r�1AP��	p�؀��#�f��lC�|��&�g��cJ��kAI�Rܜam�k���t��+��췹��mx���y���H�����Ŭ	4����I+���ti����uw�^AUg�f�Ɔ�������*%���z���)&�<$y��;��a5Ů�i"`��6�p�۷�9&�߼y,8�}x���R����`�V�)@�{���q=�A�9����1~�Cf��3Kp?�lk�t���5���ݴt���ca��g�N��EK�D{�gr�4�Pw�A�L�)�M��D����7��5,>*d��9C$��� �\b�i9�P4��)�!???zgǝ��{Sn.9��#�����dƥvV����m��шU��	����v"���񼘥���T�V ��e�l>:q�X����������8;NU=�v����_z@8��H��B�
u<3C�!���)Sh��w���~�
�	����P5z�?�lY��~{�4�>�a'K��� e �ɩ)&g�啟Ɏ�s/�p�`1
�˷�9+H8:�T�����4���(̴�2�\��bm i]�{$a�GW��}p
��q����3D]�C�o�@�G�����H,�ǯ��sQ
kݱ�N������[�5��"�ìպE��[dq'|�A� ���N��-h�ꄾS�&��$;f{�O�����x��K<��:�~��	��"ɉ}_z�$�� d�@��L�R�����������@Xp�P�wꤪ"_� ��ީ��ʭ�ܡ���R����%)��u���� ��*�#w0��
m`P2 I�5�.d+./�sQ[�k(Zt�b'�m���f >&3�j��x���(��x�j��U��ü����0�qt��$A�ĹR�G �${�4WR}�Έ�gC-T?^����˺�p�|B;٨�vV��Le���>�z����Q�)��&v�����(�'�q�+�ٶ��߻ s��\)>	*�9���Ҿy
�#qO5�fgu�N/�@�2����h�JH��ZT2^!{fgi{�}p���!�pi���A� t���'��	��ǣ/�gR�@,���4Qמ��,7(����`	dc��W��x�,������6e��e$N/>��A�Y��g�B}���]N��
��;Ƹ�^�oǗ�?�[���\%Ʋ�O��y'��a*Ùm�FMNE�<������C��U�&�rƿ��T�(2PY�
�%�~��'�Y�5M={J'����'tx�Y�t~(���1�K��a���!M(�����ɿm�슺:�A�����yh	�h�J�}��E�@g�wS"��q2��1�~�������w�Vm��5:�<��wOMLA��:����}}�f����ڏ�1���QHzz_�`���)^%��-�}-�Gm{OcUa�<:�m~���ڿ-�_l���c�J�L�]�]���0��a�����͹��J�����_��y�?j�F3Kc���ҝ����=̿~���� �L���������ӽ���k��;���I0�f)9���=�P�B42�صG����u¡K�ّe%�,Mu}�u�\y�uC5 �����~D�mM�:`>�/��C2dga%'�h��C�h�T����H�5QL��Ԋ�3�,fh&�kFhH�Q�����|�`�JՔ"	aYB�!���e�NGO�(3�3��H��X���Ã����,�I/u(�H↕���L��;��Z<<W-@�u�o� #j>���q:َ�ۋ�s6�����ϙ�����{6u)�J�b��S/�<i�{"ԗ�2ד�gO�qN!3F�"�gͽ���H�A?�G���z������n�����X���7�f��;CI`��R$!&�}�#��5���,���|����ÿ}A��k��BܠB_K�]J�>���|�Ƅ��+�0����Ƣtܥc/��N���EO�HJJ"7p��=�&T7�0�� `V �Y���ȍ<�o��x������:ߠӜ����F�T�F֐u��Q�г���^
���B��+ߕ��~����6�����%��b�D�O��?<�:n��b_%�����,�da��4����A�2�?�D;�!�"�zN��l���w���e`����!��sX�ݺET�75eLYO]���j�ϩ��C�iF�r�y��Ą�ë*�� rRO�%�q��0���S�D�^^�G/�n�_�\"'�:��Ѻ�Ǒ�W�j��a�Z��c�_��r��Tw�74��چ���e 暰����E��0Gs󜃩���ة�Ci\��ӑ(�D)�q�Ũw�@�����=�;}�vƺ�/�#��LY=G�D;�G^w�տ��zT�2�E��^�Y=@�RlA�X�9m��Bv��mܴ6��^����G�΀�����zc;�_9�}�w�� R��Lsy3?�o���z���2��"����G���{�7�U��G��e�����GJ���7��˦�W�/O~��T<�������53�.�3�ݽ�?7�1�V;i`d�owo|2L�|�&ܮ�gX�5��aYM���]7������*-7� |���Mئ6�κ���Y�� ���������u;�a��n<�鹈0$����$��(#���yP,*&�ے�O$� �OD\\{Tm�VГ��!2&�n��f�)Υ8{e0�G���1��9���U�`]/���*4�Di��B��(=v_����DuX25�-�}~?�w.�*_�t�|���ҿ�^�dT�@[�4�â{#��bLp�0�#ͅ:F�6�2��v�,�@��t�w	�k�HS��_��*���v3�%���r���	fk{;!11���J�j2�e��a-)��<uH�����u�}��ʦY�L��Q>8rG�9�����go5ED��쐅"���So[W�܅$nm.��ٸ����4��w!3�Au�����.i����,:h�khK��z�� ��d��g�Tl���c�^����D������Z�.�A�7*���٩|aC����,3'�j	.��� ��O�SD��0�=E�^GS��=�G���eф�oOt��\��1�>����Ժ���6>>�/�)�x��o�S"���D�����q���G��_�����&&�n�F��NN���T����P�a���
���˓���j�C���J5�i]^F*i
�<֚�H��z+���<~t�\,d	~85�rU�[E�c�I#:�a\ҕ�^���w�S��"��n2���\�H_K.x����Ѯ�꘩uܿ�9x�9ã�1+��j��S|6o�ϲ�]N,��#�6������j5V�hooOQ����sk�TPޟ�rs�'��s���� Ǩ��&T[~t��[�w��[��;��N��4I&1���D�����TUUU�r�T���WL&���h�p2���^)�T����{~e���cCm���^��p�X��ؽc���Be}CP��Av,"U�Ґp�Q��'������j���6��C�Vv��d��f�Ys;�"���q��۹o|�ds�<�Tߥ���M�����6����\�y�9#6��u3�J_�i4�m՜٩�C�t�	\^C(�`z�l"RRq�D����;
���HC���%M�36rr�E%��� @����vya#�PZVF���3;��9�s��LU Cze����X�-l�v:������4�L�j��շj#�N�L�����k��2��X;Kxs0�m�]XmU�8������0�'� p����ё��津�/�f���yI{�qs�~�"���7"�ƾ�fe�t���w���s�@��8�8D�E����ͮ���!�-��$M=NHDt���٨fEM�����Tt��}��	�>'�XQ��N���2��@lni�`��M}p}�rE�g���h7;?��jJg�,2*Jy�1��T�z	�^ѝ� �Xni&S&h�*��^J��O ���J�&����\���r���#7��|Ȍ��w�����`��W�j������4ў���U.?��qV���f���r�O�3��^��g�F�����-�yo��E�j�2�|���Y�����뫢-�O�1G��0��xJ�4�]C�9�~^*�55š�q�4����!�8�\u�cz��N�s��@�pZ�� Z[Ǩp�Ow�1e@s�o��k���oY�-���0-7��ָeR䟷�O��lR��}���տ��j�#8a{|痥���z�21��������U	���/��X�D��"��1�� El��-\�B�����p[S1Z����:����M��DDj�%��p��(�*��X�_�tu)ߥ's��I��:���[2Sf\ƒ1@������Y������\�#@M//ԇg�^0f����9dM��xT_|�hf�9'����,�K�p�jX�ƀ�����h�5�tD p��V�ɟ�6ǲK}y�Z��튴P�=�\
�_�|����8N�ԌI�
Z	����}'P���O�p<����RDտ�l�s�_=�9��s�����ί�_��u'Ya��c�I�Kc�@��f�5�@�(��x0��@n(���E٢
�t�ڟ�Ϸ����-�m���PZ|�2f�^A���H�DH�\-�
}�T���o�){�sc�=�(S��mtV�@�YEAA�|�z��S�k�ȶPw!%֥��Ԗ?��^�F�X
�JH���
�!���rk�:�OL|�HR��ud���+2�y���Ge���&'��hL$��E�x��%ڊ�xE_� =�Ϸ��Iwpa��dnnn%��瑸8^b��be�8ii�QMǋ3#��h��xO^mb�����7�P�q"x�{!3���b��ͱc��2<Y���մ���ӻ��Z "����p��_� ž��-���}�֌,*��G��Qn����j#�u��ȕXy4�:�08��9�BL��#q7���)�@mt��zBh���89V��E�P�6�[�4g�kޡ����U�z�v\����%��j�7ul�ʇ�{�:NN�5K���_\x/��o7V�Q��#ub��Qb��e`�X_O*��ulfcs�q�i��ti�2�䕵���������d������3C�Q2yP�O����Ԃ[���s�٩;�*�0�G��������-�;dƜ��bn�d9 v�pg;���n��e�6R7�r}�'M�Z��"�VqIު�A|pi �X�ծ%dsj󌎮��c�TAO0��\��5��w��Y�n�$2���m��>\�-R9��s8U,�3�5x���lh�:�O��HJJ�E��Λ�N�MM5�Z�GA��J��r�m�}�������-,`��ᬭ��F�˝��.�ONO�TA�~��upV����-�y�a����=�+d�P c [�|�a��꺲�6��R�:C�$$����#��C	�� �OH޾v5���Y�Q��sE��ﯭ&�g���V(t������vS�0�(�f$ԌpPr.*+�~Ґ�s�����;9Ik�#E��~��
�S�"]�]ABd+��g�sk��)h����[��)J�aSS/l��5�fjˆ�(�����iiiI�u8_301=�D@c�He�������S�G�X���Y\�~J�Pg/��oQ�,ꖌ���u�R
��N[aDd&t^PAJUX6��(�� ��a-@>p�_{C���$�)�C� �����t��n��&�Ǻ�����	*���b���ʵ,�K�[Ā�lC^���=wuq!7.��Td�*�88�y)��f�����f�-l���!�n!�伀����o/�yh,-'��&dJ�������mG�T11�Q5G::���}�O2��!AXR�#06���	�O�x�H�_�EQ����Z�NVl�����]���u}C6��hQ�aD�tC�
ACk(KSk�-XN��P�X%8����ǖ��ƕ%D)d��ʶ
|�2�痒"�),`��E>n���&M6��y�!wWm����=T٨߽����(ё}�C��z����^��5��w,����F��^�
��s����j.
�J��D�٥�f�=&���!{���h�4�`��^���#V��.\��H�h��dB 2�V�'l)�i='���sm�� �5HK�4�@.oe`���m�o肧9��r�R��3�qK6�mŖL�;�����I�r�<˶Q�t���F�����*79HyUU���嘝��F�A�'��Wԥ��i�`9}kK�_E���$D3K��|gbb��$�;H�⑈"66��_�پ���"6ddd�}���� :7�)�	�diPto�+����<��2��;�J�
�Z�!����zC;5$/������~4�}��?�/KCK/��;_�u𔑬0��U����5���(�����{F@$u'5������#��86�sGl>��7����qz.X�W5�B�vxH�tA��à�Ya&i_���t�7���5�l6�yÓ�<�v�z�0ӆ���:���ۻ@��P/! @��8L./f�u;��ʂ��Φ)4���������mRfd���:p߭�^;<|�V�b������\��O���������� upʌuf�yVC��[�5
�#J��(ɍW>o���~!�<<�) Y�<���S{ֈ�����W'�2�P�K�w@ɺ������Gk��2..�YJ���Dj(�>!aw3P�&��^�.#L_Зڜ	"�����GrS�O,�D���H�J���x��-7��#�;7==�S����P���uC:��=Bxt.�%qɽRD@�{VzG�3���n�U�����0���?;���ǘ��PĴ�;�k�{"��_�=�P�걨,��<e�B��H*p�#��0�&7ϧ''c|���k)����И�w�����閉��-��H(ѝ��j�*O�9�l���sC}��Y>ŝ��2�P� ��Eo�X��,�w�Ar\	Ǩ��n�P��n�����#�{'�q�i
x�"�kw���Po9Ц�;w�p�C�h3�(��}����ZL۽="p��>�u��ֹt�Q���o�[X���=6�]���X�[vYC�usL��L#Ξ���<I�;A<�<�Ȋ��A.-�K�C���L��Ծ/r�1���lz_�����ϟ���>T��K�7z��qH|����"ןZ��JJ��U ��JHg��}V6�����֩{�S@m����{[�l�!�lP��PQ1sV�ꈀg�z��gB��Tb�a݈�n�����Qc��S(f��8���RH� ��%��G�zL4� ��篁� �J�<�;���좦�ݷ���]�Aev)�CC����</�����W���'''9(V����O,U�ʝ�"�W�ܖ((�Ѹ�:=gaa�?��:6��sZ�zX1ݝ�{��o����Q�YQ� ����Y�4�B-@�.���rP��OF��L�E{2��+�	B:�. ����2��6f��L��z=�>I��,I�~��=8a #�ũ,�}fu��Qir񰶾��ݻ����+.w�?��o���:��G��Ȉo'�.�a�d�%�T� ��T�`kKg\�+^����)E���ghXL�g"mȐhHw��7o����w��[��LMɖ�>${'���U"*�x�����K��9<:��)���m;+���(��)i��p�����(��M�f�>ًv�xs���H�!��`f�`F�E��\U��>�--v4obz,���w�I�����Ñc������p���{�(J�c��G���-}C�[\m�Z��f��H-�[I�"�gf�il�>V��uϰ�Bs�33X�RsS�!Ob����gi�N\\��c��b8:���ݔ=����͹5�6O-�8$���/�cьw/������<�KNa{X�-��8�s%h �Z���E*b�>�b-h�R�W�*�fd+�g�H���n���G���H��������|t��!��5L4�B���dRVT�W�KZ<��a1�4� Ղ��<��@R-��b��(�g�|��</�fo_̯������o�wx���7���Ŝ��}� {���K�ȧP�a�H���A������]02�
��˶�R� ~Ä���9.���F�d<�q�) ~�;�DJ>"t��lc�G�Y�o������1�@�
������?I�T		������{����mݷZi������f���	��p��
!!!�z(Ԇ�~~��o��G8J��4����q���D�%<����L*f�r�8������&�����v�5��iL�y��W�)�F^b@|����z�7HMҩ��W�Z;<�j�`�%~s]��{���Jc������.��c4BG�ȿE�k_*Xw�J2.6Is|�k�؋<�3-��̎.�]ў��v�����.>����ohBh�k�[Y�<%FtE��3��{�CJg��Ԃ���o��ǫ�+�؟�y�AtW �F����M|^ޙ��SS7��#��Ǿ��� v#3����Kߖ#���2��^&�%����^�2k�>!��`r�Y2����i�������[U$92X%�\�j
ME@���80�kWHX��W&��kݽ�¼��_ī�d��Ū��B"Y$Ϊ���d8��AE?�'�X��"�,�~��goo�4�#��),	�����M��}��<o��Ѕ�/i_��YL�����.3iQ��z6xǨ���?��-5ukx�d�XNN��'Hp>=l�ސvp �,xm���>(��e��f��d8�PYu���c�6�x�:R��y7}��±E ���������נ�5k�ڋ�ZE�p�=���Q�,��8���p���1U�YJ͌�L����w3�PbW�����k��«ޕ�\�h&����O�&�K����0b/t��o�QeiCYƮr��j��;��d���}�&��u��7�^�iq�o���,�)���_N������g�E_��W�b�$�I��ژ��m���&S��|I�uX��l���� \YˬB���]r�!7<�D��ǊL��(T�~��[��Ɛ�ɵ��(�&���S�J�nn����o��>�{�:-���U~{�ny�^������m�XTT���/��Sy4:���Ξi*�=,�^<�:/���'�H�������6��ϮAv;��?�0ߨ�.go�yV4V�|%��x����}q1��-A��@����bח��ß��,h�J����뇷���kƏ�a8@��2H~�(U蓪[�-0�=�H��!�������Œj�-52��Q�`��[��Xpz��F��v�6Y�
�6�ф��,[O�g���i��B%^����-�N��wBd����X��y�<�wW�� {V��nDV麘m�q�5nM�Ϧ-Z�$����s�<⑨V�6O�%9jr&P�&ED�7.�VWq�"��G�gml�@m���ojo����b�:�FB����ԁ>{��'����o�*�(m�K4!�q���d�+ό��>�7�~��9f�^Y�P�?g1`�Xg�% ���߲5TL�-s�9�E*��rx�Z�LTJ��7���%:ߙ��%J�}y�`q��u�kSS2&�|?�l������
J�ͽӥ��5�z
`���`�:6>5, Zξ<���PN"��(�g��Y╹6ä�C����&P�\�&�,�'&&-��#3;�
�G�rF8^_�O�V����^��=�X֥k�dC5|@5��g�EPU`�~�p����6�~���D��m-����F����j	/�DK�Y�kd�l��QV�gy��T�*w����Y�~-g��Li'(�E��U�Ը6<�ss���������U�w�
/dM٫�5�M+�/�?z�.�t������3j �]E����^�N[���d���!��\�.������&�+22��a�V��"־o��'>�a��D�<`M���cA�&?�I�-���jH�Iy��A1��0��,)��mSH��J�/���<b��Ukb�(<���~��̷�w�xw���`9:l���1hWFmʡs:05���׵e6tlll�&R�D ��[�H�Dr���V���F�����ӄ�.���Mhg��PR��?L�e#���Pj����{�j�e-�b��V�������3��1��'�
9���=���\����A��[PDw�4�$���ݼu~��i��my>��͙1�~),/SoH�.h���tf��� S�
��s���b�(יl4��$%T�Ы9�Ǹ�@���G�x`fַ�C:��Wmk�½4����S��|�K��/g������!�X6s����L�
C���Iy��naӢu�	���p����ŰB�~n��PH��dU�g�5&[����?�2jy����6V� �_S�9�&��&Jt�v��Hb���C�f����V�C�>j����p��"��/҅sD�޻kY'�19LH)_�}������bJ;\�]"g���-��j�]���!KYYni���]d*n���c�(�w�����-˿}���nm��K��E ���Rq�y���}j*=��{}P��] ����Ĳ��û�s<6Nf����[��E��-Ȟ�e����R&�H�%�}���>̀ ���c�N�޻���[Yy�ߦF"�@$���1^Q���wf{l��zy�Z�	�N��2cj�~�%�r��Llu..~Cذa��=@�:CE�M���ٸuJ���[y�!�`��+�|^NN����aY��Þ�cçD-�V��w�� �}(렙@Y����Z�ų����u�v"��u��->�gu���
dj?�ɉ����r��9ƞ���~���[T$���zà�(��S_��tsy�n�7D��q����o9�����T�>����Pr@���X1ȆN�E��0���M�PyJ���_��p������/�ܭ�P����IrR/c;��09$c*�&��w���)�Ԗ�('%>ж������{�������\��:F��[�r7�$�P��o�/���O��9 W\̝2�y�U�Q;�x�j�nP:J�IH,�`��/T=^�wp��uμJt�D��
�������{<R-$j��*�*����,�*b��N�B�������HYh3z ֐��)�ƵϤ h5�����A��Ik�Q����e0�3���(�""8$�I���1�����I���O&������s��힟/="
���}�����d��'��&��2�3G�f�0����s;�ԉ�"
2�4�ƀ���Tt�K0����1S�1qҍ�=��r�Łv)���O>����&��66V���C�e�nP7gޕb^�	�'���J���IDF�fs83ֿ�x�&�7d�W���~3Y᧞�=��n�('}S�f�h�	7<�Ƭۈ��H�P�gx�c�Y}_�j֜]�(����cA2"pp}%��͔12����
ä���d{q����HT"]*���[N���w@r����1st���[���NJ��㶵���w�(�O�A�:?��U6N� ��|Tc�S zǈ�|�J�!Y�zidA�[9����.�:��i����C���!a� ��b���^���=k�nQ{������J�s
Yḵ����8Vm93�P��{���"�s�wN]���)I����������6I�x������*�r)���&���ܜQ�����ty�j�`m�#����9��/}��NO�+�]��/q��7,/��v!�v?��Ս�%���vpP�����\@�x/
�Q쳖�z��*�Ez�* ��YX�F�d�ۀg�E#-,0<,�030w����a�,!�}\I�4ᵶz�Ū�`�Vʉ������bh$�О�
�_Y�42������+�q&�i(����_Mv�9(�F����mU��}Ͱ���ۃ�G���V(m�ti��� P��!h\�:IojlD:]0~!E���:n�N�a�����I������8�z�A���>��#�������c�%ķ�����_�m]�}����p�;!�f�#S�u`:f	�����$�Ps'������د��F~b�a|�-��Qm5[j)/�p㖿�Hc4`Y3�1���F�iio6d�~����M!��l�-��s�}9���c3́%Aei�Q������5Z�a�ݯ�㥩*���S��SSߪB���24�G�r_�[jk���I�dƠ��"2��1���{���n�'��|�Y�MSG��jo==6@J���Sc�M��7f:���MG)�B�v��a�Z�K���׺�z�q)X�`�`�1�-[6��o���=�Z�+ s3Z\�rKOO�_2eF_Ǿ�;��G���O�.�"��Ǌ�a�,�s���*[ ;��j���|��4uv���D���4�q01$�O��xđ0+oi�r�%�|vky�b�����sZ�:����}����KY^lH|�6��&&��`�FCTl,��g�����YC���zC]�$�y�Q���l�����-��H�u���`U�����+�����o�4"��6@�������k@��$M�}.�����]=�z���𜵵G�=�R��2��Q��B��[ e_XJ�bAcctoo5`qqE璌�"�����G�u�<O����HP��d�.���g�mlp�rßqS.�_qy��p��l��ݻw��-
u�k蘍��oP����۰�����L���I���F��� ��1������CX9�~�xP6�B9tSJ��i��rI&�l�6Ǣ��>�4>��O@MQ�AsRs�u���8�8�s3O�
�{�=������Z����w�� [�ҴGɮb���t8��_�<���C�����~�nm�e���z���Xq��@[�A�'50@4`ř��ϳ}���%���C����v�]�2,H�mo;y5r�남��9�ԝ��sQ��iV��'#�R�"�*����.��X��i-�AFjI?�z�o�ߙ����
l�J
w���5c�e��>�7��n B�Ʋ*Ԑ��U�{�J��/��{����BB��Ռl�%i�*�)zn���}�
�~]���ORj��(՜.Ob�L��}�^�]JpggHRJ�.��5�B;*���6"��p���9������U^���S�r��(��	4�"I��k�q�!q����bs~Y����)�B�6�xꀥ��C�u}`Q�'�m�0;�-� 8��]&�[�S��P�x�nR�{��:�� d�Ø���)n�ܸrK�0�o���ss�6s����;�s����C��h�W��0Y�QbvvQ��ႉ��k)iiHd���=�&}_?AB,;�"��8|�l�[ظ|��J D���|������-���9#uG��ffO^h5�;(
5��^�W�����Ĥ�P�N�k۳j5Rp���z?����;�� �6P.�s���5�-��8e�}����xJ?�ǁB��#�6�g\�q�!"b?+ ������S��x@����%/}n�M}a�9<��9���`�6���~X"3�iJ<�|D���������I��	K���읚𑍎���j�sߵ8�]]�Rɭ���X�]\\|���a ���$�넪��S��z��/(�jY��|��C�`s�����&؛E�����=A�D�*��}�"���ރf�v��%�:|����Q��QQ>��0 %��t��Hw�,��! )Hwww����,�%%�������+ҝ>s��s~���⸰3s�ꚙ���*��8�&�y��{�y��s\\O�6�������1����j�����e����0�x}�����*I�۞uNd�ሇ�w��W]�[���E�|�+Ra��G�iL����-�.S�1���:��8��+��:��������K�3����"/���+��}���^qo�~|��X�}NsɝڵYՈMz�mN�K�m�����tW�B���@H�c%��"n߾psY�qޙ�$GF��C���`��]n�wv���7@��
��Z�7jǿ�Dx���ׯoQO�-��[��� �R
�����1�p'L����ZZX��O/��r��5= �J|!�7�팋��+��_�� >~=�K�K]O�ymȞ�Z=��E~I��e���Q�7��ygg�s�7�888�E�q��u��}9��_��dC@D��*-M�<��0� X&�zC��jO�e�80��i2�����H�߮�#Uw)2�{b91V�c	��^ ՟rQ��*������Η_HT�Z�6�;��ݝӼo�;�v����o^w����PQ9a����(
�}wP1�T&�
+*j9n:,2� �RsfR|�
�W�O~��3鼕<�`i���`���KY���Ip����c��������Ze�����I/�V�z��WdB<�,�6��(̛�b�w
�����cE�	��1AЇ����:le�p�����TRq����F��跉ec�;�F�1��������o�b���Љ��m�f�D���Y�����ֹA��(����yN�|�53q�e>�͈�s:��iЋ�x�'������	WW������A���G�D�L`#Ƹ�(t�@x��S"�uV�+�����1��H��j�&�@F)Ϟ]��*�B�I�%;O=�H� �c�H�Nc3�|?x#>�75����	+�
�d!|�ǂ�����?���;R��r�E����,��g9x�hV~��002����5R�lU���2�C������� �C�:��ŷ�[�t��I�С"�\n>�`d����@Nl\��~=0��������70z���	�ۓڕ�/���mm��{Pcٿ�����&��\Rbj������6��G�b�� X;����m^dވ�y�ų%Z��cu#�d��x��v�M��������^���m�s���d�kJH��3Ux&��,{�~�=�����rdك�痡�@[�T@ۛ�.;j��9������趋}@��q���WH���ncj���t���"��vh-+k���-e*#��а�����?�XY|
�h�t~�� 
�"�����l�b1��"Ɨ6���f��m��%�\�U�ŵ�4HY��������u�5�t6a+��o�j��b�;����ȝB�X����'< C^��N�§������p�^����w������W��7	
B�t�<��w�~��_G����̜ǭrh.d������$b�#(�:��ũ�3������!�����:T�(rپzl�����؈T�U�MF���`GEv�����冷iS�s>z<ݥ���v�×�6����=Iu��do��K����h��P��y���hu�`0o*�kn"Z��Ǚ/���	������'ѹ�|v�wT[,�*%���5�"� ry
��>�(3 '&2m]]��p�vMLp�D6n}�R��k+zя=��r��xe"?-5u7`�����mͣE4j-����6�ijn��E�^	�U(��96�NL.`.Ҹs*!�c>ξ_�@H�-ͿΥ�rs������%555�D���k�{���]w�=�i��B�0FX�>D���f��hb�ͅzyLR�l�=���Y��p�'ė���Η�|�Cߵ��>�����Ed�ںF���Y�{Δ�,3�)����#�wAM����Z�Р���^��ii�z��������mA�I�I?���}��n�~F;�8�ba!�/���{�ϯ��x��v_�+�nb9��GD/�w�,~i��X;8(�N�hTUW{�����&�x�����|YȽ�w~?AP�%r�rE����б%�"1�ھ|���] *�1kZgD���~,OE�0�}�l��C�g����~V���=���&��N��hK�LhK�5�<��.u:��KD�HS��)�"��oW]�����4;�dI�|�R7U���z�֔�:$��dm���ǏX+��f�<��~���ܒ�e@ 9y���
 C�X�������_����� 4�y��dNd���u����{�۔���s?�-�A�����Ò��yv���������v���cz��O��fr���f����^K��k���)��2������$���p�Õ��4�IW^���W�	&	��7��g6$��­���]'��m*3${���//C斗�Bca�����>����Eo�l�P�|q�ւ5���:J, D�R��w]�u����ggPg�чJm��������8���)�ôFl$$��ղ�ˡ�Q"uMM�elXᅅ,�ĉ��}+}�C-�HA�qS��qHk���Ņev�� Y�3�bVNL��⼕Y�3+|�?��~52ӫȷ�{k�L��lJ���8Ą������_=I�x����0a[��.U�{3������\���-����PfH�H@SK���f|O�Fsy�h�FUMG��v�(������w2�|Y�!}�O<=�
�KQ����@꣓f�&"&~jn��Ǝ+MEU��w�d�$edꌴ��avT��@g��߀o(*%�|y 2F'FKCV������IDH�Ch�+�=����𹶨g�b���.Y��3��}��q�?M��|�u[�y>Ҋ����N��<�(���	����e�������,@4�
X��	
�:���ǣ"g�[������K�����XU�0Hs�'����x�,oim=�w۬s!�����'�/?� ���_��.��1��%�y�%)yiy_�e��aY5'������a+��:w�Wll,do�9Ҳbt�>�R� /���G�����/��L��$JJ˼���A�gV׮-�=��-��^�.����~�&�� k��K����7�r2q',���[F�'8&~�_V��[^�C�dk �|���e�Lg1���;�Gw)��v��"��9���==#��nWyHп�I��f?6����H*����)_&�������#��O��?AY�:���+~֘�vD�݊��O(�����)CCFĦ�'q�	�ܻ뉰\M�9o}����.�������)I��x\�n���];�(j#����U�R����Q,狭d���ֳ�������s�C���;��v˥F��8Cq���	:���DuWv��;ᨯM*0o/C⡧w��?��Ȅ�T]�U�	l�z��%��'���\\\���%UkDe�{��&�0ɩm @�#�ĩ�<JK>궎��i���S_��s���S�hδ��1�F��2+���dm��PVc�t�l^>���<	��C�È՛j����ن?*�����{p�-�9=�Gؚ�v��e��++lm��G"�YUĞ�Ƈ�6?�
u=:$a��
#�ĭV8�B�ry�C)$0�龮���`�����V;k}�o̪�����w9�R������lh�i 2i�ث{��*F�/.f��� S�P�
�w�y�V��b�[��������H4���.�y�H/$�3}+���k�30].����Ε�����נ]����{����z�8X����l`���tTҜ���3�b����%?���@��f)Xb����? �#���yh֪s����$��=э�[��~�`	dO����q���'�d1���Q"�=/�~����d�a���uT>�1��	 �9������:�Ur��;qp|l��	��--�^�f#�����[�hSp!˄�7�'�.|��hl:"X��fb��P���Z��&Gk����(�� Sf���
��-���g��d�!!1��1!~�����R��u�W��֞��1S�얠�t�M���d��M�Y�p$��Ry�#�"��j6�P;wF;"N�Q�&���`��.楫&�遊�m�#'#�9IB��fǖ��[��#�/!��QmR�=_�ɕ8<��R2��M%�Ð�lEmdf��n�9��#� �%L�/�!�ZŠ�7���e���$�Q��a��ddf�%  �������{����=_�I���I�x/�����8��3o�æL,6����+���
1YY��v��<y�����.��u�g�=v/���KXh('�ꪛ�fm������W{�#�mZ��阙'N ^�^0���o+�>A�p�q�/�62�Xh���WM��R;��:ڶ�Y�n����NM��@����Tѭג�,�~��Ti�}!z�`p}{-���9Osi��Xz�?Yii�{wщ��0S>�&5�D�ļ�"��?P�W�8ݥV�r�g=?<<4>��ZBp"�G�B(`d� $q�_9�@|z�I�v]�E�ynz�I����؜���ٜ�+��k�}
�!���Ǚ�0/0����m��6����`%���qP� #�B���4��� �0�<�	Bb�=�©��o���Q�0-�4�����>��7��M�ŉ/;����1���mϬ ��WI���o2>�q�K��ɪD[�o��������d}����݌�JLL,i�@���'޵}�#�Y�������������zK|覫�����Eж��d'|%���)&\���dA�U�'�83a	;r5��Iʇ��Ȑ��1���lП*��rH�橵+�xP�bc���-��ٯ_�y����wŷ���>7�61<���h=�J�������� �dȨ�ػ�3���?� �>��Y�~�CL/�a�$N�|�i7V���GE��SS�����#�ohj�C��Q2cA��J\�Ѯ��']Y���w"��L��eX��=*E����/��*%��͝�����˗���|����-,��#����^1�mE�>�"��@|Q{h���#@�>h���.)-+�7��|����0o4bO�y__��49S�t�&(����
2'������QT}�� G�_���eI�������J��o��۫���.1>\nmͰ��mE;���;=]���!}�)�1{vХ2�k��~���pC�����O�:�}_On��V�'H@Q�jAs��9t��B��Ԉ�O���_���������"��>^��a��_����e��z�
oi�v�R�rM�VM0��*�kYOwoo��svZ��:����9A����#g��r�VV�,�?�Rc�Gs&(��`T��?��J�Лiq��tO��}�����Vi�y͆m��-t��Z��PR2v�z^��k?{F|��DDB� N���+�� =}���7�,����o�Y��Mo�R�~_��_׻�~��8�`�!/�z����OS���2��<5�3��8��z�$�ܰR��9{i��Ü�2�a�gK����d�6��Z�Q�Q�UGp+�#$Kޞ�.�e�Ff!Q�zr�A�����j����1/��S��ՕQ+_&fv��NXNe�8��$u����#�Y�P5���^����>�<Ɂ.n4sQ�,1�rRXC��:�cbrA���^�Cvp`��;9_&��9P�}��;y�Ԅ/���,�#5�w?8<���p����%���~]ږ�_?�h�IB�`b��e��i5=�'�
O��k6rݫ��翺��5ƌ�49?�｜<��^$"���$�Ǐ_]�Al~w��Z��-B�1|� G>��>�&\����^�'�6h������Z_�*o�/#�7�����0VU�D ��O���,��S|d�ӗ�-��w�EA �PRQy���l���+���Z�ww=�[%2�G`��@���$�#�͆��{�1f�jv����σ� f���l��	��8h~�������W���5`他B��I��O��i�����!����=��L���(��v�Ŕ�/ŃMe�_�.	�JW_����:.ٔ�
�wk���׊�S�JEEȇ���u�u?��ؑ��.�{�K�/��"�&!'�;z�X:e9�j�����
��+<�IAaa�*������i11�*I�a/��-�ϭ��;��t�ﭜ���t��j�s*WCg��*C��x��X���Fv�����XV�16��[o�_]�4��Q���Ȓ:����_o�q���-�utxx�EL�y��[ޡ��۶���ᘥ�/ֽnv���P�w����5������^��2w:��H�4����(zt��A*#����iq�>yW��n���%���/!�����P��v��3_���jW�S�|k{RGmʷ���OA�tR���d�UU�� O�Y��_�nRi�?$b��ikߌ'��g�V��辽L��MD�O��N��qS9����U�[���k�f�پi.��y��<3�Wq&O��\ڷBo�UL���[<8B'��s��-Б#o��X<̶n�t;˻����FG
0z*��k���X8ן�����0a���Ne�iAp���i�g�k�uz?�\�D����z���Ȓ;s�X~������h)������[N7�	!�2�3��ٔG��u�K��+5��۴_"�����|q��'Yn#cq��h���9�&�<��۶,�r�_��`Z�c��e}��~oo{�o]c�g��Ǥ�'�09�-��_�XA����;��q�����C�����.C������#�i�_�n$§h	q�x��N�Y�C��ε�U
�5�-&�C��o%fd��+���95t�,���C��NEm/�>���}��ݺӆㇶ	�`Fj�ɺ��8�Z;Z:|캖�,��܁U���T�Z:�K�1tOmO�GJ�^ּ�v�6ō,��5:\�g7�;�T�/�e�++��]`t)*SssV�k��X�}���Ԅ;��	�4�T^^^Ō���II^�*��-c��"@��ו�M��,0d�3���42d)T��vy��F��)?��S.8���8�v�iX
�|u�m�ǚ�ƭ��C�*�-πmQ���p=�u���}��N�}���l�X�߿��<��yI���Q`������pcjB\�㭠�B�I�+�Ծ(���ۆ�&����ɐ�}�'㵡Q�����SW�%/��;����umE��m��^8�8Lͅ��(q�mk����N�.��4���ɉ���Ӗ��[�LII�۷�i
�x�^�gO�L�M�;���7]$�w{%�GPay�v�S���F���I02��@O�.�X�Q�#E�[m���r��\OuUA�����Ɗ��������4ˁ�U*/���bk=�]�sPz6��io/Q�:���R����8;�#"Y�_�6T'W�E�?$Ŷzpr4��p��ZTzv����un��G�v�򜁞!$�$�"st����3�4)b�#��XI>��&�����=�dqi���������P�{(Ԉ���Ü�5%fR��~��$Ԧڋ���{,$9�s⯢'7V��aK�_ZKfƟ�9ã,LpP�Z��\��Ɯ����&/ػ����B��OW��n�UVpwK�&�a�ݽ{7�R��%Tij�ǃL��1�Lx��+MIONL�&��|I�-�v^n۾�:��Q,'z:ha��2K�S_(�sm�%]4b��Ҵ�����\�@�s!us3�������J�&� ��ޖBG{K9k}��VAߊ��x2�8���>�S��!1��XS>'�}+W���\;�
ޏm5d�{���(z�1�9� 
���@�<gG��e�9��L�8�%��$��#�k5ߓ+6�aJ�[:<���		z�& +Re�� {�W虘4H�X:9��L�{��RUe�y��-�Ք�����\��d�,��l6wv�����H8f'���wp꒻@��Pe��@YdH��)M����|�(��J<
���(�0�ş���*LJV��jr�uVzw L[��o���
(�Qm�m⢃���l�]�e�ӝ(��n>p<4�ʻ���N��C8r}j�>�Aqn���a��g�՛�@�� ���%w���pVn����1������n利�?M���+�sU�PF�9�df�M)4��S�J���ȽŴ%6d� >�y���y�V#C8�.�%`�ݥ�&vf��ꠧ�LFkA;q��������MϠ1�n����3l+�\��-!yj�cx`�ɒt$�����DCs�� ������
ۼ�VRߊ`�Vn~�J)�=��z �''|��P��'�zm.���އ�'r	�$�k��/Eғ�i��|��Ԛ5@M�s��Y�i��=[lZ����(�_���㝜�N���i�Q��^c9�8�>X�9Ig�j�uQ4yP�$
j�ZX������z�$�yz��p<�o7�X�����+��kE����Bs��S����\+o��#�Ѕ������gdİ������軷� G$��Vu��x���d3���4�6%&����B��oL��$B��!��R�:az� L`�l�q�L�8��gr|�a"����B�	}����or���Ń�^��E%Q>UJ�2gء�]+9�C�����!���OdI��^��������B�q�x~�S�����]g���9W��W�Č3 vAdr�9�~�(CX2 ��[�x��9��0_`�:�J(mT�Alָ���xr?�gkce�)W���Q���n��Ut��ɟ-���$���p�Z�_C�w ~-8{���ϥ8W��7�(�Zh]�5h��s��u�6L�����ʍo�6���^QR�ԭ�����W�r��L���$ʏ)*")�|���911T:�v��n>mǈ!AO�1`��oN������H$^ٯ�DLJJʝ��L����X9�`*���-.�[�q���a��`�m��i�
�c�?�*����/��D����6�ʰ���qF]]��#�W�|t$�oФؘw�Vr�HijI���v�{K��O9h�����6�&K�k��o_�npa�d�I4��j.���y�)�AoR]�Ph�݃^BيY�g�������=�S^.���&.���(S��{�u�l�w޵�E}z�F��ٲ�k�N텳�����Z�w7��,�7��$Y\$nT%�3�����	rG��wg:ն�����ǹ���5^R�2`T���ٿ˹�Gq�.\d�W/������,��Y'	����(�����|��f#���($�+z��I'���=c��|����s0��	nE����1�C� t��ȓ����r%�@���E��qKܜLK\���C�y**a�����U��/nmz�>,�Cz���k���Y[_�w�x� ����15qJ���5 ]7���O��.�껺bT)B��Nl.Ϻ�E�HYY�t(���;/Vk�c]�K�3�.��:��M�[,(�?��p���[h�9�HT)22���e``�r݆��?��+>wp� z}X����iq�^}ش��h^� �×� )�j��s���X�X���"�]74r����m�T�=X"���ź�O�����m�g�������C,x�k�\��$����Ms�h�ۂ���t��ܰ�[c�PL9<�65?ˌpL��b��o�	#╿�ʹ�a��E?;��)�,;Ҟ����2 `���#t	6�XUB�r�|���e�v�h���JQ���Z/��+��
A2J�����,�{� A�!_k�աuw����T�C�_b**�^I�$�����m��a��E}�D��ׇ�R��8P��pvu���C�5`�4P"y�'�+��A2�?<%�iI����Y��Q'h^�7�<��gfEX����C8׽�2}>ޡ��ʑj�Z'�ӑ�]��v!
m��f��^V9�����F��M_��{/���� R�lRbE0�\���R��^$ҵy��N��67���罽��L
��ϻ������뻏�b��W��B��N�sv>�z��-�5��vQ��ܹz�C�׮��"黦&�)wz��%��Y�@�)렐��8�
�>A�LgX�$~���~�s�}ޤ�ö�~���/o��U�s�r����T�#֒�l�JTc�	�����'�*��k�J|.����G����Ax~I�n�m�׽��u���OU��@���3���t��u]�G�<ԝu�Ŗ�{�;b�p)ǭ���ۢ�Ti:3���� �����]r��+���xxT�C�s4�Ss$�K(�8A�ڳgĜ3{0T��S�v���))�KF����N;<In/� �9h�(~��ߠ%FdA�\'GM(g��|/0��	�Y�5�7�f����n�����Y�)eQ�.����+ƪ7\�ZZpl��We�a�)���� ri��|!���h���/�����T&y�v�z!�O���&ݟ`������32�U_�Sg�;�cc�X�I��x���P��E�����mY��$������3*�5���`��J<��T�W�� G�Ǳ�h�_�n;!ȌYҍ���tTJ���D׎t�UNn4��ކ߭��
���ӹ�y��;������o�h����ᑥ����P�B*;�(�����n\o%֡ #|V`��t�=rӗw�9�i�V$8�yT'�YJ>�יN3
��&���\z���؍���\�5��X�Y���V��(�܈���̥%�q�">6iO�EjkZxE�}�q�L��P�ߢC�5M ��L���-s�	��<M��4cJ���˧�T�=?=�ssݵW�n�ߜ���E��n�<���[�k0��a���^�4+P\��jhz�Ʊ)��R5vG��PϽ�s|T��[�����vy�Q�Y����;�+~�)Cs&��7�g?/q���N�O6l�<�̚�3hmmc�s`�Ά���X� �L�S�G&œ��o�ί}Y��I.������\p��"����ܦ�
.�vh2��`��=�$�D��}͠rV��B���� G�HD�ƞl^�7��
Z���������@�v��'u_6~If���u�M���Ǔ0�=�dk�?AFGd��qm��������"�ڥ�5r ��ÛLهa�**$d�C��V4,_>�]��p�=��-��lNY(+�-	�֝���6f|6e�����;G�|�{��٧���?�~�ntӷH���ō�l��O�,���)u���M&�%ni��$#$ͳ�b*O�[9^����v3!�B�:~�g^d0B�~���ntX'p%�MJֹ��W$z�$�w.��l���$��� ��@��I�Xr��u�L����i�����X櫻D��.�\�Y<`�Bt������.v/����Y
w+�J�}��jK��X��������hv��E}%��2�|*l���Y�1��ϯ]nj���b�u!�ܑ�ud����:1L�����.w[@ظQ��&��#E6���������3z���=� %�i3C�%f�x\n���b n?�/s0�����~��#k�C�+͋Py ��M�X5ĳt)�/����.��g,y�h�5�/�TV����9J�~-���J%
o`�ja�H��J��2��%߷�ɒ���>��o�����*ྥ�s7���)���c?��h)�,ʺ),1�f�3i@NS���o��-�/n��*���}dJ�F&ff�P�&���F��4���z]�Xk������g����v�q�l��߿k��;�%�^�q��CvlR���B��O��*&���UZ+����ţ��Q�j�2��2�u���@�3����Vp��Yy�"�`��}�]���)V7�ѻx��\�]����7�Z��*�P�X{x�0��]�I�W�B��W��-��CMY
(�_��茸W�a��� �0��ܵqȒ���m(�v���F���d��<^9	��9��Q�8�v���RҤ�wM����b�����㋶�Q���;�7�}
���=Ʋ��y�j��������4�A���{` ��\�����x4p���hϖ�'u�V�0--�,��»öךLƹ`�"�����y�:]QP~�V�P����p�l�X��l�a�=�*y�C��>um��Ζ�C7.��m)��7
T�N8�cI�9�n�_i@�!s����\�k��m.
��Xx2�@�k�I��U�O+�ٽ��X�cmӕ��5��o}s�og��Fw����R�C��#u��*�[�������C�]���B�#��֓�%��RN�^Z��я���Ε��x��qNw����>��UW�|0�=)�/xc�ơZ���ܵ�b6��\'h3��I�k�!$�����V^��~��
c�������j��Q>��M�И����cn"���a�Rd��✌B��
��Up�jR}��E%��Q%��ݠY���h򾿌霬R��p��}
e�0
����Q�L���%(���^{�_(�$ƈO���r���7 �g��`g� ���;��l��	�z���><�߂-Mm�D�և�NIyyħOr�s_)<��qQ>~��C��s��K��Ӌ���˼���au\w�$��� D�vs���8g����b{�D�!x߁�z��q�u���sr|>c�|���0�2 ��ԕ3V��:�ȿ������D�,�I+�n��Y��q�bہ�9>�;w�|_�7}��J�4����Uw	���(������R)JQ&_ �K�D�&ZN������2��h�P|\���	����g�2�� �����|
��_a1�͋�9�cu~���Ô���tR�=� �ߺ#�2��;҂2R���ߧ�V���f<�r>q� ���"� O��ռ=���lg	c�u^e���x��q����K�(E��XAPh�mw��o^G���.��\ܫw�fܳ�1x��G���������lpmN�"ҡ��U{af�������/��4�*^��q��K� _����5/�w@� ���`E` ���f���z �/3 -��4RB�����'論��7����v�Ɗi0f�uD|�{#����L�R��S����~on��x����2''����3�X�"'�dnb�=Z�u���\Hjh���ၗP!%%%�u�8���<����rU�4Zn�y�2WT�������P�����1'�Bnw��U�/�P��]���wA��|����:K�w��YYo ��6��/��mKY3.x

�\F�w���>��K����v�s+$m6�WR�l�A����ÈF����EP�(g�ZSdʷ��,~��3Ǧ'��F\����B@�?��<� HJ��F�돕]R8����&RL��Ǐ��4���USP�M���� �
=���F(&%����Ħo]þ�g�==��T�%��G{J�O͇>5�/ېZy:�0��[�n�ZZE���6qxH���r>�����"�g�6$��ʒ#+.�Ύ.p�>"��
Q���N��xk�}�f|;��(�d�����f|m�[`�3�?��%�GքMu~{�  
P�'��Ts�7.Ed���{�#�hZ��L�X�Dd>P)�E(`��#�H�gc��|���)��3�_��	��Wt�Zt�q\�I�bt�m����W�57���)l�U*�ck���d�!�zR["(�?���t��Y���7"9���~10��A���6�ε�ol���u��.Ri��+��_ �r����E�6�K⦣��ra�z����:*�wӍ�	Pŏ����:��;g�{����qH�t��\k,�_��q��a����'C�I�ꔷ�����ɖ�����#���s59I�x�r���c&��c�ǒa�'����L��	�vG�5w	f���[�X��?���@��X	�c�'�N���5�c_һ�̿]P�:��Ԅ�(�`o�u���1���A�M���d�˰ 
C�6egu�1		Hbے�vd®��� m�mw�y��1��JA��ً|��U��;���g��je+7���Fʙ�)�9>���(�u
egWW������?<�o4��t`�3Ԫ
Ş	�m�G>������z����B���ҭ<�a:��c�{0l���'V,rG>�黑w��0Nɿ�V����sJ[�Pr˻�6ƌt+�R�Ԅ����Bw7}o�e�z��[`R �m���M��e{�0	#x.r�^���*�O�O�d60���XPrz�"��J��X?��j���¨�������܂��0��@�֯.�`�P��ɚ�Yɖ˺���� z�,���#̑��Y�4��թQ��T�E��Ǐ?|ot�\�^Y)���U�շ~��8v�/��*�?��*EH��_�SJ����p.\�� W����z�5�N���fM�B��TOȅy�����*^{X�0�*>�+\!w4 )u�.���2d�J��IkY��8]��[��a����9������:_"+V�Z��/��O^/~���F&&�?���S�rk�*��L���VMa2 ���l���W���{�Ϻ|:B�c� ��F��EG��܈ݭ��?Fڋ�RC\l������3[2�OL|4u`1<�uj�e�/N��w(�E��Ӧ<�q��`Gw����͔�3�]r�I-���F���-�j�E:�IH��7.�82E]��_��V�"��*��]�9��qǞ�C�}@�tTY��Wj��qQ��U8�7�j	�a*!OW cj��<����|�aƗyi5�B���SU*/vBԏca������� 2lԄs��P������\��"}��H�--�m��J�;g%�d&��z���RV<[8NB�4f�q3VE���fd>"�X�YoLL���]��,���g��ơ��y?O��<�v�8���⨾��=����BO{�z����b9+V�fi�>7���cô6�-�H9)��(��ˮu��	6BOO,������7��`f�?ִ2�\�R8�`�a%�S����z��A��>'�M��.�G@?\F�d����)=�r�Ț�GJZ���M�|��cJ�}����ɐ#ױ��w�\�7���Y�sؤ(A p�ж�x�ח������S�eu�+}��p��LǊ�u�=�%�J\1�"���e�"wp����@<���נMbݳ���+�Ş$"��u����59U��"K�hm.�u|���?�yp����Oѿ�ĝs�#�M��䶅"��5kkS>q>�A��z�=v�Q7TǦэC�!��PC������i����:�60S��Hg���&7
QVd��u�M?����\#*]�������e��G�ܨ�y�qF�V8�W"�J2�����m<ϙ�A������P�xlL���nN��ߝ���KYQB��`0�ϕ�j�Rh�3̝Dh��O�GSc�T�im?�8p������S>���"qu�W��KAW������4X����611Ah]?}C������#���q:�$��>H�'�)�l���'�q��o�]b�n��W)V�S�9� ��-�CFo�z<�׿&X�����ǔNb9FFF��v����`Ry��C++YhS�4�xpejSP��P���C�g�����PgD1��i�_�P6��e���8n'��9����A�8���Pצ/�{k�y�^���o_<�]�.�0Ƹ9�����
�S��cɺ<W��C/}��s�ڤ/�`i���hjiM/^b���~������%�.Q6&� $�XrO�/Kz��Ǚ�ȧ�S�pf�{�-q�P!��j���Ȳ"�Z��u�j9�2�q��Gtx��F��ň�Y��k^Vx0���n$Ϲ���0ie��J�����o����7�Dn��r�D~� ��Z�~�!E�"u3j�P؂�$���,��}rl�ϝ���sQRW��I� 3�x��lh
	qwCJp�V�#1@���a�@5���M6����kfƫ�֍��P�k�LQ( ᥽�!'�V2`�T#�Bp1�o�i̥����gBw6e���(=C�;��B{���Y��!!	�|
� M���M���Ǿ��,�8D0ӈ�&���52��(Ħ��O��]MM�V����A��V ��^svI��T>yv)��W�[�Ī��ƣ�9)����]ϔ���KƏ�� O)�>+{/f�mDh�$�YiSh{���>̹�̐$Tt�]mh�0��]��z�֯C�X%bYx?���o[��XRh'Ij�u+��x�aִhv���V���:P
BY��܂"��ɗָGOw��J��w^fx�G��Ϋ���g��vL���d��jYV�Rr����.p⸩逾��x]+���+N���l�s��r�pffF(o����Dي���X��;K��d� ``����K z�j6���U�F�(Hu=����<�"�����DZ�M�Y��<�ҵh���_)=1g���5Xq�L����b��0'�pF��������=h�u���%�ܤ !j��B�sleEJ�a}[���{�Ն7.CG"�; ���i�O�ho`���-�
E~"�	�[�����Z�|80%SSS�Dh����0�r�C{�H�����Z�x�_��'�Gސ����fU��ǀ}J��A��
.?�<b�1���ڇavӿq8��ЦXyZS�*���<oT]]��|2����/9�l���'?55Z��H�7������:f��F�����1�+1Lo��}92���������/�&n�IuF��p�o[���sb[��wޒ
no3qފ��K.�=�_��L��@ܥ�"����Rwr*� F�M���N���͕�C	Tht��9εtv��`ro=���ؘ��x����67g��3%¿{M�F����Ni���#6i��4��]~�˅ʀ��C�Μ� 5�D���Z����]������Y��u4ڎ�<@�ͤ��X��O��m��&& F�6T�̏�,�_���
'K���l FJ�J��m��[����!nD�������`��4(1h�	����S�pm���U�^�"& 1kkg1i�eKK���ץ���%����G�o�_��KDz�t+�T��*T%���Fd��3f$�N���=�G@@�n���=?���4 �&%9�\b��ƚג�����2õ����E�Z�0U�yV���#�
"N)7/��0i��2iiup����g�###�{�ȐǦC���bD@����(m`��bt��Ban�!
ms��bA_�豢(W�T���Utz�x���� ?W���x�~=�W��Y�F�����DT㼏�:��^��8>c<ܿ�a&L 귅r�LH�m(D9�n��F;6?V+�"J�,�ԏ�Ӹ
�fMS���hPRʧ��v"��Ԯ�5���X(��;
���\g/"���!@=l�Tm��,8@�4�~qd�����o�E �)�ou$�4��>-�{r��=���7���K�D$�5L`Rq a��Л��+�[��.X�5+''�kkv�6*�w�	� �x�_�<��}���gƒ ��c���'P�.���������}�ǉ�l'd�	yKƱ7���!;��{dfd��!;�^!N�N:���N�w��/}�����8�D�����㺯��19u����t�OO١���C_�,��ÿ��_�Q7������]�E�&m�F�[��Ũ r�/�ˋ�Z|,9�>gĿ�-�e�4�W�,x>ӟ7��lh|dV��A�m�la�d��7�'�D˃'�Z�dR���><�
$ �8jNDR���gk!�{ 
s��� ��
� �ݖ��6*�&?*��;3�n��.���"���V���B��7�t���T;ǡ�<ΠG���>��^�U��k-Df���w}/HD�'G��u�+���[_::.�t*��XYY�����[������G��,>#G��I|ެ�`vv�)Y�D����,jƴ� <���S���[�B��A*�Ss���;Q�{|q�%������G�\Q=������_�>�Hߩs���V�,��'x��f�3�u��Y��N-��،�y�VV�"�痟��Ӵy(;SUj&ydV��o�z���z��2&���2S� B�W+}��Sj�Nɫ����[}������i :��V�b�9#|�hK�ɢ8�ͭo�g�ҫ҂種�6�?�F�ڱ�]����"�W��l聙�L8�TU p��J])�64�����}5�>ԉR2�WK����߿/�8����L��yt��1�#(II��b97�\; �|���R��ɣ��{8�~�-��c��c	��3j��?�n���zn��4�'�=��<1���Jw:�>���~/��u���F:�%.p�M��X���6y�\7�Y�"��ņɨ�O����Uj���@�%i�]��Ij����LU��z�U������l��i�:�r��Kp�J�L�L���#e��/e������̥����E؏m) ���m2����'�8Z*u�Ļ���s��;i�P;�X���q��^_T��X��:L$iկ]Rvf���1$z�O�v��\~-�:9
���7��(ɱ��T0����w�8T�6��uͣ��˽Ġ&�ET9�����p��wehhg�u�[�wS��?�i�W��&�1�4K^��T��.s����HA�� ����v^:��u���v_Q#q^�`�R5���ܺeZg�]����A�NB��[���-��]��F�Q\�t�?-�lUW����M.��g2���_r�q�-e�ܭ`j/�k@�}�[EE��B?���N'~ GߺN����aݩ��]���ގ��n�rt]��SR�n���Y�?n���Ya�-a<pl�j�<���~� -�=�z�)p�,�<����ܹ�x/_�
�ͰT��~�2ުNZ9,��:]������M��;�t��A�\��Rǋc��3E��f�J)�P�A�?4��+�^j=�rA0k����"��Hw����r��
 �����סR�b��}�ʵ�U�Zet!��6D#b����4�XaY7�� h�[~R5 Ғ�+��gۤC;�_7J�����.�"��Fn��|�j�e��k\?�w� ���݊QW�|f ?[<�#�r��fQ���sM{i�$*К��+��q��)[A(�l�h�e�mp��Ղ�����
��_T	$�N��kԶצ������~�$����w�/����@�R�<�F���o$7ɡ^���#�ݹ��gN��g�+��x��]�h	H�Mh�޽�Bp�ɠm"Z�xԿ�BC ,���)�ٜ��a�*Nq��-��ޭ��>�>�@�D͢��$®���i�8� �2�klk�o���¤�+�.A��g�!��N�{�<M���(4Ӂ�?8Q����5�:0�*�S]�
�ϥۅ�vq{�����9�?-d��S}��r]8��I5 w6>�3q�k���sS��\��V��5�4utD���
9J�Z{x�-��n��k'"L��w�<�&\�U�bc R�M��;>��V�u޶O��t$���81�������*J4�4S��I���z���T��բc"��xi�k�W*���ꛘ�I�G�hX��'�2�=%����Q+uZEϭK�Y� �(~�jZv'����$�~�4Z	H"�jc�g��Tq/����1Q��O����Fv�P��o�X�x$7�,S2���Nς'g��w3�gO��?��wiR�����̧�m�=�e}���ݭ.>�K�}J]P�1e���j��n+R���f@}s�Ñ����b�h�������B^�d�<[鄋Y�x�=++%h���"z#�i����S�kO}�S�+��-2av��ٌ����U��LC���ƀ�|�_~��r#^ͮ~z�Ni/�0G!�>(J'���1��8W&
G5���)��ʱSCb��u��U^[K7�).�Jj��- _{��j���rpx!&e0��^��t�˝����C�����W���^ٖ�Y�2��C��YB�)H���h�n�i�8�����)��� ��{���:I�mq),Q.5X��ؘė893�,-wx�tB�� ��K��-e4dLu"?~XX��s��k~����trA#f��+���@�gty��}��F�ۻ)��Pé)���kJ�{5�zz�WV�	��ou���; ���H0����s��k2;�o�o\�9�QR�v�/1ʱ���d�U�	D	���<�ڵt����S:6
�R'���3���C8����[�uG� K���A,�60����(S+����,(��W�їՂ��N�7L��&�<@�5����g����ʃ�)�d��W���v������~��B~���jI���T@:m�G	<h���9*A�O?�oKY\�� ��b�Φ��� =������)�Ù6I�����wD�@���/H�J�^��as�Ȼ�au*A�6�Hŏ;r�w��e���-�+��:Fg������ϴ�����:�����n���Sf/pwK���du7��8�~E�,�%��Q�WW��Y�l���r�W��6ͽ�,�J%�DA�Q=�L�؉ّ�=�3�7Fr�'��a)�p�tZ�EQ$��굎 �����>햀�*��u���"0K�|05�<en�fG�*E�5q���D��^�;��/_��P�>+���m��u�aa���*`�}�ݿ��ktZ�Ŀ9��Gn�������<�7�(�>6��N�	����㱫o���î���^�*̍Ԁ'��9�窕��Kݜ!G��_�;�7��-"B����<:!+Z�F������z��s}��u�G�b��B���2Q	�h|��� ��.aP+�+�C>��V�k�+>_5�t��G!�f_������=$v��j_���-Kr,�R�XS��=,�jo�� �A��+Nt����m�%�K����Z���#�e�����W��}}��u�<{������"Ɩ�����v4� �9	�CCT���:!�߼����x��|6��"z��M����r����\���o;�`Z[���U���u-w�5u�СZ������Q�zu\L����ddG���u�@��|���R���
�j�D�5��g�91{k�/�al�b��U��=�\���[�ɿ`�=dV��cX�K:lO���Z�ë�\ę��yJF-F���c�J��KgQ�r�޽���|���"@���ڦ�U.��������>˗�|󩿜�\��Ȫ�$�(NN֔TK�I�������gF��94�S�,���*tp��aH� Óa��f%S����D���� � �z����T�>R�yc�H%P��2�x��ԥ<�GKKW�L�o΅UO����=|8zmٯ}���~���>����"5�>iT$?�=;�Ɨhk`�s3M#��荋�\_�߄g���w!���8�yQW�1@x
f�K%кs�H�M�,�L��0B�@���ƾz4���]V"[-������ZN��?��W��ϱ7��/v��Y�5]uB0�G�%uk��}����J#~�g�zb�P-�h�gVuf�Wu�˝����W��]-K�z���קD��Qi�U�*^��2MQwq�{�Y8��7	 Ua��)�Y���q�:ec��4y�xC����2�.�Wsg�o��p�w��<}ޢ����}_��~�]M/���ߗ�9 �;}����V���0B�Xڶ���Ȫ��%�Fuq�.#�ި:$�h�ͭ%��rm�v@���2h�BO.�Ǹ[cZ�J���c�+J��,���R4��z�x���Z�U���ܘ��Zgs�s��y���@,�����^�`�kT�7��*X#]�BK��5?��!��y�^�<��;��66�=�"9c����6�S�/�,xڣWˁ_Q@Y[XA��E�H�q�6��O�/�K���%&�k'
�� T�<}���}ꎺ��ܳԄ쩤�ī>��ծ���Sbb$/D�S\,W��s +-��C���tx�{q���0����B]]}Fp�ݥ�\�����A�����6%ԏ���5?�fs���ޣ��r��N�S�����slJN��+)+�c���S��7E�1ˡ�ë����pͳ�r糞�W����Z92{)��*��|�3k�4����NnI��*-Ӈ6A|�2�x���C�w�9t4 x��^�ZK�L�ۊ�n���BOu��x���cƝ>���K�j�&[$��9�g�$6@6r��_��R,R�/�)ȟu����I�-���r�!b�\����v9$4��u8��YK��x:�w����?�rc�������跡㝳r��=�d��LӞO.=�Tz������f�C�E7�����bDa�,��I2!E�yy�Zֳ�$���]����ZZ6�*D�Ti�)DpZn�M�Ն4���>[��g�35%%z�bE���_�D��X �/�.?����Oul�wG����V�b˴�Qg-^R2 a{���0�7x>����P�%8�]�.�}�TI�H�F��HFfze7H��JG����QL���7*��)x�6w���S)��h�Cn��4��u��/:w��ۖ~����,qz?|6�	"�/���:�?�"�9X�uָjo�j mjn����H=<T/�{�"89|��X���\�`N?&'�66o�^�����{rv���MC�etq�:4���8j*j������kJfU�t��d�+vv$����Q0�>7���)j�T���z��r8�'�=NX~@�ⳋ��C&�:ʥD�:՘Ca��e�ߞ����c
}33�@+{���S��찺��tߔ�u��O1]��I��0{/��Ƽ���ΰ���e�_c����'R�8�P��j���洬�&	�Q�`"H�ݯl`��~�A�t�����|,�N�9��r����
������_c.Rlu�/��JӪQQ�}K���{�'���$�����
_P�h��a�ro��}�>���N�CF|�B�� C��{���_�����{�DgM�J��jo�Y�i)|�R�������gi�"� �S�� ����~�פS.R.�8�nϗ�;}�pR�ډ]� �6��2��ӷ�}�"ovy[��e˃�lT0�I�UvAǎ6{3nx���meQ@���z|u�
$��C\���59#�\��V���v4��o���t~�XX*O�fu?x&֦�T �u����q��{U����5�	GZ1
v��Z������{?�[O�Z�O�Ԋ��WY�xO?�?K|��+�����쩼%��Ҥ:���L��Pvvvܛ�_�$����|�stp�����X;�4���&��SbB�bAsݕc�:H��%J��O�V /��S£�|Άhh��ܩ��Q�`��}A�&1�;�S�� ��n�{q�)֫����W���Gn��Ԯ�,�*
���<:!���&5���Ȣ"w�kL*�n?��l�'kN��b���	P+r��}���+G���T8iX|u���C����0^�W�mQ�ńK����Wj�K��_�S0(8{��;A������z�e?S�!���	�H�mmꗗH���xa��k�
$����a�O�S�n�G�ЖC�42�����
����vw;�Fo� SI{��Y*hȈ���4L$��s��6�����^?�ɯG�CC�nn�d���8F��� df�»��6��TӢ	h��3����WW|�V�M�2�h�
�0G�g�}v��7@�H�f8�ƒXu����5&�����~��0��pM������:�P�o8j�$_R�Z�ď�ٽ[߷C�>4����uCq�Ȣ�f��4?������P�ӷ&��4��� FKWs��~M� ��Q�$��ǔ�=�����w�3�Rq����(V}��������e�ݖ�DW7�����+���%��^�Q^p�u����� -b���`(҈�K0� S�q�b.��V<4^�m�5s����ݒ/B���R�܀7�}W|����f|��r'�8%��[�Q�xj��_���䚟����U7u+�����1V0���%zJ[z���Ŭ�������%���72V�R�1/�恊��h��*�X���{����7���ei-!�4x@`�0&��qSpg<�X�m���l_^^��:��)�m��Z�f�2� ��!�פJuA-��įr14���q� )A��'"�駏�X#j�f�[Yyx�\���������<�^{~�ͣ��^W�Y�Dy�O??;�6����H���WV���]��i.HO�������C�nğ�[ѿ��ܪn��#,ybb���x��� D��ښ�A�=]{F�D��A澎	��}2��~�S�4�d:<!��G߄×έwoO���QwZqTU)c?�L��J�kF�/����Vl���u��[�isb^�W[ٙ��tQ���xd����wԻ�c�~�-�SQ�W�4�^�yP�~|i�,�d����Ç��$�z�a��}?W�s��@�����������COKC�.8�(�����r;I2��G5����+i�_���СB��M�3��1�jC�-��T|�����<c��ub���hۆ��Yw���U8;\W���}BPv����>����O/cX�gi]�e%�r�
��TІ���_19��şs��EE����9:�����ܭӕ�Jc�0�ㄑsӐ�'Y����
"`^?���Z3�P��q�uڬ||���d���}�������B��~|�d�R�Y����K����)4ӹ0[�u��cʝ��rB�~�ܿM�&����ӈ>}{]��jGH�X��~<g���$N����p̱L�"^h\(r��.�>>�V��}����޿��i��  �Q"�������~!h'�E颔���? L'&|18�����K.ͽ*�H���m�3Ĕ��p+<?����Z|����͢J��8�4(^&��XI�'���n	�ɉ֫��e�v�HI��yJ]�j�9ƞ�^ljZLӀU��ivy�W��|���nbbr�5'��֯�L��a"��Vj����
|k �ۏaC�J�ll�����J��K��;�d*���Sr�
�|df]:�d:�t[Ƅ(^M��S�Q~Ƌ�%��x�3�K�_�d��Ƿ�?9eeK%���k�[ZOR$���ʮ`�z����ܣ�q�}��F mўA�*rZC��0$ �}S�t��=.��ĠN��5�O
X��W��ńI�=���7��i�ԃ���d<���3い ���w(ܸw�{�k������'Ζ��J%O�_?��e���P���N��'�Ǧ ���;���s��)�5Ga���*%��_��&�n�o]����@����Ss%~O�Þ`����0�5�`����}������*y�Z@Aǝ�z$\��h�hƞ�����H�\cˆ�ʵY�����=�f.�10�2==�h������h#�;������s�� W2ȉ ��gŌ�U��FʱӄP��3�����?N��{b8����h����"��:\���'���K���ޣ�ɡf� ��DS�
�T�L�8�˾������ʉ*��Z�ZUZzzay�8όh��aUX8{�C@h�\�/�KX��d�y��֡,�//��V
U`����k�ȽR�Oy,^W|\MD]gU4?Z ��ш���0?�B������!
�|�O�?�3����s����j[, ��,w�uTK��~T:�.,D:D��>��{3��x[WWW���]�Hp����+yw;M�MX���M�6�!v��������5�Gɴ�Z$0�Yv�j[��/V$2�G������ou+�Lk���
c:�`���wØŦ0���}�߹��R'�s9��y�dnJ,��a��fya�@����O�l`�H��w�:4���o���jL��d;�}tp�>�lf�L���MW;B�!&�=�٧��$&|�@�{�*ll<�Я�4���7Wwq��.p1u�����4vh�h��#x����R0�����?��i�:;_r�>���;>~atp��*Ū�B���/+�,����,��\�Ƅ>.�T�:7���y��E�g��J:������^*j�����V�d�ĳ"��8�4��ğb�w7�������1|�ňpwI*qx0��H4��mӅHfJݴ�h&�[�_��bۆR���7T:!ae�MM��GG��~���SY?��B"��]NE�	Q� kz�g{yn�x�)��uV�:�YYE
�����'_�$�'����o������J�0KQC��S��'�ŭ�'~WcS���K��q��r�Bu���x�:?02��7l[G��'P�`�=��&��ER`0�ջ�H#22���MS�;8;O��z6/�&cK�%r�˙׿����i���̅,���!R�4��� }K;���`�h����
�\� *mr�� �?�������J��!��r1 o�ӷܴ���_G�
8�o�u-|���KsB�D�	�ҹu��_��ς9Ec�d������b��jL�;O.��N?I���y����?=����n �]��r��$�g��g��z��Bv5jz�m��G�$��]�4��+�͋�z	�i�?r���7*������N/� ��T�ٹ��������z=����ٻW�|Y���#�	��O�5�x�c��3H�!�;B�v]�Qa����~�r�tx�K���}�:߸�E�np��3���iR�q�� J0Z�+o{�|.��35�O�SO�������22qn�Q-v@�:2I��i�����s��s����~�����Ch�=%�Wl��Ӿ������}���2=�?�u(�>1��k0�%L�O����;  ��z��F�P���j�����C�8�XHq{�>���3��qtU��Y8��+��+�A'��	��켼.m|WK�,yKJK��>Y�B�ዟ{�\� ��$�Ǎ-������7N	L��[�6K�`�;�Q��f2�6`	ع���v����A����t��a�/Hٱ��D=$ҧ�:�5���wP�8���̫�;�����|llF-Q���ǝ��C_��������6�.$OF����OQ,�u\����'�j�ܱKKW�mm�r��smv��2?H�w�t]�ʛ/�F�6�DC����?�z�iIu���"��Y(����/Q[��5��n���?ݔ/�H,qsbMg���u��Qৼ��-�(�ߥ���%7Imxq�{u]W��"T�������6�4uݧR!��Ζ�-saD:���/_��N����y�Ŀ��=4�S��|{��[X�Rb�/���C�����A�|'S��#���Pg�W�-mZ�U��AKO$�5s2�V7�-d�Ȁ��2��j�����32<�I������E^���!��HN<�;ې���)ڤ�d�e*3)ָz����1�dQ���00���:��Pewh�B�Y@�r1QP�2�e746&:!KKUt�3�+a(Nt�ǘ�V��a�,
D4�(���r01��5@�]Q���G�`zh�������%vY|0�{�-��r�EE��p�%���0��B?{Aף;O����W3ݪ�j�'tr?��z�5���F<�"t�ϫq"X7�4�
��o���K�.�z{I$�@��k���i�qT�k�d�������.�,�̼2��#]�?��3Y�ך,��I�}�[�3�����ۆ��βm�R2���MH;lu��Ӗ
y,_���8��U@��̀��@�Zu�������H��/�n}n�3Z�{��-G��Ӳ�xJ���Nx�Ë�����R��Pq4�~.'YnQ���넣�Qʽ}-ҟ�i�v�W�{H�#�����S�9e�h�VE�7����!]4��WjUW�]���mc���Ã.w]g�"��|дF�ږ���$"�,M8��S5�/|����s�������,����������_��B��@N���]����RJ�U�m(^�.`���~��߷�/_88 ����=�G�6�:
}�Ԧ_��-��e��I��&$'���5�_��BZ/��H�ۦKG� ��Wp����������� =$ٷ�N'��%���.0]�I�_�NOp�0�S��`X~�2�K/Thhͤ�B)��:����S��3�}1��t��vK���(�R�e�#��_[@m�~Ӯh��\����nE��+��/��Tܻ�?g+F��������N�t:����g��\(��/_h)b\�O�:>�ڡ����V`_�C�3��k?��o��ND���q�;<�ֱ�F��ڞ+�irF��z��ˬ��E�cL~)�y��	\���d@Viy`��p��=<E�b���j�}-<��e�o�/X� ���Z�E�fK�y7�p�j2��@H��
��>�rQ��>R�#��� �J�����`]�d]�U����m�*�+22n0��:�Ak�E��,�t~c����;kp0`�)�ŗ�" �hk�Jd8��2�zZ:e䦡V���Ȱ���0��+߲�<��S��w��P	��� Hem���/?������cY�Ŋ��o
Z����$t�,�,��YF\�m�I�A#�	�F�N��@?��*~�9ְ�Q�ӊ����K�:oi��]e�9��إ�zYFzK?~ժ��P��T����OO��+]ⷋ��F׵! n�rI�����M��M� �B�xjE��?������yp�uj7�blo�~��A�K2��	�̶�fW���cCS����L5�:����D��P�(E��c�:�y Ю�+ a�%>�M7�����>p��oi�ll쮭�#��$�		>���>��uK�Q�k�[�����/Q��7;e��l�V��D(WU�-
3��n��p�ĕ8�/ٿ��{���/6u�yU(�a�G��կ{X���?+��2�=�yT�;%�s�g�������Q�l�h���y��4�2&��u G���O{y����]y|�ͣ[�z`lx�8bi��SvV��ux8uY��#}曚������ͳ(;����ƿc����}yy�d�l�dS*+���n�����@�9��}�:Q�bu4���:���YC����`�(&�cWC��~u�A�����9��_<v��g�*קIV[�n%�򮑢_H�f��ߍ�u�R'2`z�k�M�}�LBU�
p�R���|� i^�(}��|�`θ�8m2�+2@nTF��2V�9%>��f�[u�a���Jm��?~0�'��@�鍩�E�{�_����{�H���-�x�d�ɩ�^��k�r�� �����q2�n�Q���NP�3Q���=���\������u-��
�n�g���O@PS�q\TA"lA����|(]��ӭh2k��Yt�	#G�󁙝�M�7�1y��Փ�w�Ybs��H@X]�8�7��Լ�[,��{6��U<ֻ�ݿ�Iq"�:}�$b��0H�k�;���G������};6�F��n^/���Y���ZY�r�S�wii�&/���ŅYT�)�0�rɓ.ZJ���F� 
(��.�߆�g+����f?�j����jɓ����6�͗�A�[t�
�u4ԿM6��Q�?:z�Ё�"p�0�:�Ѝ?��� O�"2�("Wb�~qd��˖���+D�ȧ;\�/N�8̭��1<�͍�]�-�x7c�z�<���%�L��
�:��$k$_���.Lx�$��| -��u�s�
KH��V������m��WdW����y��\Q��M&a���8J�M�l�E�;P���j['��;���O� R|}Gw�j���1���<ׂ�X�H�+�ǬhU`B�hT7��c7��χ���PH����:.����W���Ī�����869ۉTM��j�[Ȳu��<�V9��5��`�S�.[�n�-�������(@�F:���&=��¶K��tqpɢ3
��)��c����Vu�'�889e���r�>��
��� ���2"A`aQ�8Q�eD� f�k�c`|������e}�r����%�I�0:��A��&0�|�2J���zrk�^<{c���@�P�����
��I�i���[�Ӝ0E�]�x��7�*ol���H���:E4e��0�IG���+A9 ���o���b�����`ۀ;piN��P:/׀�
m���O�?�p.��R#���B��ľ��*�xW)�T E�4Ҫ.�	�]�Ks3%�B�x�M�װ�S��!5a�P�J���Q�p'T2 忬����;M>�'I�_����FSS���j��Ys�/v9 *��S<�?��	K�k�����;�Z��|�q���J:H\�#:��U��d@b� F��ʮ��T�U܂5*?~	͇�sB��;�P�tNq�]�N��n����Pͳ_���D"��`Fj�d� �ƅ�^NA��T <ew<[-^�T���ڹTB^��P�.b
? ?��q_���˃(1�j��S��r�:P�AA����`99��pn�T�[����_>��i7�_��7�ɮ�����[�����x?�`q���'����g͵�p��A|����T� Y�,]^���_����v��?n#�9hP�7y~�����i�Akc���|>
>�1��N��Z�Գ?�0�~:�\�?~���:�rr'�l���!`�s��voTq4��.~�;�npv�e���~���W`ң�C7�\&�2��l�k�_m����|;�R�� ��e���9E�S�P@����xx���Pß?#,�_��\�rܑ. ��A���^.�e8ޟ�yu�v�	���g�Q�lEm�4��o��BL�JN"����(��T7qW;��L��*.֔�/���+m)�(���ON�3����y�-�,�l�~D��* �UW��ҭx�2��ޛ�=�q7(~mT���ƏaC�Նjh����#����=�s���י.`��y�#Α�$�������}�!�v)B<��>Z 166��C&�3�Ō�ny��s���T�`xQ!�%��sO��Gǵ՞ѳ�A��[�]�@���9ܟ�����D�+q�a*�A�yM���%�l�/o,P;�rfJ���
�����B�Թ�u��a�� #X�]���6�-�g��QGy�|���c��J�Ұ�!��Yں�7gm��S�C{{~㨇#*QQ�������c������NDO�'����g�׬��C',�?�n@������^[��$�[��]�����"wi�rN����"j=��~�����nF��^�#w��e�S�Z�9]����}��Ҧܺx)�_6B���=Ju� ࢋ��q�]�B�r)w*�Y\�������5q��-.m���-w�cS�%����Z�x,į��^���LG����(
�s� �!�!d��j�h��&"#WYyӆ���B�v5��36w+�Ɇ��l�˔��K�|Q��6J@�(���/G#�;ǝ��)�e@2:�A����	rb0h�u|��=�WD�Fi����	��}hΤz����:�/q#��bJ�:df��U�t��	��Ŗi�٧LA]~!�2�W�f��}#��w*a���.��>E���L��(`f���.�	@�����V�Ւ��a����s@n����#�`��)-t��v�+yfff�9,5�F#�u�������߹߿.��vgee%�'�DC���´,�I2�8<ԓ�����vφ�5 .�G�Ã�r�s9Kܿv(�B�k��_�
�\>�6hAL���Vi�uǱfhQ�}V�i���P����Z|<��C�� u�H�F���MK��zz�b����]�ȒH�G����`��
],`w�p�r�H�x�ٷH
�{@���ׇ�4��}�|�<��d���\�P*_\��[渀]�w�ýϵ��{(,34u{����r�Ç�(u�ȥ�+X.hOf�cF�n
s��8#c�{������g�SR<��&���X<�`��nf���QۆK�Eѷ�uZA�҅A*�,Aio_	�RA*B�/����1�F���#e�s�%�+��m�
V	�Ԕ�uM����Y"A��x��0�31��5&�K�Ԫ�T��]_T�7�%(`_���5������$��JRZ:���M�S���������ͯLOߚ$U'�� 
�9	(����l���d�;	��~���vV�uJ���`B<;{&fu5����:s��\�O����C���l���E�/?^�+�Ʃ$v�VCok���Hrt�V�6�w \�q,t�Pv'-Y�_�}6�?��"��Kwɨ��8��g�	���аn����V}@�~�S�H� qy��p�kg��˃��`[�J��wyu�M��7�|�\^�r�u��P0��R��H��+�ϝ̥
wc#�k!{s���d��!���_�ږ>� ꥒ�jS�񃆴z�S��4�*���}�h�d�j�3g�J�$�����5?���z��K���.S�I�74A��j���_:��t�*U��g����n�����s0�G�l�����I��LD;��Y�x�M�����_���'�&�/Dr�.L�BL���i���ݒ�Ḧ8���IEI�Y�����[�7+$?��]���
'������m]s�|h�Ii�
@�, xcbx�ŀ}𠠸X�3M�����r������ /S�s��Z:�i(��ԡ�%�z��vz�h�@�n��s��	�rR�8A��@��ܢ�K��tt��#$�d�k*��˯��zBo�� K��'��������ᓱ�͏�>�Ք�?�pzfU�p�j��gF+�{N��5�s���+M�>�"�!|*��-�}���t���Q~�! �}��Ŷ��s��-�������x�����17�K\���ǌ���{c�9���1Tض����
 ����\�ڶ�v ���G��T�a�yaϪ��uɉ֤9ޅ�E7�.h�ŋ��Y�k�^��d�iEmUG-_�a�ܿ 8xi�6	��' r�xH7R@''eB�b� ��!��n�],��_�v	W�ԡE7�����=-�y�'�?DOׯ�x"�B2��V�,T�X�,��ӻƼL/�a�SҐK�y��ʷ�Mj �����	��d�rs�krz�)}��ٙ�Wg5��=^�W�U��
:��)����<M;�l���7���������Ҳ;��A�P��_Kl�?HU���s���`
"*��h�ZD�;�����B���o�y6LN�W0�>��4YZ1�EC�V������μ�T�.�[?���� ���ڠR5 �㮥���E�����^���>�r؍ ��>��ù��*�����v��q��:����RRj�s�1�|p��x����n���saooR;8@��.%`w�W�'�Z�,wҲ9��c���e:D.��m|}g}���Qg#�+!�n"?�q������U#ߍ��0���Sq5����?թ���v�yo�iUU��F�����Ֆ�,�rn��f{3�z\��,�<
�o�b畩'ں��� UlӒ���@~��Q�eo	A]TBr�A'*6UNf>���"m��HT��9xz���ei��~6�sH�Q��..䮮,`�Qm��]G�ބ��g)�e��U��x$Ze��<��"��ٖտ��:^sњ�Jg�_��8��:z�����>��{�z�����Z�-�c�4���+��y����	���,�LH�����ɿ��e���/?�I[��@�HgIҐq�*b%ž� ����nD�T`/���h��"W5�r�% %�NI�8�/��|l������H�x *�2[Iֆ���{3�~^�>����ȸ�#�SG�s�ŷ ,����ڒ�V�_����Z�X�p�7`'gB��TC�����l�������Vuvqc빀�[d3?�w뛚F�� Q6@������@�oj�st�$U�ht�����a�����7�@ܼ�_�8盤�Wיbm:���]i�R���R'��&"�0�gb���E�\BC~Q����H��@����g�����4�����;�����h^z�`tٝ.��+UU��c%Vu���=�>�V6�$� yn�t¶dw����/f��=%Q �����۹�o�zl՘���K(��{!�
���d����c���B���ݵ�;�nA=m,��T{%|3���/��P�j�~�Lv��݌G�}��r�1�x��P\�.��B�0T�L�'XF<�����N��p�j�p�=jѴN���'A�s��iu���n�^�I��r�[�����8�b��Z(0H��ބ��.x>��9j��Gk���E1�Z��بH��#�u��m�����A����.�bUd#1K]��b:���N�ͩ4�T?��=������FH�+ ��ۛ��{�|�Db��g�H!%<oG߭p����ݐ�������v9)M۬����}�^��eil��wVV��9���v�!hr*��,��'�3�8�0Q~��-�x��o����{�yM,�pm��K�J��N�7i-,Ĕ��=s瞧"���˖i���U ���f�S�,l�1��r�P�OF#�[(�GG��U����jsѐ��_<̿NK;շ�mc�p��1ć�bx��`��UFǂ_�'��[����0�����
�-=��_���tSZ	ݓ�ut��|yQ�����1Zn�ST?x,t�/�V?$_�``�8��Y���&�����Qq����
fhq���J��c��O��:~V��G���hR�tX��ة<ՑXċ*� 2B��!莅���! �/L��-,D�����*6��x�~!ۆ��&V�8���m0�F�D�'T�8�J#}>��f�@gX"�*-w���hhC��v��?<T7��Rb����w���J�֭� �bX���A�����b@��b*Wāg� �`)���PV�L������bz8c��۶A�����k�(OJ*5�8㩣7��/=X4�����V\����M��A��U��a� ���S�Ҫ�1��ٜ���_���s>J`x��� �Ȉ��Óv�C7�t����!X���.>/F�����%<����	��������I �� ʰp땄2��"'��ϟa�̔�m���9��B22qYYƏ���\���ڡ�K�eV�jA�<<����#���2;?~0y�=���o������ˍ�(`��a�,��$����D3��������=7���0�FH��R�g��,R�X��2��F�N\[�6�ilϥ���6p�Q(� ���\bR��g�G���8����N�J�_��{�>sf>�x��>�IT[9tt�>Y��Lm��S~�2W�>E˴�x<�$�Ѐ�H�_>�@���a�Cm��M���|6bnP1��_�F�qc��i�4������3���{�P�}	ٷ�$�dߍ5��dI�}��}��3B!��&��i��������������?Ǚ�o	s?��~^�{�{��F9�a�H���u2�n�zuȝ�����U��!r����{���O��/E�mks�7R18��+9fO��wփ�3G�}8�'v�Ν���V��r�ߤ��0-�2��*l�C��DO�������v������y��,��Q !{@�~.��g�yb:#l��~N�����м<��*sL���Je@g�7(#B�d�z�2���m)A����R��$.�P"45?�<i_IA�R� �
��~$"�\艡Ӟ�g���g�8�6b�F+��svv>n`�R(�����x~��fF~`�����6���J��M��55*d=��/�F�D^�����s���J�X���߶>�x������.�P��6.��2���Vю�Aq�#�F��t�����$~�e���,z^a���� �;4���`�̀��E��y3Q���+> ���4��NN&r�������P��.CZvq�ؠ���m��t�f�	W��FQtϸo��.ҭ6��ܙ�(l�.��0Ct	����4_G~�OYOD�)��AL�?(�&���C;}������㬷��ʚ}��{Rg���*��|����%XN莬��s����!~� ��Z��';l��7�5�9���5l��Jx��C�5F�):��J����?�\�����nDP�Y�3o7P$�e&63�HquG��
=���*U�(�.cx����k΢�a��_�$+G/��zR�d鬙�[�5``�M�\�ɕJ�W�����2Sd]�6�r���8b	�ե�8	8I�zJ&�zQX��Ǫ��t.@�Ӯ�\�y�W)V�4��������_V%�kl�R+z�w_Z[;�YM�[)j	N����O�l��q��������u��(t8\��ICE�址�?G��x	� ��l�C���Tc@̭e��}К�Tf$���q2'	ȣ�Ww���,"��2o�^��U3@AxiՇI���bH,�p�ͦ_�Y���N�S��G�����k/*[�P�va�a٨?~Yt�r���QHP��+^�	'�a񣄸e.q� ?����8Ջ|�*1��P����S�κ=�:w� ���h׮1�9?���CF1������0��+Ɛn�*+���M�(0���<���/��X�Kр�U���<��f֥?m��-��)&��� �hI�*or0��2C^4����M���q҅*W�|�!��ƫc��J�'*z)"L��$�dAZ��r�z�x�W�h�kKB{�-����,B8���ip���G� �dέ�v�@�cn^�q����ߍM��T�Ѥ��|��F�H[*�L��ϗ�Ӗ��wrm̅��nI1j��>��{�Ui����iu�<e	<
(����qޛ`�t�3�0"`V�֨�[*ՆH���ۼ����v���?oA���X��K���hdT��s:R�Y�m5��^���Q;�HP�&�e����&����(O�,:���I�����|l����Aލ^	�pF��+�-��|�7S\�hre��'����&>��=�b�a�o|���fl�)��#8�̭ˇ{��KK�7���x,��������c 9������#w�)����\/��0�M��o왛����;����L���S}ڝ bQk�8
�*�V��Sy���&�ه:�%���cs��N�"8�����@�WZ�aϔ=��q������rne��r_���mf��,���JW��٨d�
�����+���r��_�=�]W���p�_��H���E�m�O���͸w����i��͍���5;�Qndj�(�ļ�g���9?�u���d�y��W�B�������[&������H�P)KS�u|,(�E��n��ŝ��Tq#�(���T�Y�g��˖�J�~�Pv�+v���&�28Iڀ�����������1>Q2���I��lF�vg�e�g��/��C���& (]?A�bۯY��(����9<ޠ�V�B�}
�PA�H^c��M?�/�.�}z}ʨa����U�?G!�O��r|[�������J�����x��B0L�>ց��O7��~}Ɗ�=M������*����k�V��I¬eB��L
O�d�g��j����f�&fW�L�0��V��|Iq���]�C2�3<��щ�F���I�?z�_f��=U�����F��Gls?�{ʍ��|�:1�[_��|:��?�&K&���f��$�sa����ki���AU��l�}@̬ll��	!k>�..=���"o{z��x���eX}9�n4����ا��NK���b<^<?�y�!\�Il�|��5Qze�[Nɰ������F�V~��GG+���xI��ˋw��:�_i�7\U��M�d���2����3R��6��:����n��b�Q\���2����<3ޘ=�R=��,n�UO��9�~����% ���

]�G�G4�7$���1+|�ӝO����ϡ�n��?X^]MG�r�s�Tg��^eX��鍻���Dn2�_Xș���� EEDF0O9��vv.;4�>IF�B��wxb�L�� ��  �'����F)hg��,�.mX�z!��I�4N���_*ֻV���L�ĸ4��%�Y�����~�O��{-%>�d7qB �n�n����̔G����yw�rM��Q�H��*��ȝ�*�'Ԓ��{�N������';���߼����ki-|K7SX�9,-���5�qz�f���j��L����ןk|����,��#^��6UcA�U�{p��������8_�bI��x�q����Ĭ'{!E�:BO���h������X�;ifh�T�^P���r-@�`R�0@�����P� 
E��A�:*`W�f݈�����������q14L�~��K�v�mr�����@5k�A���k�L���U�?{��O�\��ӧO�i�:�7�^W�E``*��о��q0��7���5��G^�R4��]~���<M��=�v*���|�.�n$�p[����ёn©5�8�֭[��ƝD����<��<��YYY�r���c�P�uq9Ǟ�_�d R1N�H������CA]�цx����8��gN��/�S0!�OL��N�
֑��#O�����֠Ő�S����ư�z���Iɨk���k><y��/�$u+2g=Z��M\���߶�c���w��)�w%S�u*r�iK�/��]S�u��4���pټ�Qh<[k�l}�����8®;i��2M��~�4rdD��,	\�hN�ʰ
:����C pN`�hI��vt�C�	^W&��hGt]L�Ҽ�~��gda��0��x0����ٸ'Z�S}���^f����z����D�Ѥ���K)>�.(����㮆����
���T����م��c�i@��	d��[�7��~5l������)��-
�01k��'<�Ȉ�i�W�K�Ҋ���O
-Ԕ������XԒ'�n���O G���Rl�g $4,�O�@�_����_�*�#` Ύ�4�#W5���[[%�R���U��
*T�fv�%�_��/w����{��� >Ç1v#��Im7h�[�J���%ǯ����PV��]ҫ��[[[s��cO罂.���5�?1311�m� ��p�� @eKKO�����Z2�(A;�S�ƈ�Z�w��m[�v���NQuړ+�/u`�/�B*�k���8��㓗:��4�'�����-��!/ߤ��(M
����z�㔥�FX�o7�T3��@�_Ph�'s�%�!�om��Dc�@�C��ǫCv���a�{��`p��f-�CI))���M��Xz���p�v�rr�"�K�P7x�����p}/��5�����A|S�",��W�Kn�r5����)�r#��������`f7-q!`'i�LAwx a:k��o��C�i��L��l����z��S�pT_�����0>9��,n�߃V��2��S��3�=�f6by�M�o�ђ��MW��U�B���F����w&7L-,���
й��4{�w����t��YnKQ)q����ܦ��@}�ucB�-4�i�E�z�����CQ�^O�A)��	�ؼ��$5ogIiZ�~���J�*$$�t��U�cwwR����Ζ����ww��p�}����c���12q.�uΣUXT�Ġ]@F$����as�T�F�W�H�)��:	~2�B� �'��i\".�+���ٓ+�n{w#8�o���MO&$�*2�L�W���n>�!�[Vl${B[�<�U�|Z�5BQmH�DYg4���Y5���(�&ի�0}eѼ�m���C�rq�̀NP�%eȁ����In�\𰴱����b�r%zw\)w𽥯/##����իm��m--Q z7��P�FFʠ�������/-1 ����1� �A	��V��3�P}����� q_{�xf|\L�* �@6���ai�y�s@�}�3�W�3�$G�+�=�����9�	v�'>-2��eF�D^�.)?{b�K�R���~Y�U����JMtag'i�zkϲ� � 
I�"��� 	!(��d��N���̔���OL\�7�F/m�m�.}�O�I�FI��3���񀬜����PY��r��-���
iS3t���������������SV)��A�i߿ߖ���I"6�d�D-[9����Q��[�u7i,�������mb AP
ޑ�� A��5��/(p�����U��qe����/{����PFb1���s?á�3��逪?B3�ܚ�q���E�@΀a��� �dSK,ȭ�ͨA�YB�I���N�JI
0�~�.�q���4D����l�.��7��GC�5�构�zɏ.o=�>@����R�	~��s7���_�9�i ��Q�6�Wid�\����нw|R��:ghk�$0��@&=T^Mhj�$1s�f` � %Hv|��WfN�o�:��qc�8P��O*�\*��%<1�zh�-��K/((���摲������O
JJװ��l{���X�����P��M_6���o~V�H����B�9t��N tѹ��R��,^�z��Eo P E���׫�dA �ܞ�j�0��C�S�����q�ěb���2{�A ��L
���>uj��;L�l�n���?ܪ�����N@w%�h{�%l.֔�"���Qc:������TT\��X�U�	���m���<�e�fw%�I������JL�c (��M�@�ʿsA�=����婱�@����(���V�M---�zx����� %�Qkj�6��)����۶��U?��d��ٌ4�yAS7�ɑ◕7g�j��Ah��]����X_w������EՈu*l�%��efC<}�"�����:��w���Ia�DYY�/PlX�����/����*�檝澜\2���|���e._���Ù����@�\�Y*�TV�f��{-GLx��c�/f�_�ǵ�߉A�[[�X[D-�:������	ڧk�[�N.5[����屛�+w��x���[^��Z_ y`@��;6�"�9���P��X�i�����޹�^�Δ[:��ikO?�C�2������3a��U?�*�,�r���܆�Ā�M��ųC,J�T���л����}�����_�R��J�)�G]�N#�'q~��G\�<���ee�j�Q���@فcR*�y?1qh����4;��q���91��S!���Ԙ���j屷dd�US�y�/�d�;4&4�[��� ���=pۮ��d�x,p�X{����OBg'S����+#�������	,VA4��ZV�|��bMq5H6��D)VSKC|��,ѭ�4��u��'{��I��.�%L�֚<ƨCo=��E8�����gD�Jc+'�)�^�6���T�繆B�\(׮��ރW��ȃ�TF�LS��� +�T(�m��q���˓1 ���V1e5Y�x�)���Y�����,	�q�:͑��+)!��%}��<?ur�����Ⱦkn�A,A�7���keee4��������P�4\aec�9�ǣ_uYȎW@���P�ںW�}�����v_�v�$���1o[ZF0�z�Ӭ�GG� -�т�u�ϣ޾>I�X�Aw<���&gc��� ��(����?�(Y�Ir�l�ԟ H	���NQ��bQ�wɑ��٧�|�ɒz�p,7@<Cΐ|�w)�S5�TT�:����/�˃~�z��I9���À����A>WU]��6'&�+�3M>]=������ ,[Z�c���׳��>�
�W�.|�����	��|�DG� �
���nI�;H���Y�
ޱ� �k4����oq�D5������/��lF��7n����y��;�oT{�T�;:"��weUS��ۜ�g����յؤZ�Y�l?�����5D�Ԕ3�z�z44I�Z^�Q.����hdUu3O{���7t�	�Uڳӱ���q�����33����9����Ch�i��[eƜD9Q����V�E߼٢١j��J �m�v!�>�����?}X02S+Y�1���w�)(���=�1�����/.�WQQ���g�$�;h�������ttt 7z?}��A%�	i�c��\�ʾ^b$� $��n�}�10���b����Fbe�}��:�%*] 5@
_��d���oX'�'�~?G�b���֖���G�9����&&`OeN� ������L}�ߏ@�3_Dw��앍�N�´�C�`�>/���s&
'�(��+|�/��~�����>i�J	G�zhJg� @�Fi��ç}^�L�n[���:B�:��4��Όb�I11����z�£�r�vP?���������/z����˗���oyv"��e��H��-�����ݟ��8�U5���W������=E%�l�?xfׯ_oJ,	�FYY[�U30L�' ����ٹT
�Z��k�Yu��9IEwVY>}JVf/���%�ܛ�����Y�����4N66oJ�����nY`hN��'�t�z���<{"Q,�?�R���,�"�,���25͗���E�hej\%��z$���'�G9/5L��J���Z\g���$?/�|"�2�tc��Ia6&L�7B��n��}i����)iz�H!���$��o�K��_��/�p����8�:"�t'J�K-=�?�ɒ	D����{��/Ez��g��-7����9ڟ�f()��蟞fO��qE=N�<��GX;��MM��v���;u��
{�������T���]ts���ѭP��v��\�E�֭���a��l�&�{	ż���
+���&��{D�9�nf�y�k�s�en�,L�E��3�S���s�b��{Xl�,pY��Ҥs��.m��)!A�}�
p�غO\��h�;�M��Õ�� �;��+��Y��L 9��u@t˔P�����ם	�8� &$��>R��s|=|DB���R8���cMMMnVJ����
�����6��n�޽S5�ˉ>6<E��5А�Xd�����������7=�GX�ˎ�U��3�*��²�.�|���
)�;E%$�m<>՗�tuI����G�(�0�b[*�x��,��8ċQ��T�$e��fg�H�p�^�a��a+�74��PIR���2e������g��
Nj�K.	�*֠�t�N����1^�)/ϝ&�h� ���ŻȒ���+��󶈳v�ۊ�r��y��˗z?��Xs4/���Ϸ6\������-�mv����ۤ�laЀ;�\.�п�'^V�TXR2Fg�%A���������,�O�;�
=ۧ�G�w~}TЙ�W�qw,����#B�[8�M��8汱1�ZO.��K�����|����Ǟ��E�@a11���vO�&��Ǳ�����p8��A"SCm���	�H�*�~�S�)�@���ރ��f����D���+N����q���w�`��U�w�N~��f���gY�Wp��>B�B?锉��Gwg��̠�S^��<)��~�hӉ��09H�_�6��uv�N)�����<�<��k2�٨���K�A)dN�k'Y�� u�`oY�����x�_��l��1�H]������Q������|�DP֭��������e�iS�n��574$��<��jo�����e�Y1sXz�W�	S�Mm$5�T4�BЬ��RH7pV;S=6���'{p=��q��(���b�C�u�D�g'��I�Ɨ�i���?����^�K���<�0� �c�u:��& '��T�4��i�����EyʏV�I��<��
��v&y���/mA��w��}� �QH�ڻ�-�'��S�~���\J��}��	�̈�ժ�"�AG �k�K�q����4y��[=}��8��]���(�}m�����]�ٍF�����x����A���_º��$��RЌ��`h�D���� ��O�pI����$^�*��R[x1�7z5=2V��v�O�f��<�8D��������K�dsц'��4��>�u��[�w����쪪{~���J������V�r�!��v*��Q0�P��7�F-�O�%V��L�����~/H6fXի�śW�
&66hrds��ʇ���QP��67'BW�9t��̸�O���V�3��N�4�56�WU��cJ
���o��I���ww�+�	v	
",)�n�ޘ����&��� x��)��?�K����ۺ�ip^������������ʺ'm58�[�]6��k��P.�!`]b���D�z'��b^6��,o Q���A	N�$127�s�Ӣst���F��'=~Z�aX=^�n�/�����[-k�������D�\i�\!��:���&%kS�����&ʲE���R��3�p_��&7�F�������?�:͕�2zvv.�V ��UnII�V�Z�:\~��N���"9)������a�/,���	���{������ҫ�kl4��J������lp#U�$͘��mr�C�лP��A>���6���"�cx��Z�OkclH��{�\�deto��`}kկ-h�C]7���9yvu5=c���=3*`ht�{��� <���QB١1�Hp���'�<7�j�NT�{���M�a��Lh"x7P<<�3���в�X`�"�6�S����U�WQ9#�5�c��8)�aHD�v��3}@�1��
�e�J��ױ�#>��!׳��f-�g�h L��XW�_�s�β��ols����̱�v��q߷o	k;a�/0�hy®k�.G:j\\��o\��>�1$b��uo����3gPU�l��?DyvPv�}o�%S��ۮC�yW�4��Yݛ�ݘ��ȝ��X�����i([|��|�d��e��@,(I�߻�']���/EK�$���� �_0f�Lɔ󵇎8����e��-I�<�m8�"�J����L�ͮEG.z�wWwL�
!�_����ʘ�}����i����_$�HS�
	).����xK7������ʼ��yt8F�7���S&�ir�v���7  ��i0���z��B���W�R��)P��r��'t�̅�x?� ��-�w�V���8�����!V��3r�r�k�@
�'.��0��b���0���DDl��1k>��2e8f�+8Q�Z�w���n� f&��߅�M�(=���(��$"��b���IS֎_T�~Y)`!�UK����O����}�f�Ď���b�2Q��p�	��a��k�ݶ�A�u�OwyL@2���EQ�4��>@?��|�ዏWOJ1��%�ݘ����C8�fi �<���_I,O���Ɉ�?�
���3��|�+�ZΆ�����W�>)����
=^���0<�NT/��k/��9B�΍:��o�C�¨���@���!�Q�Pj]�,����D`0?���2�弲�ȝ\q���q�����@
�lT2@8w��]����ZtWJ�h<HK�⥞POE `$���^�ٴ�NL@�6����F)�֜��8���67�'Ǭ�VJ��[�Db�ЌR�|�<�����ӹ�,����7��F[#z��;���I<����`�������N
���kjn��z"�AM<(2H��9 յ�f�~㓋�e���wZtg�/�ҫ6ܜO��s��[���?��O�VA�I5��B:��򼴽ssz��d�M��8yt����G�#:��b�/��???���V��k�|��;��no��P`J�=uu��n��"dɣ���X���}�+��X�O6�+U_�}�����$$*ob�	sMq����k3B"��1���]��PW�Z�re��h�F�_ �.�C�`����f��?>����+��������)0��w�=g�.|6%a-��m0�v62	���!dʺ�8�Ā�9�zZ�/��*�ck�d2��҅�?|�J�+b�t�ɥ)L~1]�&����V^^�S��_�6KUz�����_/�	�s��l������u>��7:�9�Q�a:��⩁^>h�ԇ�^�d𗾷�"�o{[����/�m�/(���Z i$��݈�g`�a�ꪣ��J`��ǋ/8��YՕ����6�6�P�>��ݧd�Y��i����ĉ�@Uox��5�sz@���Eb(�3(��N�e:��k�5�}|������� w�D�)K��gd��Y�Xc�����NO
��K��|��ȸ-�=z����c	����-�T�f�w,VY({��6bD\��u��֏����%z�ּ4��ڵb����������<�`z`趯��w&�	 x�!���z�py@��Y�9�T4�wz�2�t�ui��\,nG��E��⫍�~G��~���j�)5�̳S�̄��ϸ����f�߂gO���1R�O�b?��'B�䪁�i^�{{A-�+M�%3dӀ�I���=x���}��xeۭ_����a��_�7��$��cd\�$�r�LCe����@\�\sH��e���ݶ���;q�܃t��5�4G�"���P�jC((`�t��^gN����n���T�A��ȟ�m��ίc��y�ɍ�#d���ji��w����=!o;:"�x�3Po[[�u��J�S�@�n���?=��w��I2v�ı�zF�;�0a'Х'����JJ3u�=��M��>��@Մn�d�P6��v�&mƶ��?�����˹[��>E�IV��_l��]�?��o�M5���hB!%����Gy�j�.�[��s�MN�8"�~��;�n��G�>�!�I-nτnu>�ݵ<�� ���|i�]��~G{�}}}�;- ���n�,]-	�۽u�(�:9�	�ek2��e�=�p�v����#`GF����O0�kB�P�ݙӫ�9�;����B,ڧ���+[�k�K_K�T�¯B�Y�0���M�c,ޛ���ZA1k����Tv��#��~��aPe�r�0�u�_ۛz;����5o���}����& �k�����Ǉm?�΍���i1�1WU�=PĖ�RP4�m ׍B/E��N���d�zU) �6�7��J	�O��z��~,$���ݗ�&��r�O��C0w�-�N�~��аKA��ݛ;���=O���s](�l&x�vk-22���S�o!tqf˻f���� �.��Q$��uu68��$��"Z�I8�H�}"�M k7�n�8 �Ȍ����	�A7y?|�4՝�d�H�ts�c���M?a)�T���� ����]0�?�N���C ��D��C#s��h�z��9�����S�q\4z)DN�<������ez�q]�l]�i �*���__$NJI���V�MaB4����ؘ?8�L�x]r����ɚJ��1��Z�gI]c_�8���v�{Fed�R�"���Ԍ�2QW�3f���8�����а�yrF�|����I����yYHy�y�A��+��;�Nn���}q�ps��&	������7J����L�~<�/r�b��U�Qss�Ǯ�T��S҈��:w鐣_�b;"Z�<1Ֆ�+I����J	}�_B�onK�l`މ��H�����ye�*%�>y��h�O�'K�'��]<���iexj>'hvY�n�h�<u�'@дw��K�0^CC��~����>�S�?�/WUU�w��-��{�N��,�� �T�����Љ�����/���d� F�2.�}�qnƞ�܁"�u6��a[ޯszS�d����:����`�x7��z�0
����^Ͳ�9�����@��v#�\HD|�@��vs{;� �	�kqqqv' �&_dd��;��Ufi����n0O��[܏�>~�ذ����d��.M�0J��o2O��d�*����_5J5�[̢�Ǫ� �+M���ݻ�U�u���J��&�>�Xizv��g;vJ�3�8nݪ�b�($D��J�yZG{�T�8�z�y�-��?��QLw�.A�쪲�%�0����4�\�9*U;��b
���"��B�њ�b�A�q��^��Z�G_74��$�jKL��R�71��M
8��B�� ��Y�M��������F=���괅��1��i�dj�뺻S�D�Km��Z�Q�\Q��đ\đ
�Z����\�}�3�`R]|���>�Y���h:v-������F<b�R�n��}���gX6
�~����;HA-|���Tm�?c�qh�R��
������W^������E@�I]Y�˛g��9���UU���_�ih�T+��uT�Z����O��,,��i�A�=d���Ƃ��o��{��j��� yz�}����D�"Wc |0��
��������������w8��������3+/�F�.Բ��zS��s���#J��%#Cf��"����Wm*��y�v���3A�.ǹ8�5���貆�)�X��ܱɰ�rۿ�|HT�Q�M����
��������!���MX�k, ^y�M�/�L�����`l�\����v�E��.{Ab�k>_��/���0����%>�Bݤ��uv������"/�
 �FԀ:y�#G��v'A���"����s?�}���Q��*Wc��u�YN�WK���R����xQQa���d2�ځl&�T&��P�<�k�{9��򧒅#�|���k���Pκ�2L}`p��0��B= (�P����Z������M����*9��-�ƵQ�
>�k����MQf�ܱ����u��d��'i����iw�`��J���b3W����iAa��.cy#�UJ��5�^��P���x�˴�H [��KXBDE�ތ�<�J�$d�ݧKmFj�N e����,�A�('�������_)�<	��!U���w����~nKe$�����Yc X�h%���7iO�U�E�%��-W|��r�.���#�`I�#y����g~�{{Cg��ꥱ)P�}�.B�c׀whh*Ѣ��z�)%��?r�0�ڲ#�'*@����)����0�
��p��E�p�ף�����ax�(��P�1�NA�aU��)̸o�����׺��h}|}[^�:w�����d��[��2�M�:#/�+Sѳ�4�d��=׸���:ć�C�5$����gO�&>R�]E���e=���[��f���8x�a����P�3
=�E��G�ȑ-S�5��hR�7��ӝAQ䫟H"�M�I��7��\�G��z�nPQ�ç�d�i&z�mc/�3>&rK�ӲE����y��X>����)ӄts���D��u�sH�߯-������v�8� �:W���W�.��j�ta�K�oe���0 �  o)'1Y�fFV5_�s�?�y����og5�u������!!=M.���9H���'���l�eݎ��<k���U�3�	3��\�����w�$B�Te��c9N��~|Zsi:!0p����9)����N��x{��2�ǫ�����_��d��! � )B���@���/������3�Q�V�m��q�!a��5QkiM8 3�\_��ˁ���"�LM#x�c��==3���.&��|���(|����]g��r�9�]��Z7�
�S���/�6a�N�Τ��LO���1r��.�\�%�z��L��fl ��wl,F��5]�>3x�M��rWUM
�%y��Sg�W�����d�O��:���	c���E@q�T�in���K��&�~��?~��k (�Om%��sˊ'�^b��u�	��{	,��?IvL�G+���pn�������a:V�����K�<��5��.�X1����Kj�s��]���󚚙�f�+^? #C;ό������?�z���L�����J���2���͒����E~v<*Q) !�	�#�h����utX=�֟p��iuˡ5@ii�G�>>	H$�EZ��Ť�Ěm4K㪓ӛM�5�m��ý=q��}�l����T�������o��v�Bv:��Na�P�:�xŴ�[u�;���3W�EP�_����pJ��~�9��X�Fw"��藍a�Ǭ���&�Ĥ�����%�?'�Tֶ�ce��I��^ON��{�av{[�����'���5�Ӯ�ڒz���	$��h=��M͍p����������2����ne��]�vr�ů�Z�v�~�,��w?����q�*'D�K`�mm�̸�si�YL[��ͽJ���̻#<BN����`	�
?Wpf��D��|P~��N�a"��-��n�V@'��5��[7!��ϳڝ������4���J{f@� �ـ.D���j�&g��n����&VU��,�F�g��ݴ����0.�r�xH"\rm��[m�d�y�a�G�����C-��q���ݑ��7���YXx�.{X�źZ|X�wq��E�#_�n������/�_G�����U�ۀ�~`�(��.��蜎���1Κ��4���x*�T�:]Ġ6������<�,k�kq���$��P�l	q��OB�e�|JnFh儓��k���4{���VJv||\��mk�3@����WV�A�?ceZZ��m�ԎCk���B���W�]O=@Y���t�1>)��uHt�R�_b,z�.�L�C|�r)�����9����gɄz*���8y�x�W;V�P/G@X8y�~��c��rJ�<?������2��n7���d;c�2)�H����@|.�W	��#��\�۾�t�4�D�:ĕ���;m��}�a�b܏�Ird�%SQȘ�1r��(8���Iw)0!�P\�9���e궡�5*��9''#ּi._u��z�y��P6�~HDY��\Dv��3s�_�Y]M�4M��
;�?�P�V���M	F�]�*��g�խ^��1׶��5A�������8Ug���I�ŷM5浳;8�b�|5I��~�?��Sp;�c��_���^j��K�F�Ts<�6|�܌Zd�v^����o��3���:�n�e� ���HЋ��"I_ 9'g"%k`�{p \|.��r�Z:�g8�Vˈ���ρ4�=�Z�Q�/$>>9�b��v�]�	N�02�	H��������,g!�1�� ��\�%�i �T�ù���^M��SS#Ħ��#��\���-9��A�2��5ZM#�cE���/����� �Kb�8�69ф��+�nL���GF٨d�? �*ȇ�XC�|ӏ01�GJ������I����b�<3	Pf�����|�--�ͺ}l����N�-��G��VU�
������F��+&��ԙr뙶����s�*
���3q��Pc,;�NcQ����㖧�5�Hd����M-��k�����Tb�kMo����i�	�i)s=Z��:�]W�ެ�e�C#����k��Ϲ9B������+"��E�Tо7�y規U�ZFOO��A^U��:Uu���(��<N���MR��`����_��¬��?!_�~�lV���n�����1�����؅�X�s����L�?���+�7E��O����?�GN��7g5�X%BSq#Z�����p�o��Hn琋$F���|B�;
i��2��qNG��:x���!v�.�ʤJJ׀.��Q<%ԛ��E�x|�|��N�H�%��Ӧ���%EH��T���Ta11 S�7�Ą�n�X>}z�ڰ�����+���>�3N�uMM��ޜ�Ԧ��(o����l����-�}6�a��';����j	P1Z[[�e��70�b�f3g��v��:9҈Ny����?I2]1@�X����L�?���������9K]�gH��Ot����Ψ!@Fn�x"���A?M�����q�f���'Ͻ��|lcC��x�/�������m����)�ay�Ӄ��6��H��/+ �֫�R�IV!rt�m�"�F�
~Se�	���.Tڽ� yI��om�/8�zn�]E��C�����(o*��;k�9;���@>��G8)��hh��w��[V�]�����Q��HUV"�k��`�U�O������iNU"yZ��Q�Dpr���CVIf>;0h5U�V�~g�i��K�K\�}�[3��]����m��i�-c��Eؓ�LQF��f��oQ;����AJ��Aj�|�߿�xN������"ŉ1)�m4(�[Ԓ3��Cx��8H�����
'q��g-�	���OAV��Ul�pE�ab�5�K�,[�48%���و���H==�N$@!S�,\�M	?�~>^?��n�Euiv��?g`@w��~/:�8�+uU��d�V�4��D>u�	�o^F�LM5�7A!!l�X�~��ۮ��Gk����s���# ��P��bY4�����Smp��g��4yU��]Oy*������(f]�{m5����ed����2-����u�z6*N�:�.��t��p^3�Q�n�^�3����.7VS[��{@vS!�45��W��}��,��)����o7 �9�z	��,,ϖ#�����[ҡ]Q��U��_��f��b\@6���*�F&���⒓���Y�#8��H|�}����������˰��/�zQg�'� �b±�ҕ񂢢P��[�ǌ@�f��w�7'ɇ��~�6x,�T�F�&���n�z��<��	 �+f=��5H}7O���y�R���Yuq���ܖ�ְ[pp�Cc���8K*�'ɩ\�/-��tY�q������7Ƈ�>h��s1�ӈ�l"�(H��R|��{�󳡶k�)�3ѕ��-���_i�bƁu	6�o����Ʈ�o�VlUlnݹݰ�������������T7�$}�KS.�;�q����S`4�˒�C-�ZZ[�zzdѺ�OM���g��3�D/y���������@:`��]�޵�����|�������M�?D���x�>|$�;��r(�������M��7���B��	�Ma��Б�����5I���ֻ�l�-E��[�t�-����Io �G+���?���KM���0����r�bx���Ðh���8�OK���JԿ:������^��D��ΑDx=��%�$� ?9��W�E^^���H��,�U�D\]��I���XZL���l���P����<x��EQ���8���v$�5���c˞��G{�D	�Bs�̌��$��t���Cg-:�'�����$�w�������1��(�@<$,��S�4:�H��O��'v�V�=sB/��p���,�p��L� N��#k>@E�h��j���sH޳�wN��D+�R��	A@P�.���Bж�5���?�a���r�hZZ[�a��mTU�荥��3��V���&q���sgr��~��7��\�K�X#33�cV�E{��]c��U�*�b͚�O._:t���@��������}��f��2{h�ÿ���Xk|��<��z�t�ʁ)O�s��EV6*n��<A����W7O�AQ�-�����gc�܌U.�@������/�"t��"�|M�Hq���	t�����;�����U���{%$I�$3\3#��M���2CٲB!d%d�nH>�n�^)ܐ������;���sΧ�_���1������Q���5�!�ӿDI�k��(�<�u�l%{dR�@�k wv��e�,�y�|�Gmln�9K��#���ё?�9��V�G�.J$�;#�����N �U��	 50�x�93oؿ�Y^S��1����O�9������ݜG�P�z�V�CxK����%؞�-����Ѿ�cI��II���'��� �8}t�r��Aj
����p �g�cZ�A�J���봵�',�%"ۏ2���4:6��4�?h�w���!���U��+��:�*|��o�d�~z�|wbU �};$9�t6n��������O�Ngo��N�����E��M�������&�r��d4Wrӯ;)���n	�R�Q(m�;��ڴ�K{�a瑱<�g~�*+,�>!�u�.|���0�b�`��B��C�m�dzd�`j�<��9�om��w3;�xbbW��]f��T����g�i�J|��)�B�L�@��1���8�'ov�l nq�4�g/85�B��Me_�R?�9.���7�i�fp�Ε}���<�mNW���-2�Q?1��n�)��������w�y�� ]m^^^R3�\��H���0���>��`�}u%���ekP�!�R�Ӗx���|��o�$l?a�� ���m"{?
�ݤ.7`���+W�"/�XqՇr
t@�qS�n���,�7z��2�5���*�3�  M���u�G�z=$��g��vg�Hv���c�a� ��O�<���T"22!����ܾ[( �0��g���֯���D.[��ȷ�W��buea ���a.bktG8��ݽ�A�
�@���1jd��6MmJ��{����hpe���dʒN�C���Ы�b�F:ѫዪ9fyvF�Ȭi�ɷ�	 ��֭���Ȝ�)�??�<������uq�u�����m?�^�����G�W$��~�=�v�UM�*�#--e��v�����~�_,Sc����,K{]�E��nD7
u]����;�I2v��%�eNO����� &x|\8�P�vv����I,rqwl���E*?9�6Y�� 0TS��Ҹ<�&S��I�Ɠ 0r�sH�gyJfv���,�e#����;&��X��eȠ7��agdp~�r,1$,�Z�W�߀!��WU�kϬ��:�I�Sn�؂�4����ME�$��Z�|dZ��rK�~wãQ ��$�yZ��������\TX2�.�X�:/���I �8ھ��G��W&�N�:/.5+���v�oo�H�\zK�^J�y��h~B�ϟ?5q�{��dh���K�o���������aQn!U�4B+���_=�+��U=����9����EHkF�*�ٞr��\��KO��1���_ݏ>�SnS �v��\�0J�R��"E*�o?H**x��������?�E5��S��!�M~�#�$;3���g�����L�6� �������ָ�g�8�ƆG'�?��0̦��k�F�7:��i̡OCBdt����U�SX�����N=9
KWu���P�e��m��P΍��%�w��׌����:�~K�LI����g������x��y&Ck�yt�}�0ir��Se�׺��Uޫ�	b,��w�1{�����nJ��k8��J�}�k�gC�5�﫾S��k����H��p�W�[�(�F�������~�� U���!��۪��J�Փ���x�v�c��s�l������Lul�g ���N֌`+ߌ,�;;w��D=ԽLɕ������j#ɦJ���_���m{%,��޺��8�	|b�j�9��^F�l0b����|�y0��H�V"�-]�N=t�t<�� �^�-]�P��T��,Sߥ�kM���F�ǯQ����=�Γ���D�mZ�R�L�z�J�RZ
��/LDq����}*�ぶh�������9���N��m���/@�T�We����"/������@N(����Ҳ���>��l��y��X=���tɓ�x� �'�))���8� �{�G��4��q���l[�A��)y��̾��A�ZW>�XH���EA�$/���R-��X툚�1�����l��l� ������s�f�0�L2��� "�K�4_G�P�;:׌ � ���T�{z/�����n��_��֮=��i5>`5_�{q���g١�Hp���ל�V�76{�����ɞ$yf^9ՌT*�<k)�ci����ǓZ�9M,���^/9���x7�@`C�fc� )ҙmiiɜ�>f�c�e9Q���؂��/	�gh"�����D5�qZ�&7O�q_Oxl-aS��k���f ����oO/��{s���$����� �<�T��mdnęH����BNv	�
�?�����}�j�N�404l�ￒ<��v߼{�	,��R��*��;���1Tw��B��W5��O����c��,�o��u)n�z�:s�F��^�{cN�ڄ�����u�@�F� �2s�K�LW��d���*�9;XI. �*�1��/�W� �m-�<n��%4���H[˦)^5�r�w�ܚ�����(�fg?�M���!N�1�/���v �>���B^����d}&߽�$������6ֲ�u��:5G��� �n�%e\�+�"P�y��vوt��/\-��*�0�6��Izzy}�wwD4�R�%:��RRR�<}A�F��L�g'�y�c��4��Ȝ-�P��q�<>h�
w^�y�_�;_��]Mu�`�����uk�YRz�4�\V�"�������S!�W�2{T��ru:{zȁƎ�Oĸ��wς P�����_���G֢�����'��gs��Ą���	������y>�Oy�>�lV9�aLxc�SG��u��mEE��~�����(t����#c�|7�{��	� �JC�#�����}ԉn�/�JA��DN�����JI4�W(����c��A�OO����ڱ�L�)�'
�ؔ�g�`���jӧ�T5��x,�PW�aLŲXǊ�m4]��uD�9� p��[�٦������Y�l�ҿ�* 4�A^A�:.51m\���T��O�)�V��YZz���z�-�Nك�}���[4X,6��LJj��S�����扷��6;w���83�I)�Ǔ Z�[Qt.rGc9F �輦�HA�J��n���B���/"d��+!JR5����ࠟEȜ�e���)�ˋ������H����#5�m��LL:eY΄�A�zIf��&��2~���������k��*S����CBv�����6�o���A�N���N$ob�Ջ�����������j�'�����s���<d��X��s7���S0�E_2L��^�}��GF����w���u��^�xWT8Hh�L�+�ã�����F�~��D�r\�o�6�t�b�D��٢'�����w+(��|�^�G��~�X$��a{|�G��*ێ�ﶴ[���p�<W�2�D8zE���� ]�a���婀�`��b�>
���*�V�Y\������\�o�r�����x��w����NMq{=g}���#%>ʧGBAAQ{#�V���s�t���ŋ_7L��i;W0��?{n��|䴜(�������2]{{/c�x�*��s���C�/Gy�A����%�Jj��3f�ra�ü3�Cn���V�sTT�Ѩ���4K#�q����l�P��e�e���1��s�F���U��9F��ϻ�xn�\��|@-$�vB5~����}x C�a����b�,,��e��m�KR�(�*���646~X\�!�m�c�䔽l�5gZjc�㫏}�r߻Շ����y��x�O�"�Q��H�'�]�ep�x`�k
9��������������U���y<�4��Ī�1��Ҧ�,�I7&�J ���}+��s�ė���Ռ��4�[�� �v�[���d��9i�̹&ɋ�|��TȻ�s�K���b���R*X���265%��?Kw��ʊ6G m����o烠kD����y7��y�#R�is�o`v�ɼ?�a�a��a�<�I|��L����8��r��)@f �j�'4�%���+�����o@?D5#ǲz�Roƕ.JI�ț̬x������<S�`��D�w���5.�9�z9ǜ.�l���r�8RIpf�B�������������N�����	�~��͸��ѿ��UUc�>_c+�ȴ���;�-
5}���EϷ�4o�WWF��>���<�H�[���uO�I��n8К��h��SBʿh��o�9�v�5h��?>M��/���?�\<�p���/�k���m����d}5C������k�^s!F�$����0+�T�'�}.]�|�E�~q�g�̟���h:�@ٰ�*���5_�(cQ�f���d!Q��8MM+����C��^��E�q��&���5fw�\n	һz{�*�Y9yx�]k}�������zڅ��ׁ�Y�����+%��9q���A:g��e���e��Z�W�a��b隠��E�W~�YK"=A�_� �s)���e���nRbG �[8��)4�]�9 �x׏��F�TR�ޓ�^��QCJ��T_$/��6²			�{x�#m�d�\Q���������U���/�C���]H;�ݩ�##S��*��-�B��>8_߆�=��66���ؼ�j�yyr�K=��ov���9^��9Q��=�_��i����ν)�Du*U��"� CT�U�2E��J(���E��2�ْ9���=�-s�N��b{j��i��H�B�
nn����+f�sK����4װ����#�����-�QQ�߽���e[�ջ���S�k.�����T�enl�tv��Q�� ��:��-��8`~���͜�������y7�������%���A��6��*�=+e�W�0�6�Ry���e��>�>=�8����0��kb���[�QiЖ�Z��6*EF���}����C���PG�;nnoj�&=
V=S.��1�z�Ї��{�ccn��Ky�"��eqӝ��?c���� ��=�8�B�[���i�zԽ�݌vـ�G8\����g/��H��殦�Ȣ�x�.G)��˽��֚���yԁVA�r��el�6K@M]�DĮ��[�8�u���9�Z�����]M�]�2fBY	���Kӕ��nm�9�ėX}�}�:��af3���U���8�2���j�VH;D�zg�1$�I���A���ʥ�OF/��ܢQҡ�@#����i��(�4�M�9^�4H/��Q7[�X]$�!U�n��gLĢ$n��ܹ&ԝ� ��t�jgz�[��ϟ�yIxU�\w���my���^ǶࠐPwnR��[O���_��PPs�̝s��������9�i1"%1g ��P��m*8�#�a���gyKԇ?�:^��;Ҳ�(�i-�(�pK��z�� ��Ksi̓���C�F>aR�����|�P+�O|ӯ��1 y.����j4�hT*.���{B�# $�><��C7;��~�B6��=<2H$wN�>��#�?���J��5:4��G�E
��C��E�� ��I�����4�R)))EI�{��d����\$D�h���������=��=�ǫ��x|sBj1%��ZhmP�"L�G�)��N��./<$��]{��t��C֡T_�>�B���K��Zt��������YH���:�"=犟5�Nh�Z(�����@�{{G�oߦ�@s�Qf���r	��9�
h�z5C����3 )e󍅭��(���σ����c��4�5���k;��X,�V�M�>EH��m��͹n�&D�����G���q��7�ϥP@��AyO��H�h�9֌l-5�)ր`��}���7�;8��2u��RV٩��KbL�=�)!-=9q�\�����p�~�4����e�|(M�k� �e�\,1�>>���Q,����$3B-��}TY��_\��A���ҕ+�[��-w�غ���H k����6J�4����7#*#ceGM�_o_��kv�Q��5NR�R��=�\��a!UK v�����Q6���� S.����{�I�	;qV�*�����*OD7�SB٣�A�M��M�����V��#��7��s�\�_��p�^5d��X�\�Ƹ66$�)���Q��h���ZB�z���z$���A���QFbSW[��d��IͻZ��ݵ5aaaP8�G��_���S���$�����[?9&B�>�o��=����<==���Qዽ�e�]{�t����������:t��L�u�q���#:�����1'��G��>�}�B�j�n�	��� �=�3R����a ������υ�U�n͹K:��d�y6|�u�h-J��R���xb�sm�,��KW|��%�}�*0p�Y��e����@�r��0J����c��}�s�gg���~/�olz���
{�T1t�E�[+g���C_��L�v�V����w/+�˥�h_��������4J��5��*��������w�ZB�<f��;���X��!mTH�>�^�k.���(��������7�7-w�@5��ǿ���#>Rn@���@�H(gB&��"OV��4@�ic������.;i~AW��º$f�>���A.߾�b�����Z�k����NH�G/�H֌�,.���ArK��ؘ|e����> Q�f���>s�o�(j�C�TyW��s�Ld�:a1�S6���R z��￮m�������^H5�%��B����
z���c-��-'�r7;��G�o�Uv��	7�����*�ں:7�lĿᗝ�*l/�-���)�᝴ް	��˷�2��>�zP�|�� �l�	@y�X��}�Gi��KK���"TU��!m�ޥ�p��4ܡ��m�d�{�Id�����Ş1-�!R��~����$9�}-|�:@���a��c�aM!�s�^*]�Wn��Z�R)�����#@O�L��a)�Ť�qx�_�,Ss�Q�zʅx~��`F�؛�n��=U�?���<��E����o�\����y&��Ũ*�
?.���N���������+Fy*���c�y/�Ȧ��Yq�[[�E��Ѫ�÷����U�I��u��P� ����s����ES�����9U�'�M:��.����٤4�zђ��u[+��G��v��� ���fz�Z ���T��@yK_Ň�4YQ�F���]Z�=Bf���~-��op}x�<ћ)SӘ�rp�A$~��x"T?|��43cFP�W)���X��da���7er33��"dܾ[~�ڽ`�>-����f?R6����L�ES?���ݾP�c�oO�����c�㬻$R�5��ܳ!&$DF�;���B���泞��mmr|��bY�AWFK�*(f
�>��=�ҟ��.,��i�Z��)�A<�\�$�$�+A��~�G�(�DA�4�:�J"��k';�@�0��R��TFF7���$���]�"<GW=��;���2�F%^k�M�̻�#|s�<2�$���oi
y*���'��h�H��yb`4C6����b�H�Nii��@n��ܿfQ���}x�A��F��{Ș���T�}�3'KJJ��~! �M�����]<7�B!ޫh"x�� 
aD\\]����r:�y�������<T��=�n���	�S=�Κ�G&��p9��U�u�#���7�brk�*U�#�%���~���X�������X�[�5���|�ds��n��p���t�xr�?,zZ�۳tYۛ'^�ʠ�:/elf�;�D��R�Xy��aN�&&ӿӦ�r�=c|�gq֍��W��'�z�
�o`��D�x���(��GB��J���8��oR�OI��!�82�2��!�k7<����9ɩ'�	]����Ty��z@}�$}^s��k�y��컦��W9��7 ֢v��=  ��[��J:ߩ4�EɎ�(��ۄ ��]	Cs�R*R�Nf5���0����sp�Ё� +{�-�Ħ:s�θchHVe t[�%�[��}J?}DL� 	Fy�-F��4�$RL-��>*�ы��1q���jtRAq#@����ne	���z�,�Y�BiJU�C���p�����1�v�� ����O�Ɛ��~v�f�L���eh������y����s6�ڟ*3�`h﷥Sg��t=U"�*f�.X|���oF5��h��=+1n�s��*_bx�L�C��"�$�Cx�\�b$8i",�	"sd��l''�9c��ûl�!N\��~Gq������8IZ��~�=�m���%�Ɏ�v��=�VW���W��vV��lXqqw�X��W��>|�G19Y(�]J��ec�r"��KH�W��b�P4{��y�Ч��Q.��T��3
E�,i=��'�� � k�E�(�򬌅�<��lA�*º����)�����Q^��Ł�f��e]YFrĞ�|�)��n�43����#3�����uY���%�Y�
&''��peh�L��F�r��ǐ�Ώ���,.CD\".)s��4�3�U�xe������3��	���'!wh-��Z�+�e�h�.�$�\
�@�īv�&��)axg�4��T����O���q}��q�g{/������3e��>��^;;�tE�̛7®�'C-��1ǋ�$�b/æK�v�hѓH��<� ��:�$s�*E�������'��^F�?�a��:l�ӊ���v��z�#�s��q��R�����ݷ�Rl2�����{�	kB��Pc+�|�T�0DɃ�^	Vlo�������b����7��P�'����k�E;�O��{r�o��4G�Z^PS�ݩ�w��o��:O��5Uoj.544�\���I��l���n��HV?��ə3���"�CG�!"&6v{5��^��M)ᶏ�:h	6y�T�C��͆��B��~{�߮����>��k~s�9����ȧI��5��hWuu�X��߿g�G�[�]Y�.t����M�Q��1r�q/���ĺ���׳F��L,zZh � ����9�a@kԉ�y�睏n�v�EEӻˁ!6�v�Dw��!����,^��_�
"O���:�X�]T$!#3%>�҇���)�cP��.�8D����Fˬ�r� �%ؔ�3�!ӓ��R���Gꅖ�Z�<�<���C��4�R���w�������M���\�m���B�^M��r�q��jN�@�����ͷK|à%��7d"�SX���	�?�`��3r��ǖ6��� c��-1-�	,q�>$�2���;�H� �}U�\>5��P,���pF3f~���	���pUk�� �r�x��p�U�u���G׸yKyK	����?Vy����T#�����8�3���i�9W�T;Kvzgg����$���hŷ�q��?Kcw��.��V��͜�E��.6ʷh�!:��`��M*b̔�P��"��2ҩ��pv���a򡜞^` R����������'�w�^�9O��i8x�7w�T��9��{�/=Z睟Fq���>n�����2���=;���ަ��C��g������L�W��|��������(�&?����ɮۓ��T��4���%��n���8��-����E�Va���?�{b,<R��<�]������&T��� il�Hz����[;:�rtVO/7��?D��L�λ��_�[�5�����sx�>O�P;%��n�����v�(O<)�wN��Y�D�|��T�'
�,T��\�G��&)5]>��A�g4+�%N��S�A�٢]�)�'8���Z�΁������wD9cNV�~] � ﲽQB��qj��y+(����	�:�C����}�� i�gC�K+k.�Zh�I.C�V �o���H#e������888��{��E��/zά㮸H��>J��95uĭ��J6���f"���O�������)�S��-:�B��������lP���q�Jf�Sǵ<�y�����O�Vb��z�Id�b�h�A���|
l�>�MX#ˉl���U�(-�xd��/�=��7�.�Ą"ύ����A4H4s����hí�Hv�j%��7�t�������O��{���5�z����` uδ]��;���;0_���&�g�z-����%~�Y��q%����TĖ�ϻ�f��>y��٠�/���z��}ґ��V;�����r̵�����������Q@@�C�"�y��BUTē���_g̱5CK"i`�44tϟ}о��ۻubL�c�pZ��aO�q�B�E��/o"ۓ��Q�9q�Χ!�V�N꘿!��ʊN/�<
#bI���LN�) t3�.���8��Ku@6�5�#C�u"�=}�/��!Js���S��{@z��y�A�K��a���i⯬�!��H5`5dB�zV	��,�_��	2���</���ےC�=��Dx\���c�9+����˾&��m]]�����ѯx-.v�"^���u��f6
~�N$2~6H���~0I���Z���yņ�?�H-,I}�IIdΞ��Ӧ�bO����<�_�/���� �x�ÙF��V6��I��Gয়:\��G�i����tTU�Q�Sj�.OMj~�Pe$!)�j�VBi#�\��vQ,���\��tsg�fcD���)���>�6�`y	�{��h�LT�[]��Őc�f3*>��δ�(�w=��^J��	�u�މ&�X_����s��ǃe-��ς�cd���TB�l-*>�Դljm�ս.Rv�H0�~�y���!w�X��sN׿iaF�d��
%On�N�x�\e����L��|�KW`�*S�a�l�B�г8���Sǿ��c��5�V�IR/�H=O��3t�Q<�������\Xa�������S�-n��\��B�K��IP��m� �&Щ��n�Ik��*�����fV�J\}�����/ڋ~�+@�7��Z���YO��便�����c��<vuuM,$`�1r���T��O7����q�$]S.�NN/�2s���7dd�A|ԀmwƟ��9�zI
8kA���B \j4���e�y|Ȍ���Zc����+a	�\��}>���~�T�������i�D,1��\4'�B/���}�{�����Y-/���u�H��0�Ú/�n�ꨈ�+Av�T^}���BQ����v7���y�����W[i�RI^�Y�:= 򷕫O�i?�G�5�nʠbxi4� �HIz˿���A^�#/+<L��M,tl'<�4���7�Í�!T�1��'??�MTÆ&�����P������b��CflU}�Վȷ쾡G�}��_�`6��Ў)�m�L��dP�l0�땫�����Ӧ9��`"�;�"�֢O��k
+��j0$�<O"��!��S�޾�s�ϖ̴����7}1�����?��NI�7�<&{��W�Ξ���>���d�tl��\�ׅ.\��?��r��Q�ԉ� uP�~vF���fcN���h�j@ �ܧ���0����؉c��n�~�7@��MJ=��t�9opm:'�yXn��SݹS��z��YGW��:���g\y��;�R����	�D\Kq1.��s�$I���S典jl�����%��0� ���n��R��k�w��m�`U�`s�3�	��~�3��ٯ�x���G/���&����vv�/��z�n�0~���m͈��RH���Ej`h�;���,"����R�.y�;�������5�Ҷ6��C	�4Jհ�{�����$(xk�GH*\�l����ec��W�b�����FZ�Jj���ʚYX8E��>�z��x�-2h&^�8Gb4FP��
����.շ�HQ��l�>���"��x�-��a���?G��k!a��*=,�oo�HM�Eu噒��^s��1w�����Inv�}J��꾪:$Y#_�i��|=r`�.�F���!�h�7.9��1�"�߬
�Q�P"�ҡ�_�UF������XGU��W�����uf�/f��?��[^�PzM�H!��އ�O[��Q�go��x�Q��2�T��t��鯤[,�r�$�>,"7���i�,ˁ��(oﯸ�_`�C^�s��WINՌ����#::4a��P���������rW��k�k=%W�qd�����\����WMmC�"r�����:�v����^���2�Ts����GAlQE�k���y�V���3�I���B���3kkt~�Y|�γ�z�1S�Oo��sʾ Zg�C��*��d��������-���M�E�*M���
�_(i�1�W�eukF���}���UK_��y�x�t�)=ނ	9�����e�0�����s#5oب4rl�]�F��p��eo�Y�]�v�%t{��j]�������l`Z.�o���-��7YW�)u�L���\������f������(hPd���Eů�P�8��Z�k��A+�ޞ�[X6s��xK`�Vvt�u�[iX=���;�]��0�u�p�Je�5�R�`�b����oC�cD=6���y��2���;���=��P�u�,7EY��~��x�����U>�o���/�5W�#�7*�k���������U	�awo�T�q�=D�+��7Ǘ�s���=y�|h�ݳ�-ON��)+-��̌�+��;��=bb.t'��ݖ��ܼZ�zQah��E�W�TJк2������Ӡ�@��K��T���ہ����:�={
�Y��17E,�xb��0U��lxg;Ǣ�Gs��QXC�3�{5Q�9�G*+{�H�M����ÖG�G�(���p���
"}�;�ǅ{{�tŞ���c�
����>��9�O����>�^K�+�����E�����nHL�`x@�&ҽ�`mxТ�����K���-�t~˔z��ݨ�w��3�W��]>��y;nu���e^:w����ΉrEZ�u��K�<�9�>	P[��ޛ����|�'ǈ�(��lq�q�2�����O� %>*'V����r�E?��Zv�
A�񴂲OȨ���u�]�7��S��햮�]��]Ѱ9�!D)�y�i#uL�4�C����|o��	�����p��W��ǎ݇G6�Gf��<4�U=�r�)��+&"��O����4;�l�H�D���BĴ���ciW�i���׉
�x����������g�w��ߟ|���E8�y�*��e��b��mQ|���nT�2u�/N-�8��DV/e��AV'���"�\}(He?�0?��U/��h��{{{!���*�_�h��~��? �X�s�����4���!W�����K,��o���dc4����]�o�s��l����mFDs��+����{�p����e�
�������FZ�x�>Ř��V��$Z���0I���Hѕtr��o�-D캦�<O� Wf,<{�l�:���KQ�2����kT:�ݳ�yx;��q���<���v��5�ޗ���=6C9�C��"o�p�Ցa����i/�}��Ἳ��NfO��P�`Zj�@��S��� l��3ٓ�|�i)t�������� Dy$�����|�)������2��	.mB��u���ۙ)t�#=����O�<F��S�64�Vz�+�/]�r�P���pJA���&Z7��G�x\����H��2~��IX�&��Gם�TѧhTI����KR�F$�n{�ܫ��&8h���j��I��H�C҈��a�P����bKs���~���F?ۑ^5���*V��uI�+r���2�K�����n�R���w5}1�O���˛g�a���/o�4z��5H9o�>~=�&���,��Px��� o��2�E�Q��G�nRo�qxyyk�X��p��EZ\�wɊg4�OM�/̎:]�����Jn+މ:��������w�Iꖁ�e�
�_�4�^o�X��n�
����`m����(��2�H&�p/얻��ȺϾܼ'0R W��x�/eV���&������?�f=��۷��aD�VUE(L5������U%�]�+8=9IDI�D<�̂vE	՟3T��)Ar�W�1x�M:z��k��M���1=n��ѱ���|P7+W��ip�����o�Uo~r/�ū"ss���i������w����_�V��m8�-,Ш��L����뚠���'&��+���yΫ��@mz�z���Ąb��ڛ����{�{�����|s�5L^~L�� NZ�f�a��]i�^J�I6NN.��nd(������|d���:� @��o��ze�+��
@Q�������:��!A�����/\�;�M#��I )Ҍ�)E��7�cE��+;��Q'�F��_�9"�m�����J� _D����u�N�E���*?j�����;�W���qJL���♖���ݠ�Τʨ�9`�����tQT������~=l���)�+^0(�&�g�:������̏��e�Q�i��c ��Ҙ�G��� 5�mn9��FY99Qx�~������:��ӛx���xc�֖�Q�Y�B�?��#KKO����)���u���m(�#�R��}/}	ZEW0`yZj��īu�3��6��ܱ�u{?��!5|;�n6x�����vM�v��5������=ы�?.rTs�$�W�c_Ot����)��il���T���]]�^ƾ��"�;�w� ���nD����ؕ�Ţ�kj�aD2K��e�p�U��i;��:���gM���Ź$-��$�Jku�⩺^��3�$1��Bl�?��z���d*$$��^��(���hۢX�*� 6�;g@���s�u-�_�V�2R�Rg|��W����߳MB��I��I��S��ȝ;��)�ߊ�v�L�)@w���E1�wm�I�b¸��͚fW+�t���
Q�Ǐ����)���O$�4��#9�3d���Kg�#z��
{5����G����DPQ�Sh�0�	#��ߵʄ����%�j�D� ���2����s�N�~�`0����$}�.]���U��z���t�[�9m�\$��p�����L,�?UԿ���X�ۂz�;_{U�
�GR��`�k�.{���]q[�!૷���}ۋI��J�N�Y�S!d��v*111��@�%�w��}ԥK���w��R��� f���W�kk�HP[�{��rpU~�����D�����'we�;�z�4�N��F ��g��$�D�@�-�ȁF�*���+�6"W��s�ĄM@t{n\�_|N[�+/.����Dn��H�%��Fw������m�?�ϑ
!n �z_���fN����e|�E��&��#��X�(ص
h�aV����Ǧ\��rb8����8���ъ����0OS���&��!����ܡ���`҇�j/J�؆��>7+I�:�����ss�Oό$ugSFK[���u<H�M����Ύ9-�CJ}�m,Q�,ӡ=��u�+�%D��p��(�_��k�T#w�c��?�b�� �i�3֯������c���y��꾖�>/+��o!������S;;�

�E4�\�|�"s��<�c���%�ʅ��J�����:�/����L?WOb2�m�3ر�x���~�mK'�B.�W�������r^[���o�����D���XkÎ�i��ץ;>MOKKc��3-��Q�m�ec���k�����y�k��F7ve��A5Ci�&X%�k-u��H��.iEE���N6�8�UK@��ܰ}m�{$��I~��󼻅��1ᔦ�N��G���Z
�8�<N���P1���/�Z[#.��	��TXݞ\ߙ\��>�V�ks��)����Wo`���J���Dk[ݿs�_^��u��l;I�fH�~u�~����P��}�]���.J���g�J��� ϞR}���'��\a��)�-�<��Oy]��/F|�ȝu�JH����/���tt}79@���Ni��`(;A�;�����V���|����"�O�i?[&�raF�@L$�W��!����h�-�?b_=�q�exD��ۂ���(�F��]�M�[�IE%+M�ڙ��3ݢx���X���\<�y��<�FĂ����W���y�Ju4��}E�_�9��i�c�ַ}�"��%�,�H���ʝ��e�̹�|�c��^�Z���Ž�IT�\;2E����w�D��ӳ��"�X����!
�	W����T�B�`@0�~J�YG� t���Q{~
'.�&Ǚ��r��w]]]��7�s����_"]�z	/zץ�$[0V��9؉�L��n�~��ѣwp���]Ԭ.�}��=�]T �$$>�\������*�|>�#��`�x���)��ڱ��ص��BLV�����d]i������Ab��臃��XIM� ��h������3֞�gdM/]�ߗ���С4�vF6������q\V��mU{�'��������I�'��t��3�7�cPZ؉0��N�c��#e�&Dp\]/h����� ��5��:�g~^�%�m�N���'��R cᑟ���m\��A��,����+��Ñ[$��CDi,�ߥ9���x7<�	�`z�+(����_��,ͧY�t��������w��.Pdɲ�lr�NM�$��pwo0��u��{��A�&���Ib�-��AY�-�	�p���v�~�f���Jm|���xE�C�3����g@t'#H����Av�8�At�.�7u����<Q����^T#t�Xms���0��u����u���v����*nv�&:%�raEZ���XX"��=�42��8z]A�rԳ��^��Z�gh�[|�.p��_��֍̒���y��#�!�����.o{�n����S�Jr�1�<8hFl-0'ӻ+%!&�}��e�g���:�$ȩ��ܾbm8Ψ�j�h��r�EE#����=��"���,"&v�� ���O��{=A�R�ib?��_�H��YA�����{�1v;o�G�Ȇ���I��e������f�{y��;�op�f���2���� �B6�^�s�~ّ��7��<e�����)-�	9���W�V�TBT�p�2���M��%�����nu�x��}@hη���>�����rn�}C�2xl�(���P���?t�r���pM�I��a0�	�)�w~���ș�r*��I	�+�RS.��G�%�Ƚ��c����_�x`�X��;��4䮫<mW<�5�[|�h��F:Eѝ������/j��
[��O,w��H	��*%vv��6j�s�S{uC؆�Y�<S�ck��f�y�~�5|���Φ�<��^�3S��>xŮ\�-/���+�Qr6��/\���a����`8vM6�siI�@�k�M:����&�鰥�%?�p������8�[qY��r[�Vg��x��'�U��ʫ����m�;�-6-� OZ9��:D!�
\o�ȢӶF���3�;/��g�J��Cdx^�8J���"WzO�UfP�m^C����[[��(�5����s�d"��G5� %��(��R|���ff�k ��j���<�H�u�xOvw��a4�X(�GT��_@ɛ7C�ẂIo�֩��J{�^g=l2Ev}�Rz��t��)~~T�P���t��]̌	߉�U��"O�W�l�;(�|��WO/(�u5�s���s2�P�V2�7e1�X��1�{�+��%<2��!]<7.���fy�	&���QdG�h����˛�"�����s�\�	�����;`j�N*0�ȃ׸t�^�ڎG�1#�/�=�+�cs!(rS���3����yDY��ڬ�"8&������S�j�Ґ<�;<Lb,�R�cTYZ
D�⇶6+3s���wl�pT�ֳw���q,��IVK V��.�ۻ���18;�?\j-���m�dvfIɩ��$ǈ��rs}HYF(8R��1(w�'*1!b�NW�����<��-!���}�(�FӋ��!����"B�g�H6��1����=�0(�XN9��9GxԐ���nU�Rd�ϩ���J���(,��b	]�CFA�)���� �m�����!"|�J���I?�A��0�	�H4o��-=r��Ŀ5GF���!F&
�"�範w�x�P����Ҿ��\�|>�Pط_�fz�7��5ց��[����%N{�'�u��}�x՘�c�z�S�]0�{��G�TBQ����ɭ>d��t�1̾Ѻ�a��)�@YTdi5�Tڵ��~|"��0ӶL"k��Tǵں:e�$?����O ,����zx,����RBe'�HI��PJv�ΖU��3��
!{e\��I2.�2B�&�����|����qw��q����|�q�gˁ�\s���3ˮ"��ñ�/�w\�WN=4�[�w���R<��'�Ali�-q��4L����3����|6����w@TN���9?��� ܌����y0>dN�����F��&���FZR�j��j�`YV�f��;��F�N#K���f͆ƞ�ж���r|��m��^��_��2X��C��/,�X��z.���=q�k���^��� �voHepӷ��3�x�ȃ�PLg ��Q,�P���Ґ�vp�L,IbO��~qdL,�KS��&�J��}��e�A٣:LE^���9�M Q_����m��
5�?x��="�#d��BYp=�+Z�`4���PUZ���v�A4���!�Ǉ��>��cR�jV�{2ȫz���?�T�K�d󹗭2w��i�m.���z>{���K�P#�=4o���c��?~-`��y▴x��%-���������U�pk׺QP���b\�4�4�̓�At��nq�$�>�͕�f �i��&�`j������!b|@��N��F h!�$�.U^^�`���[C���!k8�l���%'�O��[�΋a�m���m���Ӿ"oem����76���W�F#x�F\=_�����w����t���;w�u&��/���v�K�w[T��e31E���E���j�|.*J���-J_�y��I��T�)5������EZUu�O-id[_�j)�U�3�N|}|�l�o����qV�:55uNSK��er+s
��j:5^w����ъ�H(�;����� ���Z�K���|�P-0=��HNª�ȍu�z���5��G˩Y�þ�ö���>�y��A�UY�����J,L��!R���E�ww)���l�������MK%u�F�!򞨻i�����JDee����ʜ��`�N{[1H�'���������n�5��[��0�ڃ4��Kn���=y�����6��>�	!!�@u�����i�����t/�3o�s�}�8Y��<{�J(�%��Ը�*7Z��[]9���\��~	D199�S��	Q�y���R��v!S��U*�9�
�ZR|�'Z�WV��T5�3Bڅ�b(�op�BCK+��r�P�ZUٝ�D"QRZ���W܈JW�1��rN�QdM�!��pCs�-�"�����$���dX��"TZ����B����������K-��e�@��2U�8�REȗ�j���q�w��ՠx�&�@�Խ���%��W>��^���.��q�W"�����S-ky))uuyEEC//�荏��ے��<uby��+�HZ� ���8�|�SP�0��~94T��f��=�<O��{�m����	Uh��J�G�Q2��)(��3Y�er~%�ć̜�;��"�Y���:F�~��[.N�W~���r�nٶ$d����pF������Y~&|����|>>�s7�̧�q�*.��$	�K0특gm���u9���?M;d(�6�u
0_C��eSE����}6�o7얦L�
�x��iS��
��@SWiJ�����\v��^��sp<�N���U���j�?�P~��ia��+O��-��25�����&�yq�U��\&�B	S<m��^����[6�B(MN*m���]8����F�tӃ�����K2�$��������c�g�$^��*�ѧ� �xmz���̪)���sN����ww�L��]��DDD�5�\WTf�F����cU��p);��$�p@p�����N�y��h!a��ؘ�	��VWC��h�=���h /��.p���1��:���
��^��ӎ�vT����4�?ͥK6ږ4w}�AF(9ٞ#���'���������k<"���J��쑗�ކ��a�ݙ�;�� ������S���l�va����s���_��U�kb��˵M���|��t�+'v=̵-���8�M�\�)���I;'�o��>-�a�J{eZ�����)i�2'��}d%���}����I��Hq�X�ֳw@w�.M��$s�t��Ȋ����QQ��$'add�g&'���O�Mk�f�T���{YR�W�5wF�-@���TqqqāV�7T+�I�_o�y G봺#������$��'�sJ�T��a�F��-P�w#GG|4��>)�Is��^�11~�����1ί2�)\���ʊ�Ҥ��?���V6n:��(7���<dg/�{���'o�%��5�!��Tʻ|Zr�6��앹>�� .	��+���L�}��z���7X<l��8�%%B ]V������~%�lX��C����Ńmg7~�,���kHE_�xꜝ:p�}_�uO�C���$��_"{5��	1����ȷ|o�^ ����"����T����Ez		��R��|�����^��an�]:)�H���l�3r�we�{m�����Q�VB����nq��A��m*���|/{zh�;��j���C4���'^^'pUL*f��nz�9F����Ĭ3ŝЖɦ�=����555� r&%��.�J{��+�Tc3t\�*�ML�,jci��,�c�{�3�\�o��ɮ�q}�fWÌ�����g�e$㘽F�=���va �w+�����ݼ���l�Z�т��?�W'�[��8�WT1�!�Ȱ����`��d�9����nk�׊���C{���OC��`���L��ߐϒI1ʂ���Rk풙�N����v��z�e��zz4�y�苈����~W++�Ț�Kڲ<�	�]��Y$���5
.ęV���*8�3�߱lu�k&?-idH�'Z�ᄺ�5�����;����ыp�"΂��}vj�7�ODw����~���iE�lZ^I�	���3)K��ic'�5mkI.��ܶ=�)�=�g"���v}=���я>�vN��K߀͵4����B#L*,=�B��R&��R���ǋ�~���Y�_��,���[W�h�u^��Cd����0�QX	P�.Jq�?��F�%����t\�����������L`�]f-��T��l4Eh+���)��cS��Nlmo���|	i�P0���܌���Z�C�༕�O���wR��`���X"�e5)f�e�_ߚ�_��M�	)+;Gt�Ѹ�6g���X��pUƫ7������eh�/�dO@Q4�$�U�@`,�0�g�{�Ė�(u��߿V��b�DZq<Ԉ*p��Ar���8E�����Ld���g|��տ�o:L�SR�R�?9mh����y��ѳ4�ŵ
�X��5�����������É���(���I9���c�gY��}�*��*B:�8��\Ƨ���H�F���!i�̺�Rb���P�|`�a9�
��DK�2�簢��%K4%*��A	��L&��hå􋗵T���6��qC�� � ,�L�
��J������+�}|RL�1���R�������� �k&���Ȉ���mP�ᛢ�F�*�h� 	�~G���5<�o�zƓyh*2���+n6%�(�v��Os"�:����{ɼ=���k����&����wn�@�O�E@�����3F�vF~$Qz��Y�C��u���4a0�_>q$E�E��##�^bʿ[�fp��j���uo9�a�����~*yy��<69�V���!�m�\��ː�N�r��)�cp�
�2硺���a�H􋱅�0�b	��3Ǉ�,�c�ojQ�_a���UP`Y�8������$f?}ͣ�ܿo��[�%����%�>3c^k쟻�
$�0a5q���e��.i�N�f�Ezp�B�|��	�]r�O�=:�$?57S2E/C�rq�B{>G�B�����e wIEE@]�a4�rU����kK�m|��DғQ���-��U�B���>�h��K�։�E��P��''f�IO��FB8%дϘ����Al�M8%��v��X�3��׃�������-���*�gs��/��%��5LL���p��p��T$���ߗQYdi2��:4tb�2눣�H=$��MW"0�����i5�X�,��ȶ�:��M�_J
���R櫙6�5#o��K뱄w:���G�������)��኏��yn}�k-ųW��3���W{�Ï6_K� |�����Y4&ni:<�,�"ě�5���j�@9U�g�O�S��S� �ύ��E�����Jd]�G��ѝ���>��k �fg�(�Wf����;�YJ��U���1S�Ǝ�b}��)�����)���]��X�P�;��T��B<���Tʏ��������6q� ��q_�3�'w����"���������6��"o��V�3���O������s���ع��𞖍�9M�<a�������&�"	�-���|��������H3�G2.����-��<�И񆔪�)�����-�m���x���y�mN$�gς:%�e��p�/Ҝ�Rcޫ�b��u:&������¸�ۧ
پ#�b�l��--�	<D6x��.E^(((�Pp�pc}��J���o����L�N~_����e�<�?0���;#�Z7OO�p#F��8'�$>�������M��A-~���uH����{�Pc����.&PE��9�����`ck+�:,���hd�YpQ�A��5p����&#M�������V!e_���YV����r�C		:�p��d���K i�093OS[�y�����B�̵=�Ĝ+�����*~6Zŋ����W�/e��y���)��t¥�qN�j!H�"|��r�DW�E�Eed�t)��4��I�8S$RY�M�-��&��B#�Y���:n�I�����;YP{1��zD+?���%F�9�pڱ�i"�<���@RjT gW�~��c:�{V�%��?�2v�U�+wŘmf��o������n�{,K�WW�<"C��ea�gf]��07/��8��j� p�&p��vYv�B�z�"��ee����f)U��^�8+�}�`}}����`}��S���n�"&Z%�#������rװ��J��݈{M�]�����}9�ސ'��E�7[׏P/Wʞ����9h�d����2uOh���,שHk''Wfe��rM�GGmm/lz��_�=�{�-i�TR�i"At;3e�EEnU����_5�KQ���w�;��_J�zQפ��MO
C,�k�Ȃ<���m��_&+r7<�Yc���^~':8/�M� A�o߹���� ��UfrR���d�$��q�l`��HZv��U�Z�8FO�hp$��u�c0�պ6ض�翋���"�F�̲R|���Fl������!�pr�c�:���5�Wȉ�����*�yuD��_��1GV�tum���j^��X����O�gCv���kR�lF�^<{��(�s� ���������zv��6)�� ;��6p��xa����l�O^JJJ�V��D�a���;���`�y.�������i�Mtܫ��Nf�������)>�vj�܊G=�� )0Αw��UU��&&�ߌTES)T��+!�C�����*-��jT��#�<L�*���)�Hez��� �<å���p�������N�R�g�E6�W�<HrrǟXXk �X*+�f���Rm���R���u/�2��tI��+�=�� �6����|a�&�71�+�!��KM?�����=��xz�u6���'1����tƏ׋�/Ʌn�Fp�.F�������C�D���%%ꁕ�e���ihh^��o�Պ{(|������ERXz&y�W_�"�����������%)�x9��Kr�QPϨ�i�3�扅�Ɋ�����5�ɯ�(��~��$INGNp^H��#&!���}��i6����DF..���g�(��S<'~wZ�����<���7O����4���+,�������T���3�&t@kt��.����1��M�M�N{����7�$δ�J�N�x��85?�.А��SKs�_����"��of��QSS��HX3k!��+$h���4�_o�ޏk<����<�3���<�	�R���!F^^�ف�4*h���m
��:�.�DHJ��%$������?Ń�D �c�^YAe�̵��&�4���r���5�E!Z�m��)�e����n���aLk����Y��[�3��ӧK(=6K�������kP�/����L~R���V�&���-�sr�*�0�k��t��N���(D]o��P&򛚺
z��I	^��r>��I�`3~�C�c0Nը���*��f�+}/�\�
��Y쑻���HAZ�3����j�BӃ3��(X�+<�gi!�z��Ċl�Q���u�ѥa����Su�JO��+J�#��m�r�8��j���� ґ]�Z��R�����������'�x#�]^�+��69>0 �IOjlmݲ%a���(�96&�cn�;M1�,{f++�%'���B���:_K�p^SV�3H/|�u|���xŞ�N��V�y��M���[L�L��Q�y4�EE���s���cb��y�6:�;�����}|��?p0s����X�&�J����=�lj�N�۷�9[�~�
而,���L�0��[�Bݼ>fO�&�<��J�V.���Y>�n��	/�=�r�)s���:�Oc#��oss<з��6Ų�N���fv����kA|��ڨ�ff����­������C��xD���M��jt���8_���P��nz )���?��w�ɓ:'ffhw�OQ"��>������,H��3���'�,P���,�g�cۦ>���=T�rt0�{���,@���iʐPă�\�JII���M���"���E}$�dʧT7��"���b�s��|E��g��D�C�k$n�9���a��S˘&�����)�7٤�Y����{{�)\��o%Ì���R���=ill�����\��6	�C��	�q�rDF2�-(%m��[Ȁb�=ST\�Z~�n��Y�%!a(�Zy�B���R����;	u6z��n��@��X9$�n2�����^�z�(R��3�*mx��(��\��?ҙ�oXm#8c�Z�l*�	Z9���f/�H�B߇���q��ȭ �����L��
B�R �J�L��ՠ2��ui����ћ��<���������z�:��I���٨#-�t�0��{-vB��/�B_�v\��'o�_���O������F�*�P��%�v�N_	D�� *�l���*�O���/����9�5�4Zt��;�{�VR�,��lZ\�`x��x�FQ���s��*�r�O��t\�5)!Ư�(������<�:�p*����Uف��?t(z�[P��.�O�-���R��`�vBa$n���6͸��v���+/͌������[g�Lx	>��y��FA�����k�����rvKNⶕ�������zI�&AV#w�S�����CK�s��H��",/Y�@#�a���ڃ�s�� ,�Z@X0��>Y ���B�)1Y��"V�;���w K%3�Og����w�_��q7�; =H����1�/8�wY��`z�E��|�J�t��8�=����n�11UG��݇ ��=�����~�0߆c��#�m��uL�z\�q�(��"�P� �olj��0��+)+�J%32��T��(����-V�`j�[卋=��4�.5�Ԥ�tC�Vh�TU݀�{#�|�uйL��e��Op���E��B�c�d��^Bn=�*�`@�����g|��'*6m깭�����> 9Mg"�_@%ي�d`��`�F���3�?������IW��Hj=z҂�D�p!K���
D�\."g��j`@��ޗov�f��~�>��T���%��JRg�.�U*��͕K(�?f�9�{b��@z06����M�.��K��O�Ѕ^E·P��A�AZ��4���8w.fe�_e�A�J� 2��Йc�7N]�y�� ���U�<i���nbHP���%��|��C�؊��y�!	�_�F�pM�i�aŭ�w�^(��#�?ۆf�s	$�6�'��A�,��/��-�Q�p�9-(8� #U�e�������oz��=�f��7a�_K_������?QXߐqcm�^M���Io�Z�p/��$��]R�� xV���w����>c�6�AM�5�bi���FE��40��Zx�	).�|0����ܜ:�o�^�_j�=����c������׌�����9
�x�~�
K��{11�̔����g"M���(���Ln�9�Mc�~Kg�<&��Wc����������{)��B����OMx�e-LpuC�8 H�:e}9�|��Y��}� ��!����W��}��P���s�"��+�U�E���
.�K��)����_�6,Z8[����_���U �&��[�5���GVS�o5���/��n���x)���;'g˴C��������o�QxX�e���������,�����b� g^^��	`�I%�~������,�_��sml�d�eO�cض�\n����w!]ݩ.D�~��I�q�:�L4�^��n���H&]^'Z5I�1?R ;���4 ױo��֊�.'Ϭ���G�]���b�{����ͤ[C���n�B>Ͱ��r'�z���G�H0��&+�΢�x���٨_�eC޾=�I�.�磕��]k��|����ܵ���f�-`+߱�X�_++����Ty�M����6ge��lnz0 ���b��Â��=FE!'"��ڤ���<����TŃiPc�,��롕�pʑC�����!3
Z	6��^��Ky���&d�O[G\�s:^{N��a�lY��@�^�"+?Y�*�F�]SF��o��Uy�(�Q�H���o������^M�n�S2,�����w�l�9�n�k���ײ��w�";��ؤ�B���]��5	|Ԋ�G�}���e��.CV!�%�x��#�<���%���b�nP*�d$-;��c�����bg� ��׷�������C������:cp�z�<�����Fl�C������!,*�C�҂�	B;��`��)+�I�_�g<�z�_W58��Ç�k���w��jZ�n氞���<j�����OP�e����E�����h��p��m�$�H��-1~�������n����Ai�r����E��.��ۯ���sd�m���c���������H@^�`�MP���W3�K�:Ս\�S$�S��SPxc��h�
0P�Q�c��;�!òq�ab ���	��h�ar�������>��b�:#)a��p�c����e�,�ۮ�����''��E�(��;&���#�z��:�d%X�
����8�٧�'9ȉ���/Ȟb��]Uf��qQ�SyCHpT���
�Wk�G��u��ō+�!��u�Qnb�/p���#�A{��4���)�������<99��О�(D�-�s,�FR���+�x�����>�A<w�Aĝ]�,+��q&�2(�X�6��-��.^��x���:^43��%ӯ�]��:3C�l\��g��E�[��N�Җ�9;��)�����ÇLADp�mN�e�����%(�y۸cH0,V�h���M[n�բv�a{+��g{���שiii�"r�Oq��_�@���|hll3?�؈���f�����ψ�l9�F��������������/�yT;�t��EE,�����O�-�B^J�Q.> ������gx�3�J�����}����
��.Xw4fiB�bJih=��z�2���h�O���nBa��o4��?�a��Ɏ9�r/�{���/���z�!߀KKE��v��/���ǧ�	�RHT�iƅɃ��wf�Z{��ub]���xO��QZ�Hx���z��m���5���
��vřI��˽σə.R}J�oB�"�O�59����f���x�Y��*�1]�r�HBB��K���*�b}��i��i]e�jӨw�Q�K�^��O#s��w���U�:��yǆFqr���(�G��%��lB����hV'�$j�0!A+<�qUkѬ����嫸���Ĕ�����f����JW��򔒞2,u|||�>}�[���,]N߄�>����d(ѓq�7b��}}=<��95����~���ͽ�Fu�d��ޭ�t{����G_�-<n���̲�?��8�חUe�m:���XUUPX�I�{be$,<���7�3�x7�`�G�2�_�\���B0>
�C���$
%
W|Դ�q|t���VA^���#'�ؿi0��CXD�ҎM����^[�M}�e9mtd���Zr׫�~��[��ܹCKC��{t��UX��ܯ_�Ϟ]4-��&Z|ŀ�$��������@.��4���]�|y�,�ԤG=wk��*>��Ϡc�$--o
���*�^?y��cs����nAX觭�[�����Og��w�ccMk�<g�+��8���XZO�Pf7�F�P�K��4_�i�/ڞF����0��lȷק	��989y�\�$��Z�֭2ڋ�M󲲮Z��pRX�qg���n��[2�������ٳ�j��h5���x�吿677���,�udb����j>�� �7;�Q��N��p��o o�jaaa���IS��6>A�\��H�������HZF⦲_B�:*��N`������)mos�H_��:;����/��1��@����� 2{��˃����.v���I����D����d̠1�Ztt��<�4�	���������)#P�%��
:�J� �BCm.�='�Vx8:�7������ѨD��!n�;KLOkkM���򴆆���\o�e����u_]Aޥ	�0_X��ţ�>S��3M�0��.������P�������z۾V��(��J�O(�D����{�g�x4s�s��b-��g�߳�$zAp��qB����=j{�>�����L��D-��jt��pr��-~�x�r!�38������������Jm�_�n�*�ȘL\�7M�ѯ�(������m�<�e%��0A�fMNR��E�KaW�n���>\���_�H��L�:�B�s(��Pn�Z�I���tQ+��M��柩_�Z�M��t�k����on~aUWi��:kni�*-D"G ʐc�;�ijJ��ۣm�tG����prv9�D8�������?��>EH��V�F��2K���*�f�^ΨsO�wNI�d��J�u��Z|<�;����)hp3�[P���ټ�[衡�	b�=���h�O��iR�^�=�
��	v+mMty�w����ei���g�f����bi����z��oB3`>n�����`�%6�ʍ���@0��d���P>�C�ml���6Qh����v��-�҂�������[)ii7�;f�Gl������_5Sq��m�]�{���%��ޛu�==ʘ�iY�D-	&n�Z넆���?��-��p_������P�[y:
F6L{�*O���sh��`ajǽ�L�v�P>%%E�� �����^����d�~��O+g�����8�郛/�'J0e��݅�?��ƣ;�~7�1�+���}Q�=�C��jt|��k�{�������3с_�<�����͵���'%��[�m3��y�oݔd�ʏh����G*(�ڑ-+s�c��?��t=,��g�:��A�B��ɚ ������^��:�P[��z���Z�v�+;55W�����c&n�LQ�� J��Л���3�$2����Պ�1X,�Ma���W5M˴@���@�6��~*��ө�h�x���D��bʪ�KR�Y���z'��	H��s�M6^����֖��\!{Am|L����������O�蒐�X����_��o���D�gQj�j�� N��M�[�S�c�8�`|��ring��?��ݿ���L5� �53{���M�a���k[_5r|9BQ��E�X9tq񣃃����.Rny��c\�]7�N�Q�gR[�yW�lY�������#P���ng��\���v>�)����+U�f��
Ϟ%d�8�f����޾=0?�����'Կj�LUG�u�������������-�9�c��}$���O��.�v{�!�K��/loG�G�c���
��+�-]\[Z��sPٔ74�ttt0�L���+�ݏ���?^u�hnP�T�,�����B:!�j��R��������
妧�� �]3rMR��|b��[S�a^K�kk�o��&-�������4mu/��SM��u�
e�{�Y�\�A�;�GE"ˬ��VE���Tء�.����< �,a�蛿���7sww>7�����:��|�}t􎶦�0o�ewwwEC��z'B���\�^.I!i��[d�N|��ޞܮWj�7�,Ĩ�9@�����^�6��ֽ��<t[����p�*u���[Y8����_��>7q�"�ry\��1��=F�<���O�b0��yk�g�t����*J��ܤ������>Yl�v�7Gu�����r�1�CV��1˞$���_�W&�3��w�����.]Rzwʧ�����*��Ν�b�s|�Ƿ��L�=9]otO�����?%J;�x4<�ZpY�Ҝ����uGh�ڏ�o��ߛ�
��e���ki�g����8��N�=޹�QZ^���:��~�]/����u��FHHI͝�����@�۾4+��誷����j
G|9�>��t��x�#
�4��d#�9�V���ް;���:�34�xL�6�o``	��U���|�<����f~U�#�Z�̯!chǅ��������݇U��N���e���l�pq�tT 	��j��WA�m.��tu��n~#�l����]����30�|1�N�9��a/`�@�A�g���ٹu���k��;;9��֮��>B�{�vk�t��M���P�S�9�T����eQ�:>O�{ob�UD/�蘒��6�j4+��L����/-+�=3�;h}O8ݛ&0ci�&[�~~nN�w-�	ZYT� ��v]����*D�<K������#�<�JC�mv��ӲoO���z9y���=��oz��-�����mm-}}#�n����R��޿%�Փ�Eu�w\0Ԏ՝b��v�h��f����W�����e,��~�>7��d5�L��8�#p ��D��N��~c��v�����>>`
E`Y��� &��E�UU�vv�C2��H:J��6�+�*�Ch���:�����EE6�</e���h�e��:���������w�3��i_��˙zv�p4�o���v����o~��d��!ꕝ}M+N��륿<�������<@�aw7ak�e�'���X�i.��J�d�'��}��T�Yj�����.k�YC[��z��_<�� ���xl�4��II���ISB�,>z$}���Tέ�'��^Pp
�H�>y9���ޜe�c���]u�dT-*�urO�LOgsrq�(?�/���f����Y"ş߿���p���tvv������x�V��/^������8[.;�![�>Ꚃ���v��"�[.�����\7���̀��uO��2""��-ncG6b���C���,�b��� ½�ի�����F.��B[u�<c�lml�XG����`J�_��I�2�!����݆��[$[��-���w����f�W���[����/���{���D@P���4��~Q]�Ս�'tttFۜ(�|		����uH�FD��9�O�������*��>3��c��oΤ�{�)�q���Tv�KK� m�F��D��2F6�^�g#g��<�=�Q`�*}N0����ښ����z�O�}S��/�VP�od�آd��ַu�{��z�mQ�6�B���Z~2��QM�; X����e?8��zz{u676����M��:��!V�����6 ���?���`�L���W2+�Kl�\l\t[�����`c-��~~Ǩ$�u�A#C�̎W�Y�����nL�j){��&x
���;����E.�mP�k1z�b���4�lԡir�U1cg^�	�l�6s�����������z�uʔ���ط��ֽv�f�I�n߮A�ʋ��z733�?��=�s�{���@
��� ��)����b�HW5g/r|m��t���O����:Eʔ�8���*|W�6HDŞ��������?}q9���&*���C�c}�%�ݷ�&bZ6���s����#����s�0ߜo:wLT����Y�^���2ۘ�2+Pc3�[�)c�}S���l|R�[y>������N�
����m��v����:5࠻���l�N
Ed!k)9�Bv>>E�����ʷ������z�t1������(�!Dun��fB_�w������b�R��ۗ扻���W_�<��N(�յ�?4��=G�V)�M����7'"b��L�3���|*�y{�u�,-E��n-�p��X�������:e����ߝ�FGF�4ٽ�|��^TП�Eu}؊�M���Q���iW�ieH3Z�����Cչ�i�c<�Nnb4??�Az[ |��M~@	� �[������ŧC[3��-χ��G��1::���j�V����nj*k���5�0��11�4GD�]��G��Ć"�Y�%h;��{]}31+����?��������4�i�Bh닻>��nm݋9���ɛ�ϩ�[��f��#�ml��lwhk�\�Q��d��h��Лԡ޻��"oІ�J�{���,������9y{�_����,�l�:��8Hp?��^oqii�1��b`45��@?�S��}�^���	/j��6��p2�����M�+���BU��Y���«S0�;���Hl�1O�Y͵&�Cu�$���
��ؤk����Z�qi;������|h�
7�V
�Ā%@|8ڪ�P`Ѱ�}�ַ�>[�:g��}����ʬuz�6Om����3���K�D���n���N�KIK=}6?d?}svvU���l5�`�I3�>�
�ʚ���/���:,�>�1�t�����B�:�pkfx�=x��iu#�nm���:^��pB�u�0�hbR������sxk��ϝP�B�����υt=S�8�߆�W�WG���Ū������Δ̞|%��J"�T����x���v����.ӭ�QA���[�@ ��c�w_D􍜤��{`��xs?"��k8���\���d�a|�5���s���X��  ��,O�!~��G��M�d=Ī���`S����}�R�m�,Fn�g��x9���SO�)��f>�t��4�ql]�kae����s&�J��0����
Ň7�{�5�7RM���.JK���v?7z%A[Q"b�=�$SU�o��K�?�r�l{���.��H�/���N*���W�F���x?�8#*���8F�&.nl`E�y���뷧��{���Ò��������G�0�-,`�MdJ�i��Qzw�A��aPH�����K�>�/_jI��ha�ﲮf�>���33#�}fB��*��W�÷�o������q�	���;�f�>.��M).���Ǝ�x��0 ����j��a�&�|Mv���>��*��OPK=����c�ӂ~%TV
����G̗��=*�L��Tp�CX���9�ow��O�[��ȚJ�	��z9D]~>pr�����fJL�@&_���1��P�{^�q�(��w_O�J���_�<����&�sa|yj�0�W�Q��a�ٚ����J�?�@�WkiG^r��VXK�ﻶp�h���1��UP��]�S�o<�0l��<�:t,+`S��׍r��Y��`Oԏ��d�6�$�!��sX��iqp5o��Ȑ�]j�v�dis�$`�K�4�t����eͼ�M�qw��侙uo���-bճg��^������p�I"�90H��Ν�tAa ��ը�*�|�IO2�%�ѱ���}0�K�Shl��@?/�����֝e�,F��������{ݍ>:*G��� ����[^4=�P��U���d%z��5��@/TBˠ �����%)L�d��M�lt� =���w�2?�̈&$1VƩRX+,�a��<6E߶{�h�
GG�ӚnN�|�`��`�H�F�(F�����J���o/;9�����a]��7W�#�������JC��W�C��D�����_��%��=f����D�M��>���:F\�r����]� 7�\�v���r���sЫ�;��*�#����y��U�UU���"???�63�lYK˛�c(K�����?|��ԣi扄���=VTU��ؠqw�o��~:�-c��b����6�������!��k+�4�h3�|7�M�C����,����5��l��C���I���J��ɼ�|k�}0�6N%L���i��\����L���P����7���ia���Ðe t�����-�O�(/P�8p�6,�t����[�D)Q}���*��ޤ�3n�>�]]7.E��yg(��ڒ6��uV$�����U:��z��lPx��כ �Q��Հ/���c���O-|�v�4~�݉�a����N�W_��!�ܹ����?v��)�M͂7�Y��1��R�:%�~�S�}˴î-��PK�qW}��B�p��nS:�� �=8���%`yP�{�d�� �vb���X���{Ga���$��d��ՈG2KY����h�Q�ȯ����uQ��؎�0�l�c;L�[>R����=ZM���|�L{�=��յ�����x>���&I���f"�����vgwR��I���曒YV+XVA�Ap�F��SB���G�q�5��z~I���뜺L��À��1G�%000__�3MDOo��-��w{zEEs'>����p,BZ_���3OL{�T3��5%�J��!�����:��E>{y_��`H\G[5�>"Q��h�{��!/�l��w�n��}\�嚱���k8e�Z��Ύ���忥�+�U"���

0��q���zv��(:J#��c?o%"}��[����>�`Et����u=+^�����1_jO��D_O��LF
7~A��}�'��fDDFV��+O;�t͡&�i T�r��LӉ��V�gCv�pՉ3��+�펙u_�^�<��W٭��T�T�J�7qŨ��)_^P�����L����<)׷��M��R�\�������)' ,`�^��&�T�N���B��8�1nK���,ů�Cs!Qp�a�K���Q�6gL 
���VA8��g7}�����Ľ�:�5�bdp��-;*n�ɶ��ib�}o��P�q��|���`����W�*��>2��8�~�E�a�q�+�+�ݣ�_�����7m�w�Y�O����A���I�iy*BuFpxlL��Q{��MV��d䅔�T��Tm8����R&3J-��N���VaD�@WwwEU��2���:{�{��8q˄�~�}� ���G|���^lb%C׬���a=�y��I�++���B$�H������<�g0��R����h���uT�|����FZ��b۷����E�0?V����r�no[$���SH�ˊ�����s6tZ������x�K��>>��='}��

nn7�b�Ġ�����������[
뗉^U���6O�X�cŮP�����Z�_�
�ۜl'��v����7�~�!��:K�I�"�!KsF�7t��..9��=q�G>Պ߿A;]�&u�E�Ҳ�����g�Oy�^���0����zA�t�t�}�����L�?
5��AJZZ�f�%2�� ��j��e�7ݳ��)وL�߆����΄W�=�����8+++�X���`����G+77	d'������)C�?++�����M�,E��~̓�V�.���o`���U��u�^�Q7p���������Q�k浇˾�/e����Xp�	��P *M�M���>��^��[lS�SBO"��	���L��3�O�:aa������:---�	T��~��g�&�9� �'�q�-*Z�y( ��O�o�R-'!%������f��8�c�4����c:>y�A�G�����e�
a"T�!ST��G������A]==s�]S�~p����{{{��" ���2@��;�\`����:vj��ҡ�pq=�ڜ����Bo+?{�c�P���q��9$L.W�Ȝ�g�Y���Wou�������Ւ--��(Ym�e!��,c��F����졲�J�&T���(d�R�&&��3s?��������ݯs���z/׹�G^O���sD���9��E�.�*�O�3\�V��j��Մ���历_�UQ���K���+��V��������ˎ,{���_=��E�/�QTT_YY��Rl�Pﳼ�jv)x?����D1�~�/�W*Y\<���7%����22�~�2����4����'Ѿ
���0�&��9�2�߅���-3M���]z�)�]V{3'�{{꫰��-Y�9��ⶀJ��K�.��R鶰��r�2 T�^��	}���k���� 9>����a�O]ll����A���ꔕy%�����_��[�{���Xp� ,��t�S�2y�-���,��]ua���}�m�����r�b<��B�{��Tx�W�_�q))))��w�}Ꝭ�m`�+W��}9^SS����C�g�����|~{;*+����|����?:%�+vra����T!#&JO��������
H��
�ujW�*]�P��+�Y2�p�.}~^9����73���0�qQ�"��ߔ��|�/E,���'���c���=����A7;�+m�I����"��::��{S��K���k:�(^��+���U��4|��S�@���:�;^7�����p��>qږim�{Ğs�Xj�aƥ����ɫ��I����Kbmdd�Y��`��������hЮ<�oh�������5O������?bt]�,LP����q��k�+�]�2	��rͣ= u�!���ӝ��,i�M������
�v��y�i��޸Z��ձ5�HH��-.$�z�3o	*�E X���.�������Ӄ�怷�#T(�**Y��K��꒢�֙��vZ��� QN�������}��?�޶�6���ގ�Ћw���KAA��ӳ�/��MLL��[���q��2��銊�#C�N���nh��\"��{�fq��1i��;-������͵SE�Q������O�������_^W�"'��[ZjUj�p�MѨ����f��yiiihK�b=$Q��H��
�DM3s�?�72!c���'��2ԗ��@|���OmҸ�066l�5%���f�Bw���e+���5qў|g&= µ5�?XKѡP(��5�o�!�����ymx�p��l$�Ç�FG�8��GG/�$ܸ���V�d�z��ŧ ��b��*�"�Κ;��;Y$r�n�s��#�����z��ŋw��U׉%�u�%z�&|���;32�]3��6�[d��CX#��D$H�۷o���.�+�,����;Z��(P�wv��Z�5���ɯ_� jÂ_�|��5�p�۷m�&Qs�*��<73CJ�=��4�ɨ�S}�߭}!))�� �o�Q�}��1�Sh�o�^�ݽ������Ҿ``o'?�3�a	��?��e��l-v0]���|�Ȧ��@x
N(�!��v�`X������
>![�}=:%���nm}xK��L&������L�=�������	���Nb8����Ƈ���3�Vig��qx������,0�

�CC�0Ň���A����E?C�.�з��|�&s&�����D�=B1��4{��s�LDf9X?:�<�/��h��t��@j�0�,�iei_��終ώ�<���Ó'������M�|��u��09�ap��	Ԣ<��87�����G�\R�UQ]]ޔ�'��hk;�Yk=V��NGG��ԛ�R8�����@�������� �[s�G!�Ү�@F�FrF���!��x��7T���ҩ_� �=L��!z����V��I�^Z2xQPV�>�U8.s�n�ؾ��0�ea��O��+�k��]�|ܺ�r��M�ߥ��Ӱ���w��"�t۸O���M��C�2��
�k���(ͨ:������V��`p�"�_Ł�{�Aw]��vq��}.q��e/�`��,oHw�X�M �f���1v}HU�zWV2�lٲc���	��))�9D�bEE�#5�K}��Ve��Ь_@J���ˬ}n�"-b��vf)R��)5F�W�Ė𻜪�T�t����__Z^���Br�Qi��c�kA�����h��

K>k�R���atj!#�4q��!9ע��J�By,�|�=��x�&
����Ԕ�W��J���J���[��S^GmB���h�]����Ꙓ��{���©���:��~������������쑻��`R�{Ǩ���@��S�ڟ���li���R::n��t`�c�� �Tq����]���&k�Vʘô��ZYY1nsb�h�/�#��`>'k��+"ӿ���o�){[Ў�!<TH�s�����)W\W���n,�ݘW�=�V=H@��S2,��	� �<�L1���AKED�uu�u�����q2)D[V��O/L��t6����EG�J�j����{D�^��KJv�)w�L�0�4j3O޵�*��Y(S�{��;:���ז������6�6�B`��jk�z�vlD}*���#�-
Y�f�=C?@����uk� �\+�L��C4;�U�6`_���65|���!�w
��Q1w8��{(D�b�L�T���[�0LQv�� |�!e��5c6��t�4�5���yy=Q��Hyd�<�߭T^����7���5s��^p��|��D��kW<�:���p��UL��O��~����穽;7�C�D"m�\��J�E����d�ě��~z��L�4�ş�����ǌ�|�߈�SZ��yә ��Tb����@S��]�9�W�Rk��WU/0��4鉠pɕ�G�w�|�j��/��:(0���̚�qg�g��g�m7�a��X�%�5ƵĞ�ޔ�?i��&󨝡Lˏ�y�v�)�@r������5Sy*������<<�?���}�f�/��Z�����ξ.��;�@�?T���n������y
f�/�eW������g�m��K�C�>.++C���С����������ʸ��6%���d�t����P���jo=$�h���=F��X%_��1Q=~&����a�������k�d�`.6U�^d���ݎ�svt<������TESS��ݷX���+`bll���+e<K��ikw@J��\��G�@vddCj�+�Ϡ�g�Ev1�t^�"��j�ݨ.�Շׯ�AG��=MJ�(GT'�����>���s	�		����$n���`�+�3X^^���7\H8^�����,wQ��@�#:W����ݭ�<�;��\^�����ޓYz���J[�K].��B�Đ��/J5�L6i�.7O_����K8���Ŀ>;/"�J-a�A�}�Bz�ϴ����Ctt��W�u����=�A bl��ӂ!�]��@>�U���!A����)������1�}6{LZ:�'�i�a˵Hc/���B@x���g��<�e�W�d�V�}�n����_�E��ߌ�p���FAnL��!?�=1���$:.�#��^�{К[,�}bb�Drr2D<�$�fvv���t��HN��ڝ�||�R2ݻg�� |;6�t��7�fm�XF�쬀�nW������� X�o��c2j^qB=�sq��<Wa����������r��q[*jj�XXtoڙ�^�	G��%�%v�"�������>H�������+���5��MMi�~ yq8��dgg����±b�.jycc!�H|�.�D��{�d]˗P�@
**�4y��s��^f�F����J�v�i�s�U��Ó7Ng.8�SVV�+F`ejzA��%e�0��b�d���-,-�&&�d��/���H���� |,l
{�C����	��wM��?���tO���6E�]��	c����O����V����O$��~k(-z�[÷�e�	�y;��o7uD�[�=b��fV�<�'P�B�Y�Q8��������������ń��/ttt|����.&{��,.���xT�~(�}G��}!�*G�Z;���)*�d7>a��oĕ��E���̻*?��P%G2[� �-ZP1��}t��E�I�A�D�-�Ʌ���#������d�=�aO\�aXX��̔O�^��ȫ���^	����;�NM�*�`�r�n�gd譴&$����)"MAV9Y~�� ��_��"-�����\�<�ڂ�a)hz��)�LFG���SDFN��sDD�ĸ�qEg�V�թ�隁 >}����w��<o<�������z�������6sPt\���$��X�剠=��L��_�jt�>Ä�K�;s�L���d�,lXEʃ���E6��uu����M�#�[�����L }J#^���8�rkhA�ð�N� �z?[�q���

f����5��o�?�:�se�kj�b)O)�I'����$�jӹ����J�[���D-��>)��7�#����t��&?F�ۭ��r�9����W;���q�������,r� �9����skFx��I���/��5,M�
���LO����ֿ�Y������� 9Y٧���)���T [*՛_@@4�!�p��T:rĜڥ�诗�)!?r���VVBo��F uAt v~f���E|�^MZ��3>o2��8	wx�P�腀�]؇^t��$���l��5��8�dť��@||��ܻ�x��w�2����h�����ݳ��J���[�5�z''ol��0K��|t���jˆ���ٌ�ޚ���#;���1�SS��q��ZG�3�**v����nn����̨D:�Y?�ևd����0��\-D��]�#�f��\K����XU%rcC��$.G_Qe��	�_����m}��5^n��E�xo6���G�Ch���z���Գ�M���::;�_<M����7JԬAz�ZAa[jZZ)�D�ڜ;������heȆ�mш�+��C�.��m���fF� �k��'������ͨ��sX�7�5�y���߾��vC���O,�0ͼ��:L��\�q?7�!�H��������6��:��5��J$t��W�ъA���F�r���o�v9�����J$&0n_IU��ř�!�'���LH[�D�XI�|ӦR�Tb�{yUU����jH�e4���*�tJ��qb|�
��WS.n�=59�T���9C+$��� |��a?�`
0 �D$�[u�-�2���P��Ӎ�Oʹ2ܷ�	�korj٥	8�~�bOb�^�����N��j��G��J>�%�����ڇ�w�UgeYC��ޝx:]C{����nU�n,<Y4��'x��llc���,,�@�>!MHެ�����r� ���͑�ԓ����岪�� �@�����n���Z�;I�]td��1��ە��8��i�����埓�Ew���3WH�_?F��)z
�~��������G��
��/xB�u�n̿�w޿m!�W�����)馼/@/���ܕꔚ��A7�+\ve�Z��C$yAډ�cJq;l$��3%*=G73�;��"� �	�jɐ��)�����#��tB�����l��]s?kj�	d� �A�W�N��,`��D�@�E����Vk��p�"���I�7T�WL��?U[��t�����=����'�v=��u�|��>`�9�H+{�z��^G����Js�4Nt�څcF�>�z�x@�3@����h���!y��v�����o ^Ss���QAQq:t�y�y���
��:~nYi.|`&d�E��BC1���J7{{cF7u�8��b�yA$\��G����,�6���Y^F@���<r:���(s	�����5)��,҇������Nn�k����2���V`H!e`�w�И
}7a��1�f�Sp##6VV=�O� ����|��,++nh���c@fQr��T��׮�G��i+�?��{V����i�t]���Jim��ٹ������7�9!~�RߠB6�ÚC��sO>޸��Ѧ���������z�({㶤{k�Xo:�6��7$��ܢ2�A����{O��$��-a9X�BJ��h;R:GwA�0������P3I3�x��rN�;��gf�7]g:A��`r���]J���_2\co�599�d$V�����Oo=_6��p�v�����/I�\޾��ƙo�jPaֳ��M��>pxG���d�\��1;��Х��ߜ�XN��\�066�;l\;XRY�bĹ֪�S���=wA*����W��oE�*3�}����r��4�$50#�o�Ĥ�z�/9 �c^�`Z�	ߙ�zQW�<�����RJII�0E�&���H����V�-z�O��L݀4ٱ6tt�j\����۠rf`�Zh~avP����K�pkg1�D<���~��ZQT���%���gYJ#�ޱ%Ŏ�o�j+rC�.n}��ME6lx���{�S�AV	�]-'�uSN��Oт�F��ԏ�)%d{�6t�a�	v���L%����'��)��C���r㢽�������s�4���KP��2�y��qE8���DF�Ȭ��^���w��?�V@r<P��`�*~c(��N���]�P�Ha���Z��ZG�i���u��l_[	�eb�0�D��c|ㅖ�E����Ś�L�
,�ȹ�Y Ƛ�"����p���q�s�"�g��!��cW���P��d-kC ҿgOk�D���������~~��IZ�Yu,`�v[�,1F������2�6�u�̟Ǖܻ��:��B\�Br��I�G��ϮW:�2�󖽽D8,,�Z�F!���׸n��+�i쁥�-�(Q��� }ĭ�4] �[���z�V�%w�Rː�Z��l\*����kᓱ��g����96�|�%����ŏ6X<�E���l�/�]-+sY��Z>oh�*O[φ���kR������ʪ����=�X32.���+�M��*ͫ�2+ޓΆI�ɤ����L�� Za��W�����f�10�P^�P���s�E�U����ʔ�e~!���a�Ɯ�!���k��9g���̔��5Ct�(��Ҹ ���[Nf��=_��Í�6]Q�"���#UC�huMv%e��(�Q��-���Y�w>*�B����Srs�C͢N^�:�?VfY�g6cX�����=7w����Ϳ��F�
�K���ۂE��rso�������77�k��L��1����L)��]�h��7�C��o�ml�7����O��p���9�fiQb����v�.ګ�`"�h7�}�&�&z����75S��<:�a����>�7[�����|�5Kˍ���Z�m�S>�.2� 5t7ĻU�������\f��K:v�chu\P@�}MC@>���׶��dz�����0�+����+gV	��0�W�mҸC��Nx��]�^�����.��^&�u�Ndۍ��b�8�@t/;*"� B@����i��g�b�=u�w2P�N�Wl�tK�\YQ[���DY'�S�rqp8c�v0 SR��v���&��gx���Rj;=6M��6�`��1#�0�q&j�F�rei4�Ce�C���(����Ak*�̦�Q�_�}��Z��C���6+���bî��%?�h���>+L�ܔO!i��Aw�s T�8��X)���_Dݚ��n��N���3S�!���:�hr�mr^���O2��͘6�,��~�X�y;Gkk5���3V�.Mt����z`�>f`�s���X7)}�^�	�4 =����P��)9T��gJ��U���֞�!�S��t	UCh�e�n*����E&���u���3ƝƋ����E}�a�j
ƶFi�߭�������V�f�Я;7`φ^I������wz�T�o���?�5_<�o��E/G&hΦE���G0�C��ֹ��e`^y�2K��":��q5�����\��:5�n�5�@��1/�wc�rr��_��q6���]+==R���{�ď[n��NMJJN����h�^=��<��2Ǳ������C{��q�}2�m�r-���ʦ���T٫�cHe�m�+w�k�0��#0���7n�)J���3�*���;8�F-"Ħs���r/o����hȭ��.����~N[w<���>a�6��)io��I2*%�C-�#4��w����l��j�@ ���-&{j{޳�[�qnra��bߘ|真��C�J�1�ƛOi!��7���F]\\D�q�W�)us�ҞI��;[��p-z��0�C}�D����IY@�����M疖�����8�2S���r��i��=��8�D }�T�פ U������;ZVV��\��se�:�A`����<�>�M�V$�-������"_*���}B�@Ƭ@�!�vG�$j:ySo�~j��q���ő��+�l��.��HOTe���+ �c�����aG���u�a%��u}����믕�S��B�DE7��I�'��.]
�pJ��A��r��$v��W�SqII�t~����/3@�[8�S |��0\�M��*|�n�J�cY���.�`�ii� �_^~�Xp�ā�5V]�ڰj����uto}�|y��[TjG��TZmm�>��U	,��ELh"aLV.�@29aD~�bX�`�b �]�6��e�:��P��y��ϕ0�@�ܜ��񮾚�ӻ�m�ҧ��{񌾝g76 �p�ڥ.s���;�ZfV�a����lR^^�����b��d�9C0��kj.��RK�K=��i�ZQ�����WKU�.��E��/$��LT��/��~"+�B��Z@/�8��[�JKKKM}K��㓟�^5���9�^�m���O����v���U��S폱G��ۻ��sF]S���4�4ݹ�.�Q(F2Zt��Op�%)�Xi��kf[й�v�E	�@�Rף�����ܫ�Y�C�=�u�N�1�
�K�4�AG.4-'�!�zN�88��?�dK�~Jȇ\\�Q�o��`���3>|�&n�����s"CxLsi�Do���`��E'ｉ�}�d;���|����	���J;�'�!*QG�l��������Հ���Fy�S;�uܧm� Ϙ�u�4��= R&��{�%�WF����&)ɫ������e韸��S�v��U���ң��. ��<��3p�x��5] �\�|�6��D�iiy�؅�mQ��wv��u�$��qT�K��A�q�%���?��y���08G�(SwZ믤����!@|���b1T�;?P3N��K��9��1��S܊C�xMmu�����
��q,J�5J��6��Ӛ��q��;q7�hGSN�r��&\��'���4��^&1ݵظ�v�y67#��r&�{�P�m����ڔ7u�u����l1Ցv�����C�.������1~�/�:$�*<�FY��d��k����g�v���>|���,V��<G���7�5& i�j��8�-�}��ݘ�Bc_����iŝ,������ݗT�}�0$����^<�Z�x �8Chp�0(Ez�9�,�h+�ZLzH,�fo���Z���;WVyP�����v`��#���R ��VK6]���w�0��u.�q���� 	oC`�{�f�$!������<���twOO"D��l'Q���c,��!��`[a�9�.���:�1ݘy�dB����&$���RrM7G\>�-��]�g���}��f�����x^�S�X�*���=lڷ�������d���ʚ�/$`BL� ��>��J��,1+>_av��l��זa�'S�?9 "�q�\�`�fk�A�z�Y��,/
�1��q��;�����UU/�	
���h<��4����6W�A�'|��]�D��`�7R�b��&h����x�L[n���g���j���]}�"�����*@7�����>���4��:�Jd7��n������
ћkl�젛z�Tk���i!۶�����K���;�x�U
��M�$����7.%��(J�C\�i�Fu�����c��%���܍nd�d��-���d�[�G�Ú�HOc�Ʉ1�R�>��jm�ҴB�	���Xp"�ԧ�Wt��r��Ҧ�A�����E=�E����9�d��������r|���$/���ri\0iH��{;��o������C4��<�Ǹ(gf�\����2��w��V�Q��
khr�6n� @J���k`���r'AX�@��I�9?�O�YZz)R|�w���Gx)Xt�'������(�$��E^�%"���[�U��9��[t+��F33c�:U�[潉}���ht϶5o�M�clB��4��_Z���}����kB�oO���O�-|�p�����y��l�{���}��@�6_�5rP�w"�5���99cl:֛���~Ϙo^�.o�T|�}J}R9-����g�R��G�:yԨ3M�XE^���s*��ey���l��s�M�=P�2(�/f�8H��ĭ�%��	0^� ����:���;��ew��˩����&��5�8h\��6#W������VC����La%�kgJn�+}hb��D���C332�<�'�~i�)��c�*e��(��=��X�^p�m��q�۱���5�� H+���>
W��V�O�������N&��}m�0|������4d��n`C�1����Ae.���q�2s:=�$ȭ�o�B�3�!r��3�w�A�,-R��Mpe��=�o�9���3ss���'�85ni�a
l�2��K�d��h�({[t����Ύ���E�@���^W�1�5������
�Y�by��rG;W��+$= �ܢ�XƩ��y�YX�x��죀zL&��U��͗_p����?�щ󀇰��q�\��<���������sv_h�t��>���,lP�q�D�S��8$���+���N��>x�;��A�AW{�]s��e����T���d��J�ߡ9��:�q�
�v|�����ƻ�A��S����6��Yw�:�ͦ���^  ڊ
|q�����׏291q�Ҏ����637'uJΊ�L}����F��ٿG�CW;� ��
�gE��P�V(���Wң���v@���	fffIN��كt!PV&���y{�-����2��`�
�3!��4z���!t%�r쟋IŶ2�5m�k˵�3�d~Y����yW�h������ҟ�h��F�sC3o�V��d4��5=�\�%Zsgٙ6���<O7|^��$�\�\F�(�d������d��Ø��O���~�T���}�f����Fx�};�����nP�D�@�M!v��s���/�kγ.��q�;��E�!��4��4�.�(���w9��'�Pҝ����#�s��<�:PL\�H,�A��L�o!��)ߺ�X��1����'g$�6�����M�g�%�wSb�'�~�V��o��
�u8�����lsj}�����G&�=��<A��-7G��`�ڗg(l^��.� .yqCa+}�y��q{�ν��ۿ-3$t�������A݌ǀ �V�;�K�ݭ~P�#��b~����w��_��,/��qQ�b�M2������<Ig^�Zp�`��lN2KZ�n�[�¤wf][��9��ZO��x�B=Qx�����q'��΀�hH���	P�Y����(�����Z-K������������;�*w%��TZ��m�u]�P��-�R��4�����i�����չc�k�ux~|]z�p�9p��۰����II���~y�����x#�5�e�v��qp#' �ε�*��`=<,\ȿu�2h�L'^���<um�^⋧� z���;b(�\��Xb(���?������S~�oqG�kٟ���:�+�˕�h�4��t�!�gȜ:�JYWCײ7�c��!t����D�8��uj���N�� �v���n�7�H�*;�U�0�� )ɮu�t�8	�_eG�bz%���S����㲣�N��|�B�b5e�ŏ�0���r�; jb����n��ә��Fe��
DY+6�ymϜ��	9���f�q`sD�I�u��AjzzO*�ȏG�`?~�����h���,J\P�Q4ں?�b;��&k	 kq��e�Ly,�Er���_	\��2)s�o2�����������_K�#�9�#�K���p���S���j$�<�y�:|�*���9KP��� �h���vU��׮ᓚkC�Q�?���J t������1�W.r]�^i�!B��oD$�ġC�\��Ls�T�n��U�e���� ��fN��E�V^�j�D��~�5V���&�����oZM4c����+A��>��)*Y����Ό&��0�X�V# A��|w�3�%@��Ж37��Iڂ�3o�֞�����y��Y�k�-�ί�P}rle�3O5|	����u���9끭,J� 8}}u���9G��(4.��!Ϥe�(7����?���J��Z��芠����:{����0�A`7�؉��B�Vu���H�Ufe��հ\��24s�;�xv�j�������o�)M�� \��]e.D�Y���,�Nf�iiğ?on����s:;��Ԕ�+�ڿ��x��������]��S�//�s���rϟ]�$��ӕ�����rU���	�4�ي�G��--��X��be����z�w�����o�fΧc�J��@�x /�$v:R�
�-l^��Ҡ{�b"v�!3�����o�����mm=��$6lW-YU*�Lh��ts�� �5`(�8㤩9��Z���@�}��� 
�Ʒ�A��!���wa�-�4�WwG�����]��g�7�Vڟgi�����!������!3C�!�ˡM]sb�^;�o17f�m���(�5Ue��V����V�n.�v@޼>�!}U�J�[Tw����G�Ywh�����4GF$yB�V����C9�aa� ���X�ΑN�^k���F��+�L+]��-���<���T��F�.�h ��|��>ey��1�ԑ#;���5U�3-K��cϵHߒރ��A���Y�'���++-�H�C���3M�C��ۏ̪�qO�����
a����m�7^݁Ef"SYE�y�B�O��i��ο/�X��5�?��c�wÚ�-58�Z�B��E�t��`Q�
�vʗ���N��fo�\{����ǆb�! $���D1��,�.r@a��A��d�|�zUI�[�Z����^����1���[�{�K�5�������]���A0=����f�W��J�3�I��ip�-�]�.���d�RZ�R��j���FQ��k���u��ČP��T%K����z��\�DS�h�-�ٛk1??w��Ѵۊ�>��AyT*���M����S�����<5N��e6�y�w��ø��'OF�+�^��b?
�K�I9}}�I���=��/H�w���a�Af�"A���JlWzcB�1�D5�|�0m���(c�gc��
�]��.̟�����Sc�ĳJ���F�)tE��5����|m_�z�k�.Ձ�#{.�zVVZ}����2)Z�M:��؆�'��|)/��[sdRY���9H�U�h��uX��\�B�(�s֫=r^�@�Hs���0����_��α5퍤->��/4��){���s��c���x��C��Z�#4����Z��'��)�*��sd4�]� M �ǋ��X?"��'5p��.�������.�[$퇒ILw��X��U���Z�\�\W���0^�J�_<"�D�fr3ƾ,�̢�����]����� �{ᅬjӣ������������11)~�)���v[d�S@��|�pXj,������V�6��Ufwth��C�N���N�����U98(#���a���6^6t%��c�&
��$wvv�&/�i��>8��ЛkJ��&{�f  ���n������Ǭ�h�����ކF��Y	�Rf0e5�^���J=�����Hk�ng\r������my�M�'����B_"���B���J�⇗/Q�i�p�Z,�FC����Ds� M�U�C��0��$�������VW?��R7��W����Ӄ����M;c� �%��i�5�m��ݞ������p������a����Ԇ�����@�y#~<n;��񀌡��b�R?���M��I��8ŸS�l�J�cP�]ӓ��(k����[ɹ���^�@}�~��L�<2��.�%v[��ac�+���s�ݺm��D]G�J7��ס��C�bMJ��^�2�	��������5�e�����d\�y���(=?$"�g�9Y9��TD����}<_���W��r�J3I�j�ݭ��A�'''W��i��{�T�UMi��*G�`��n�����4�Y������ik�	��._

���u@�������m��\~NMi�����d��<q��tq�f��A�jN��n�uJ�z����� ��O�����7N
Ƞ�Zs�x�~;WsI��yq�����>�)��r���������v%	�ր*	\����M���֞�Y�Q==��"}	��r�'3���J�nd�4}�jC��q��0<�f"�D�A���m\��rǿD��� 99vv2)g�H�rg�$�Ҷ>ał�`q��z�P�Y?�+(tO:-�⣭�&مď�y3I��d#�D�c-�^)������l+Ã��}�ωce��vn����]�o�����t�����n]T!��Ҹh�9��kg�~��6~V M~���N�[<���c�0�����h��e�����(u3�(��������������([�ͨfT���Ie�[������R�m���l����!��n �ԅZ��*�F��!��\ߢ�������g�a.E@CӤ�>S��xJ��Q��nk�5�"��]z*��QQ�wƶ���V����?ɸ�q�6��u��[�P��8} Q<��Hգyx�;������j7F�Fe�#G� H�
�v�~"���J���Ξ��
�>�����f\5N�;�0�Q��V��W�{�A���Y�BY}�\��ˢ�����g�y�W�ä$c�NP��Dp���[�0�̏��ԋ%��"�
�7`��ϲa՛Z�Qsr2
9��p��P�A���;(�9�h7��[���~�n�Z�1�]���^av�_P���X��/�6T��.4srw�\�;B�3'�3@���y`��- U{z���ڭ�뎁PI�y�)����\P��c��3��RJ��J�g�^$!�D�ؓ�iugD>~���dT$*Ǥ�+�5���=���b<�qnrtTz�Fߺo-6cg�����10A�R�U\"5 �k
>�/���p�����$�M��\{�p�am����P!���/�xoo�}̷T���
�5`$�L����7��C�w�2D�ls��)��Vq#�!!�>
���_jY�{/K�ڙ*6΅	߰z���<�j��61x�Z�㌧֍�ي�Sb��޾��V��d�TԄ���֩M�b�������\��h�.|uǺ�L�κ}u&{�y�����[Ǵ�`C'��PG��c2���2Vӟ��$�ס��}�P��lǙ�q�u�E�c�zn2V����ܱc���IvʁMB�E=>>>�
���:.��q#�a�gM�=֪=�����o�B&t0]Gj��^��0��*�U������/0������!�lSB0D���$�!�
�	��CV/K�U>��r��ZL�st�Io�Q���C��ds@DE���N4���|D�1�5��߆��`���
5۴�<�����k�M-A��Q��A��a��:%E�֮;� Fǹ#�z_<�TrZ�w����e#�>�����l�㲓���7Q(j�zg;����(��7��C�X�	���1�����Nv#�n���7�rF���^��"مn��h��B!�r)�\?���������\�Ʒ[�^C���m]7L�,�Gd������� x����8v�C�9\�k�����	����ǐ�Z����9�碷v��q�l�֣u� �y��Um3�)��b 0��-U�U�4�G���p��ZV�@$�H��� f��Oy�|[�X؃�.=��}�m:������.0{l�.�˥������c���d�36�:�1�-]R���b�Je�`�z܌�`k6��7N�)��^�э�������Oh��� i�:c�Z5: �k�4N[�)�W`0*"c��L��˗*\�4ow`�k�)+�����s���}zB��I����	w�y��|^N��7R��o��,k� ��U�tqq�a2	�Vh\�p������}������m�D|}����R��.^�0��n.nn���v��u��i?S^�8�G<����w�R'�_`:s��a~~����?`eE�<��UD�"�" ��OP|�����69vv͉.�aQ:�蛘\���F�ȃ�2K�S�����%jLd������C�0���s�r&�@f[:+`�w�f�=��;7��9m(��|Tʨ8c�W�x�~.�4�s�[� 7�~���>���?|Bt*.�8�U��' ���/7�
�㕠��7J̋�ኚ��A80̥�	�:�②,��4�[Xs��<3�~7���>W��B� ͝;�t��88-����+�p\�e#�g�B��Aki�F��㘃=s�7�QbQ	i������Dͱ�y�[ֳ�8�At���KF�K�Ҳ�=r$[���M���~��k<�F��1*q�2��c�n��ݳ uԙ�[��w�:�`g�I[Gg�'��%X�(�O��W�i���M-ޝ� �Xt�W��K�����WP]܄�c@x �#qפ<�����]W�p�Q���cF!@���5�.| @"Q�T.ϘY].-��X�'�,q���1�5�T�]�anF�;��_�f��Q�Qz&)�w&n����&��kzl��[�8��w෕3M������3���06�ç��f�K�b�B�B���P|�N���Rƅ��۝
`��v������ �=�	��:��j|c��߃.,^e�OP|����Y�&��M�S�!�.��H�B� ��>sB�ݎ�(m�?}c�%D�M��B/?K�5�}B�(2+΅�;�|j`�~x�qqٝ���u��!�f@��e�/���þp�;@�g0�-���4��/�[\�#4��x)�XѨ�؀�~�|�q)bz���ʹJ~����Sx�u�-ҟ�Y0]u��KK��\{y!Hbb茰����Ў̡�!�I��n(���#���B����'��`�:J�ŚW��}�0���9���#Gv�%��s�?A	/<$������qvsS��&�r��o�f`�T=�L�?s��0�1x�b��~�Z`%�������hJ�K)��v��5]����u?��(@��.?�,ݽ���!P,�Δ\Ђ�7��@'2��SÇz
����	T�� �~�����[�\��k��'���X,�?Q�"Y�L8�7 �p���Vp�LD3��f��>9<�9�;��4W��#�L)�Qƕ��1�j��-�k���4s��#���L�2�����֌"*c#
�q#�$X�Qy��q�0;
��55�M\�,��q�����M��L�������;{5�D1����ʨ�	���H$�!�TNO��X�2�����oYZ`YJ��E�k���qS,Q�x�tB��=...�bX�vZ�)�%	Bo-hƑ��ҫ]^t�gU��k��\�/���A���HT��\��\qu�Z���a>�J��I�.p牡X�ҕ�ݔ��o9�RYyq�ѷ�k�H@�_&A�+H�$�eV
-,r�;�"�i0Op����� .�����s,K� :�f;�E�<��II�PNٕ��I��WĆc!@kڒ}.��=^�8��y<�x��Q]�\�E��dŏ>[�/n$_�;���b���K�z��z���Gd=d�_3�&�
�eR�>�@������`�ް'��?���B�Ƭ�2�X�����ፆ>ˌ�����յj��u��kԧ�

�¨4��q��	��^���p$�r��<���~�J�!���r��IT�ރ���OF;�ŸЌ�b�*������Nˤ��d.I+��c���U/��f�3�2s	�ڨ�Ь���"�8ϛ����{��@~M�֩+r`� 3BQjFR�Ad+�0����2��`�?R�=�-���V� "X,777:����GT�7�x���h�,�p�ϕ|�quA/K�P�.�Ԣ���QQ:�_���K�&]�|��n�W����=X���$�1�ƘC��Ы�F�p�y�� �.��E��9fm����B����yfI�b�U0,Z$�=_OT,S�10�,�p} �_=gUE48�Mx�~�Pnn6\V_<ѫ3����P�v�p���G�C��!!F��S8�@/�CȰ��-�NT��zL���1�`fON���$������XA��_8d������u	���y��f�9�]#S��v���_e�!ͼ���0��N�8u y��w�j��CѸ��r>�D|�E%&�}zFy&]A��Ȳt���K�ܸ�`x��K_��2p�jlKKH�s7��ǻ���^9[���cm(└�aP:��C��E�.��Z[�����������j�����&�P�o��t:'�ꤨ,�RT
5!kG!Ր4��![�]�%ˉP�J��,�ݠ��11֡���`01��~����_�N�>��<�}_�u]�������ۗ�((8�δw,4=�.��=��$�\|y{g�e����a�O���0c{�%�x�,F�Ըs$��E���R�l��W�Q����r��������O-��|�����zi��\�ḟϟZ�{A�˵J�.���ik������s���@E�n@gS�t�`t�@!X� ����Ǜ�C�y��⪗[�)�feC�-S�j܏홥.}=5�D�rd�:�͛����_7�;R�)���%u��Ⱦ�~����pW����R�"�<sl�`{:�M�����WV<O7 r+�vt;�̨p�|r{AW���V~��SSץe���־P=>,���ޞ�5<-���-OR](�f6-���۷����	�R_�1{�X��7��_nJ5^�>�Ӯ���J��<�3�+������<#�evzl7��@W�69�G���70p:F������e����Z��h�����1����rr�룭ee'�O���SPg�ٯ��

f����������w��XwQWA����|�FK�6�%=���B�F9�Q���{�[�,#�Y]�o@ա ��=~���D�/>���V�����]R"�����$�v�;,~�|�Xh��3t���6��i�'A�fG�g�K������sↂ٪<I�%QI��Q���V<�����Cm�4�\t�� �[��i���R�tH MW�WB���5�C�j��.|ln֌m�.r���8jh$^����ء���ľ}�RS>����S�G�e�L&�������)
�*X�'��w��f��)Hצ���j�������4N�c9�[��xI�!4���b��,L;��u�ķ+�/�?z�YN�۳����pp���VffG�u�Msc[�t1GG��%e=�����a�U�p�&�m�̭Z��õȘP)�:���9))	��?�,[����(�R-���fJ7.q�r��9ʸ��vv����m���1�����^[���Zt}�����pެ
eؚl+(�SW_�~8[�O~�������v�e������Z�~[qu��އ����K3�ns��?�u��b(���Ņ1���hsf雛��,f�v0����g!�j�"�k���###���ή�.��t����IMYy�C�_}s�����a:���	K������ݾ��a�_�md�#ި��Yd�Ht���8��_9���Y�y4m�T�~�&��J��x����(����w�;$�������=���[B�ޟ6����騘��`��zT}��61.�W�CrHV8q.׽��ͷ�\���=�`�-i��9X�dޢ2�A�|!��(A�R���Ɓ��Wx5p���npf�N�pi�:1��?�z��4�[;<�YO���E��Ix��xD`���S�p��kGr��|�2|�x�Kk��77��n�*���5����NjN��P�/�	�<�4&������u_�^��.6��w�[YXD���wvG75e߽���K��^S`ЕV��a_�����z�����l���@ʰ���6-]*<�@�-�y����� �>�6��|�H�R��iK˘��8��	(�2���٬�q5�[�'--���"s*��|���e�Q���[;?_�����G�~�C����P�Z��yʱOK?'c�Ύ�e��4�طhƔ��o���R��Pz�c�$��Q�W�� bup�a���2�C�5Y�)r.���崲��
boedd<c�=�5���7�v�Z�А:&,�Mv,���~HRrr����Ǐ���-NmF���h�[�Q�=���r����Cb`���!�)���4��@�q������RY�
�M�n�%8h�n|�eB��sϘ\�����p�.�f|2�tjV������m/Y)�>��g_������cr���K��_O^{�89��oK3�M��܌��6�t{����T�E�����X��|in8�l-�"k������D�zW�3���
7�#!w�،gg�ڶm۬���{u%kQ���R��y�����Z	�?�lYDӂZ��Eg��H�����^����|]6�hhd��=��T��\_U��Ko�Z[�����w��e֣tg�,��|ƹ4�|�e۞"�����ߠ�V�雖�qȉM� �0�:�N$PW8 ��h�L,��ޕ�{�Ïa��:0�f�!R���Ac���Xܥ�
ڭqNDЇE�gV��F�@�ViQ�W	���0���t5.tuN?�JN��@�XC��Y���^׎��2,]������V3�����d��'IrǏo70�� ���[M�R8�����l��ƺ<L�-�WU��P��)��			��+6s��D�IL�%����;�E�=(&��N���>���dCqS/s�����J�?c��sP����֣T:;������������hY���Ϫ����0���Z1ˢ"##o@�y�єS�{rt˖-��L�SU�]^��8���XUmWvJ$q�Hsw��w����2,�Ѕ3�_�t�a�yF�7��7pc�r}���l�zuXfff�
D{zzt���_8�X\�rNw����Q�|=S�z�� �d�d)>R���5���֜V�����k�S���ựE�J�<��*O`��cTaٳ�P�x%�V<�9?�s�+�[B��P��c�j��$�ÞL�8����2:5�B�l��V��k��Uה:KO��?dv�����`�[	^���E��;37�M|���g��[��p/Ǡ�6�������+պ_��2�s�#��e�G@�rG��a�.�AQz�;�A�,c�˩��=J�o[���=Z�һ�t�@�inn��X�RQ^��0s�<�Pl.-���
�D��ϗ��G^^�ܒ�B�
��7|�S.Ek����ˢ����������I&�)�^��aw�SL�Qi	)��C�Wܥ������j.�	��#��
��a�{��ֲ�5n�w���=5���^ӟr�'ME�\�"8}AJ�Q��=E�gr.Ͼ���7�{Esz�L�˾�	�~�1��|���|�C�A�N���ȗ���zs7O\7fT��MO_f�A��sK�烊�V�����Oɖ<Z>H)��TMQ�H�25L���p�L�� ������ĪP�+~s�`ƫ+�g^vwuE�R�lk��R*�� ��B��w*A�����$�5���.�>��� �v��s���e9i)K�`�ҍR�08k�2�������-�3����TmV)+�B/0�, �Ɖ� ����rn��l�0�Eƪ�I&��!���/��N}?�O�9�L���V�4���)a�2*T��*�Lf�����C>��kв���]̡Ξ�)�㣇ɉħ�q�'M�iqd��xƩ��L�j�Rǧy�������.?��fm�*�F�W��p�,�~Y��,#�J]_�\nt4��֒rPjh]�2��΢l&���1xi�f%�(h��w�GHY�T�>�x����2x�\ӂ�2f����n�5���ӟ�j�/.yr���T"IoY%��T��\lU���k�rD�a�N瞺Ky[����Њ����2G�S��p��[@V���cJ�-�B�-{K܃����"�A��}�`��՗`�"������9��p����|�����ԪR߾��O��b~wѽ2�g�ީϕ�+�y��uW�*rN���jf���ܣf��@7�|h�2�:�m��Յ�*��Xڂ�k���,��#�RO�H<��*�k���9_:F�O�3��)�s*����=kI���*(آ���أx�����W	A�QI>�����L��osCc�즞=ل���3�VG�7��I#�=��;�TD�2���!ђv�����XC����/�L�s �a����\���(����s�jn�w������@b��`]$sr���I�#���6�/<�COZ��X��z�������e��B[�;�@�2G�=K�2�[��K�SaÚ� �~J%���a�c�lq���C���ma) w��5���<��p(3�e����=v@k�"�Ƈ����82$Z�h��	m��e���-[Z�1��L]�H$Yؿ[�(����˟kn2����j\�A�����c���LA�F��m/���'��Ř]����D��s�'m4���z7X3���a���[AnچZNY󷵎�C���y��Է3_
������-b^�=YM����y�:{�!_��b���ӜRN�mW\Y������f`8G���2g�e���=	0����9%�)�O��LHS�T.����fw�ݐ����m����q��-� �GOY�,�ฟ��HV_6�b��N撓���e�Db���@�<v?�����{��i @>"1H�XD���qֱ�̭������C�f���e�\)0�K2���_�4$�I�W�xE��ѹ�)�֛B�ۘ �M�����nT3�͸�����2�K��?����-G4��b�`�SNqUK*w)�v�dh�ق�T���6��C�u����*`#X�DhEn��E5��O���aҞ9kP�Tql���bs!V�v��L��f_�	ij�0�|��d�j����* ��N�����6u� Z�^�U
�ۜ�rg��ԡ�%�'�	�8�Gų�����&���.` K����H.���TR*9�[p��MLMá3�b��R�u��@���$~��N֧�ݽ��a��o;��]4s ����zCS���qw���<���v��_N3c%@_뾸�,�OD��b��<d�%|�Z�):T�v�p��<�߼\��B��>7����j�CP��{��� "q��Gԡ�������O�×b ��_G��Hj禞h<r�b��5W��7jj�3)� YasT�n'���[ ��T�$�7�H�J�`o)[N����2(=:�C��T �o�t�|�_vhµ�m��r�zL�_�It�����2YdL���kC\#&�l��9�lOm�*L����^ ��dr��@�6��nr�I]�a#��TJ�\̣���M�l���kn��v��}�O`?�n4�.Z�C�|�i���+���>th��� =���[���mFSa��m��b�ZEg\������"�*���� �F*�ڷo�$�t���ڛ|��7�d��������<"'7ݩvwQS9/��i�&H���7o>CH3�K笡s�|���Oc�\��ي�x�߈�n��SZ^�G��On;�I$��B�e��{`�}u@��+k����֣z�ia���-_�0�����D��8Gr0,�e�,NB�ի仱�z�1�:�?:::PrZ�*�҇o���;xh5 �Q,)K�c��y$�K��y��α����H �|���;i��=�֎8�<�u�\�>~7��r�:@a��Ī�Lt)<�+�x���~� -<E��� �R������byH�f�}��Y�|�C��I�xQ��Y�J���4�+�,i$����S
K���S�W��oa�⊣�j(�&#騸=���O+�6z�2�wbJJ$�!Ã�:`�� �H`۾�-����хpD	����1+�4�M�N���2O����u��g�`v!�.��).��ۚ,�>�>�`��򱱱�|7�V�$#K Gndr$Q���s7��b�r��x��i]*�Je7]I��E�x�w�I}�Wz�r:15�#)�M]�������13wF��p`=Г��3�i�R2J�1S�¿�Bר����3���B�u����y�o�P5'L⫂"��m���]�,��@]���0����چQȭ��m&�v���!U�!I�f��`%1ϛ�� �E,�wמ�c��WeK7�\{:vba��v �yq;{ج���?�li��c9�u'� ��7B�c�I=���Y�dO��������z��\s���I�Oʻ��?Z�K��(74����k��T�Qn>�}�Br�aXL6C�����|
&�3��s��;3��u�}2P���q":=��v�Q^V��KKK}���,g�H~>�Wu}b{�v�Um
zڷ�	= ���~łf�녮}ŉ�Q�[;L����Id�ʞ&�9?rNe��ɮ��zG ત$�)8�F.�K��R�LAO����3��h�ݦ���#ebH`�����"����8z��K��:���z�G{V&a��	XCG���3ؑ��Z�.�.�4˱�è+��0��M��������v..j���ٓ/K�MU�}S5�[1_���+�W�#����%K�C;OD֘�#���m��0P��]���!��a�D�m��;�`�ı^8�T�¼,B�}=��T䕖����S;�r����

_����\�F�x�� �Db��-�h��ύ�&�/�{*��O'w��+�Qp�+��ܽkT'�!t6�57߆a�?�n�	zMM����)+<��s%��zx���{�0d�=���Ѹ�M�!QM:�+H�Z�����H�=B�l�ɧ���C1��Q3��*�>;Zjll�C��~��JA3�$�U�B�E��o�儭�#Z����x>_��aAg��+��5�<��c###K��T6�
iа�U�b���#����_}���s�OvO��)���>����)��Q��xC����B�PŹ��ԎLIS ���y�>���i��D	�P��/����t���Z�2b u.�mx+���Yl��ɰ����9��C�o{��.��
I��j��kj���<�Z�WQx2%\,�cm��h́���Ka]�jʽ��� 6}A���0�O�ݠ���UZ��[�B��=ox����vQd���� �W"P��h3�9@�%=�T�#����0C>���Ta�|�d��^j�M}�r���Y�9�899a��Ә��F�1�X
��`�,��,08j�e���PV*n	E�5;kh^��� ��U"�j�权�i�f�!;�)����d!TH_P3���<o[D ��r�-�F�FTH6泲��f�� �~�x�)d9h���9i���M-նe�ݓ�0c�9%�C[�b��~z<�9�3$��G����+��J�*��{XB����"<�hg����7��p�֜��yR�2"�,�� �u� |�`��y����j���g$�%LF�����3��T�RUZBf�U���l@^�����?�^2w���$tK]������T��5�������(Rهr��S���f��$�J|s�^�jtv '
º�x=�I���"�Vh���|~llj:�t[���X,�6=V�Óo8)�^8zKN��s�$u*��1�xE�:$�G}�A�nBЏy�ׯ_o6ʵ�ʗ����#������̊1��caX�"K���̈�4���n�=vl�}Kjtfff�A�I֞bW���X4��c�[#r7 \C�V\�,A��XZ�,��Lj��
Z덠��ĭ��{���8:2���y�b&�8�r��_ϣ�t�� C��ya��Q����6|�y�Z��h�ژ�J�j�E�@X!Ơ�<&�~��VӜ|*Vc����V�^� �Q�YN�·cV&O^�P��~�s���IY4�?[؊��h_��v|�'ߍ�,:-�m�oIݐ8ӴY?:�20 ���fC�7��ֆo��+e�`��ڮ'+y)M����T�
����/n�S�x�x��	u�s�E7��+�o�)sH���!�����9tfu~�C�����$x�fc����jV|�ba��M���5����I7��9�4�� s:I���C�S�rH�N�ޖ��o߾��"K}E�\^�>Q$t�v��f���b�(�~-���;]}A+e���0��KE��*r�:��y/�]}J���R�2��6k(����������L���R���v������dȰ���w��[�l��z���R�.E��)���o6,���a9,��7��B$@���S�uN�eW�5Fqq[Щ��W����� #�\�<����^��ȅ_�Nf�*�z&����8j߬�ډO�*Bf )}c���˧T���`�4����XaKٱe�"���J�����8�R���oR������;�p�	��)�mԕ�L|͗����M��������n�p1���-F��s�[w=���([x�5�O'F">>~�s&��B�2���5��F����GPS��AW|��C�&[�Ғ��1�� ��QdmAA:�U35��4�`�Mi�v!�`�m�t:=̙����B�oN�W���A6��5P2��W��7��ʨ�8�J)	�7��qO48I�?T�6�Ec�hcc����G4��XDh�UB'�h+�3��ERw%FW�?# :p��e��
l���VM��;dGd���i\���"�����BM�!��<�ui�4�s5���H茀'p3���j@;��$�_44��y<L���cͻ�I�<ͫ��]zْ� �D:ج��n���P�����<#�V�L��y�V���q��?ʓ��v���]Ͳ x;x��bL:O�4�=��Q��crr�3tS�n߮E��$h�Tx�q��?���ؒ(>�	�HRH/o2�c~��@v�T�4oA���H\'���^	��!�]H����CbKx��4x�si� �N� & ���W��6� Fwz�����ox!�&F�!�BO;�8��: mU��7Qh=Fʖ��H&#�����P�Ԍt������1�W���V�$���|��s(YX���ί"cf*��5t/h7:x���E䅈�16�.#�S���A-̙^J�>���Lf9%�=Üa袣��>�45Q*�(:�g/QW��0q _��M(P[`�1�����
7�hr'�Zy1ncq�}���N�u�OCCZ@�� '9����^�ɕR�Ţ���5��+S�'�ƁS-�4��ҭ�b��9���IJ�7_Ns ��_����.�Bi׉e̡�)֪���f�y�&���^�L�@(�̃�e#[��P�fr��	��"y b�k�f�_��eY����嘬��
�Z�4N%�������M�����m��vq�CZ�7z�,��I ԠS��Lt�-f'qH�*�ů%ڕ��~���UC;��G;�z���9�rj@�rf_8�= �f�G���A�Xc�<𨁽��ކɛ�/l֋��ފ�f�?��&gp�ig+�\9P:1hah�5;�=��a�#"kdFŇ<u6���J���&S�SBvb����/�XRv$%�,��ma����5@O��������\4̥��Kۙ�T3h��9]]o��E!o�d�-���"J�W����8����s��nʽǏK0�@#/��S(mIc��)�=M�7<��;��M���>��mz��P��?JI�RZ=�����h�H�N%7~=e���J]�UR��ۮ�V|Sq�3�T -C]�_s/��`�����o~K��ޮ�d��F�2y��b�*_ϛ@TNp��T|g���t��>0�a��ѶPK4F����O�@�%P˩�u��ϼ�Yӳ��~j��fP�~#h�5O)�A�T���n����i��}�YUt\\,��S��U-6D^���Q�8�9l�'�zQ�����h��0����l�/�a���|��R!�E:w�k�I�$���p���K��ߨ�	^�[����"�^t�O��nQ�:�B�A�!��+A:��)�Q�a��&;Í}���%��Qp�����&�B��;w_Z�0p#�7h���1���[$P?zb�$�X��k��5��e�sO�˥�2�`wQ_;O0������GS(�a<�t=ЍX�ޖ�b��c`e�)
<2�c�s�}�����Хu���o�ai�2Yq3��n�T�k���x_9��ߑ��]�Yn
� ܔtceF��w�=���M�͵��HZ��1�_��"]�V��KA��"P��,�^u����T����p.�*��$�S��St߽O2���K(�| ����u�@�I�����r�ѫS���HA�V��~zQ���C�Gmm�������^}�x-�8'��\�A{���z��۠�pG^���K�7�>|�l|����q�X�k�pE���*7w��5��&���d)�7�P�P��*�P1�M|����Fݘ��XR��j�z��9x�L��H�m�͈��sH�E�֠�"?5A.�r���̲�O^����04����c�S=E�x/p�D"t��vO���)�^�x��?��!څ�����wM$) K�q���ec&�����!��E^5;�����ҫ����?�t��B�o�������]�x�)2%��/64 ���3e|�	���A�����z1ϛ�GC�����##.=��G�����/b\{y�,?�`�\�,ggϰ���@����՗24׶��~K�s3���c�-��Ik�=XU����JMЬ3�B뻌���8��P�v�-w��<��]	�Ç)�Og�^8$�.�t�-�Q(*.��G��-����L�R�(NC���Z{{}9=I�����A;v�D����������s�J�/_�~�����h�J8��)?� ���������@��X'�W{������]��H]��`*�`�w;g���ƌ�/꿬����I��m�蔾������ݻ���-BL-p������X;5u�իW�����6u��F�Tȁ��pHe���
��D�B4��j�p����P�H瞲��ȪJ7���%��_�-/-�$�3E��"�* ̹��\geŶ�2S	t;���`l��7Ͻs�s�:Q5�q��-@��K��X�bYK���9vnmoo m?+˹�9�K�ڍ��bK�� V��s2V!1yD&�c�>�k]�N��5�x���ɬX�R^1�Z�F�������Zu�Q:3�	���^�~��T�nW!ڐ
�\���'�G6˹	��+�Zs3jg~�����[����+�͘܅�n<g61�6ta	��$����ccو�����.SB�p�!����:�ؐG ����h�L�S�W�����ܻwr+�30қ�lش3g��Q�o��H���B�~�7��hȏ@g��gdr�uO����h�kE�Q�+&t/���##�%~l�a�-X��e�*��6 ϰi3�Νhra�N����Wхc�>%wz�3�{�-�D`��jM�A�D��!�=�GBSD�%ٻI
�5��#����U�%��ڧ�*��]��#� I��� �%��Ӽ֧�A&i������Wβ���Y�>6�8�T�wuإ�s��?�l����>�D���ߛ�9��׎<a�Q��M�_����p;����۽��?;�(⢏�,ge�rTC�d�2�� ��*��꛷�p���sO/{~?���?"|��X4z3�ہ�
����m>3����?_�ϊ�yV��ܝ
.W����ꔃ)���:K���!e��Ȱ�Txw��^8̏ѹ�H�� &�<��c��D�B��I�J����Q@@��H)w�������X�EC��Œow��P��!�RjJ98[�n�Δ���П;�a���s�8~�:]��f�I�"�8�NH��ҝvr���BX^���� ֣����
�C�������j�E�tg~�G;ٞ62㐸$�������6H�v#]�82�)#�5Ac����Չꛎ���zE#���`4�"��(�`~��{I3��L�����~�ey.�{������-��7�m�\rڄ<).�G{Z�M�t#�k2�O�������eLUnWK�R]i�����MU�$ü��v��BS�ΝIݝ�S�᷿ߕstu�SpQ	&s2�]�^��s]z2�x�9sje�A��=���Mr�M�IB��M������
�.|�r�K}`+�S	=c��b^{�\����>|J�8tW$�GsP���Fv��z؍�]>�6�ٱ�ŧy1p�S3���K\�'.	�L��+GZ�ǣ�omTA���@�u+4͆�k�?�4Ìv	Y��j�/6 %���-#��|���J�}��V#l��R"����wd��[�{z�tzΔJ�b���
��{+H���c�9������^'�\��ܾ��QϤ,7�aC�]2w�N�';��/>B�Z�E�h_�N�w`Wa��NN+R��������E�'~ExSY���D8�� ���V���3�6ю�I)\�2��UA��?i{����	�m���6�^`��o��In�n��Qx���uQ�:��D����F�k��Đ�נ媓(tSe�'P���t��y/3��ր&@�(�;�_>��/�rrr"֗|��رa�����W�̋��{�tKWBRR�c�O���{n���9����V��PwO�U��;7�;�r^me�����ߏk�/�<��`����$�#|x�tc�u|<g���N��d�MJ�AȞ�	@-GN�����)� �pa�2t�_�^��"��'�,C��r�c��r���P���1UN)����u�^���\]�b?��("��]�hq4�B1���V��)�|V/p1��7�qP��Ι(~/��3��G��&�!frYJ5gn
d�;�6$��#�--U&$G�T���ff�f��K�B�EEF�U�l��~Kkt^�z��"��a�ֳ�i��Җ�4c%�Y.|���3ߧ(����Q�/}2��F;��:�\��
7z)��q�v]���?f���ţm���q��X\?������t��'�Vm��5l79�R��e���M��|z�&z��)��+����>S3/�1�Y�?&��R����gc�����,/X'ly�����f�#`yϮ[v�&��Fi��X�f@>B=��u;"��I�CP�I&s'0*��Qo�:ۙ����:2���^B��@*\��q���O�+���pn�F�W��
q�_��閗���**&f�U��Q����z�ZJ39�K�Ts�\`N�xȹ����b'���I�����LL�@ЪƓ�����2~���H���ZVU�BȎ3x��Hj���p���<C}3�X�E���ˢ��<cI+�K��D��6������i�;���ߚH�Q��ke�u����O8
*xX���	��cޅEEOu3�D�[G@նB3���޾�i�0�6d���
��+UyP�@u�D����'K"�N�O���U�i��	.7@IE�V����O�f�|��Q������!c.��5�1h�Es����$1v���Hl�e${�F�Yvq곲,T��d^*��vU)=镏�o�N�%�V	L�d2��# ��W����Q�τ� �i�>~�W:�����3�1�Q"�2W}���h.��Q:����ë?�%KiM��u/[����-[�Eƞ+�"E0�*W����B%��3Ϯ�KoIN���g(��t����?x���t�N\H$�m�Y8�Zdg5��q�\�^6=�_����XwL�C%Oǜ�s�rsp�Y�b?�8d	=QZx0���)���j8��/�~q�Ι���͢p���(�#k����W�*�Pt��v)��0>��Z�^�r,Bn��=(��=�_Rx����&��_1q
Ӊ	��T7Z��aip*q�t$���rv�0�砂}>�lX�����?.Y-.�H����z�'�B�	���Urhׯ��i�t�A�l�`Gw�?�꯶��I���V��'C*~я�Ȩ����?�qk�>�c���ۓ���l�5�D����������H�j���-��S�5�Y|�|�)�1�/�ʸ���o$���!��l�J�Y�_��M:WEW3���58yV4�X�q��������@4��3`O�`�׀P������� �
:12�-��5�:ѕ����)K]�;�k��!7_�ۤ-��k�˗uLx��U��u�^�;��ļ���d�)9v�=~�0�i��/_2퍝��M���g#x��(��4tc��f�u�F񈴽mD�v�gm�[Q��}��7���`�s�5(�LG89�?5��U��N������acɢ��k�[2]�i��PU�|G؆2"k?�,s\\��/���j)�Y��B���9����P�#U8����G���J7h���#��1 1�n�Ю�H%�Ĥ���!���ѡ7�dj�<p��J�Z;�s�qo��tb���i��_Me�/���e�ݔ�D��������+�h�Q"��T�i"I�IY^��_Ey�:3`��xD���T`NpU�ڑ9�[���̘虱�)T"�#a��k}�[b%�2<���{���`hVX��?|	��-�kO�&S�{�;S���~Vԍ�QMh�BT�̠8�X�g�G7��vVcmFj,i8 L�3p�	{�x~fpvq/n�ߤ�Z�z@HH��K�{���#3� ͏��k�{N�bA��S:mxbq�An1ɻ��)�αTV�.}�xU�*�l;��^�{�	�Z�ݱ�H�|䖛Q��Z��*���;��y�LJ�a|p�X�cEs��L�i�9�Q�֓�>�֚�}F�wtgH�[�!&ּ:s[�s+�_A����n�O	����Pȭ�d�����~��ʅ�OG�;�L��A�ڙ�`���_j|o^T\|Q�6�a��W�H���o�2����ATO!��5rg�)1�/?L��ib���z��k-�9��Kh>�	��&��Q��w���P��#���Yo���W�������RVl����Vh�X-�4���q�+ב��A��N/g-�mpz�5>]9r�>�F��i�M6PSxI����a��y��DED~�E2�s�a��Nc=�~�		<RWٲR3R%>���d���\�MD+ʾ�u2��$j暛�knް+x�%?Y�!1�����6;�q��c���w�T�gDl"
:��9KNMg�+4p.B<ƑiM���ͥ2w��UL��?Q8t#�_����*����6���!�����U�u����z�Դ�y�pAI��ݝb1s��Y{#W�4*�	�zjiXƏ�� l���)��e��az�˯��*8;��$m}XA�0�����*2)�!-�$.eF��q���L-|���wo�h�Y���%��A����&��\�]��í���t>1_���_^�ˍLL�������Pfo���/!&ځ&���D�����(1*��f���ڕЂK�x�U��G��3�q��o�	Pu02�ӗ�B���G����DFOs3s,,342�h���\�P�q;v{t��ه�j����]~HNh�+������^��G��`0��E��G*)��绰8�k�j�o����vI������qP�'�����䐩&D�e���37��By�L��@��ԙB�B{ky�����]��0�"qkB��[/3X�]�-T1����m�**���?�)B�m�l ⫟Q@no'�:��y^���rv�(Y���"���h�o���05�r<A|$ݨ�T����4������2���Y�mA�\z{��D�Aߏ��d���ޮ}����R��n�7U@C��� p��Z<��GF[5'3���k9@���L�R��Wa�������5g�N�����u�۪�6��gƚ�
FNW�&C��|[||l�V���L�np�G.y�V*�d _��Hx�g[ak�p:C��UNь�;!��/vrқ�_ p��8��`%T=�{u.xI�7�͕�͠CSf�V(�*�
�I��;��@~5)�V��ΌWg�Ţ�;"�;6�1�P}����P�3�o�}�^6I�1 �,��p�T�m�޼��Ј��� ψ���͔s{+9
u?Pl��L��8k��&.D���z3Q�w�3���j�3��N���64�scn�������j�Uq@v�U"c.-n�FX����+���}k}$�+�q`�\]�ſ��q��)ux�dT���}�D&�x*��+�w��^"{�����"���$�y1���)�e��|,�5C��l� ��_�{Ї==Y��x[ۈՇ)���z��|���#0F��٨6<P�ۗa��J�-`6�ҭc$BbH�YC�9��VV��o�wc�x,�,������O�9N�G.��m�꜇��G�ޫ|��� ~�� ��]�~�����7���k��������Ti�s�b�E��	��g�����H|h��IM��j��+��#�mޠ^���&��sb��+V��$"�R�uw}�O��X��+wwu�{��+��ۥ�H�~��.�]ۏZ���99�ҍ��s'�t�:�XR�|Bn�H�?(�f{{�����aJ4X��\�m�Y����Y�T�򾧟�֔j@�
é�Y�u®ً�ń������Qr~�����	n��Dl8s
�ܔ�EF���X%�f$����͹W�ޣu �촥Д �r,�P��!���^SKsprhs���9�JV�	���E��/�w��|��o�>�����	ݼ��§͋W�8�$��k>���!�]DJkw����z�a�۫�˦�M>h�?B$��6S8�	�TyV��G	��ߗ*�����J��o�`�zD�5��@���zb(�+φ=�}������G][�T�{�uM��N�@!{�F�׍a��99�����z_�^�g�rή���qx��K;ِ?z��emܥ�yU`hha$891�;�7T������"u�b�Sл4��mV��@/�%tE�[��]Z;B(��^�����_Gw�Ә��������e<��.U?ې[�靀2�ҳ��$m��,��p�o@��q\g,�U�q����l��,�e�]���ЃR���ǯ��?8c�$�Tq�_yU|6b��K���4"&�S<d��s']��9I��{a�mxA��u(��t�3�IVu�Wb�/Mm8c �dw6���/[��A�o�\����1i8$vZ	���T�r�[��j�,h�|Y!ˏ��Mꄡŷ(�N��L6�J��/�T���s*G�Q;@0 @Kj��o%��x@�Yz�	�����}-lu�]b�Ui�[��Gaq�w�H����љ�%�lH8ʶ�OrPJ�p��x	�6�|�:�4��8�!��zkڧJIq�:�r��'TT�q����f�a0��ݏ��8۫{u�lv�2��i/Oz,=�������T���Ф{|�%�z� �j���nVk�cն_��~&�ދ����l��W�[ �)���4�1��V��6��Y��)�k�r���3��-"��|R_����aa~,�7)�	�Ώ��m�I��#��v��I.p�ĉ�]�S@��kmZ!��?g��ӹ���^F��,����]��uRJ*&��(?K/i\�3H�#��M�u�_�EK�ZG�p�HÞ��Ƭ�Lf��s���B8��_x�NH(lSpo��0���o��be�!������Ew��֛fi�O><�\�J(�㶷�z��.��+��8�!Cdu�.��&��ۮ�G%�=�m>6+}4�B��.��R{�C��
�:�$G�/8�dw���&���~a��^���]���\�ȝ�j[�7��Y�O\��@�/f?���lk��m��}�3y1m4�SH�X�Ԡ�ڮ ����MQ�����+.��3��:�A�I�[�W��>�󭤆~���3T]G��Y/\��]�w��^s:����iOq��Ch���^���w��O�4�S:��x�k�~l�?�
T�'4
�>�|�Y��7-�!��q��\�8ipN����Us�m�c&��ܺ ccc�!!zt�;S��na6��-N�7���3(�U��>g�jao��1>�����r!�fuɟ..�U^=�k�/�s����|���G\6�?����W��ЇuC�#R��G|�-	��S.�/�*��Sl,\���1\�d���"&O��>�F>����[�5���ĕ������==���$�;�4�7}K�k�^�P�NP�)�b���$~�n�͐C��}Ƞnۓ��o m��|��jϭ��#k��gf��XK�г���|稤5Xy���'��kg��6�9�E|��*�#�:}�(5���U�YG��W3��+��nޚ�˝�!p���1z��
#��jj" a���S�f$O�̩����$�Z��&B?ޖL�>��6�Ρ1��<��k>�J���E�2h�p�@�1��� ��'���mU.�e�Y�A��ۛ*���J7��$@m���DCcm��>K[]\�q-��p)� Mv��B#�0VCY��j���S�Q��5�lIrv�H�K7�ןݾ�G*'�-~㙣H���\���z�:>�f�Gn,*[-�����z�K�YR�j>U���y0��t̷+Lp���?6o��ٮ�uUQ�܎���MiG�!�1u��ſ%��Vt|�x/��6��ݕ[��,XGE<李EO�E����/���_T�S�'[��������?��b��j��i����꼫]���WK��,�z�tds�O���ѥ%J�y��lՐ��9�I�<�R<��\WG/�8�z������Yͥ��&�EUà]��^'F�����T4��6i`�@�y��NO��w��.�{dš��>���&/�����"
�����o^�cX���;���&6����\IA��q�O}�%�CW��<��O�i�-��t���͐���2��B����;����7��VPGA��ڈ`T�`1"��A�����Ju�t+̈!��!E�AJ$JҤ�B��|?����u��de�˓g�g��>{�s��O�r8C]]ʮ�bRB�깡��ῒxju}	Q�y�v��b8f�������g�����Bj'�'`�ď�4*o�J�z�Y� ��k>����\���w�i�VVT�}m�_�Կ��������N���H���zK��dݘq�?������̄=~^���O&R�@Җ�	�Z���4��5*�m?d��`!�)��<xw����A�Zn9�Wk�rKl\N��ݵ�%s��T�U� �ݒ7O�'�x�Q(R��!~	��6[q��R���~������ ��q��m@�F%b�C��"�>y�x�n�ҫ�tl2��ϙ�� FN���i���,~T��U��e������ߞz����Q�8��E|Ɖ:x8�" �h��:�I4����X�UV?���b��ҡ��X����g�r�������g�M�i"6��6�a��7�G�S>�>Žc�P�w�ι��r�+�/���pE�����C�����+��8شc%�Ĥ�Aȋ��f�M ��S�+_��^�2���KQˇ�"�yp�j��Ɍ�d�({E�ZˇF���-)��C�r~Or���]v��
�+l���FVq�&��\�/�8R�;�Ԍ�p��rB�"�=�_�խ�)KWX���B�N寅t���W ��Rp~�5�(~v�ο�4�X/~�Yu1qI�'�F2��$cd@��)Z�^0h'_e��ysGҖ+�ޢWazf���q�����++��F_,N��#In8�&��}O7H��J��#��=*�ͯ����Љ�2d�������$��~��NP�DR�k/9y������[,&���$+9�K�d�xV���aYWU���7?vA���։��|�`������m��Q�J��(�%�n���Uv�Ck�i���1u��Q&�w��>�(�Y�ē=22��,�y��zE����@�az�
ӗ֌_*�N�#/+��1����=A�?�������)�F�  }�yW`5�����7c����ٸ)�p����X���������ū����7 8���,�����7ъVnٹimSp��*Bȍ��۱�G��J�g�d4w�f��f���(ﴃ��"��@ 9{[���8y��f�/v��tCQG��B���j�Ҋi�	�:�
M��ϰ�q�ħ.�Q��,��e�{��
�J��u?�L{`��-(��*�1)��ҧ\��$+�� �J��Z�5Oe�*5 �)��p�
�.�8{҈�!X�J���8��b�%���P(^��?/�]h!EC���H�UͿ��T���]�@�d����t��?��7�8��BFX�z��)����m\r��� �dL���I0w7����A�HUA�eV4u^-���!��`�Bk� ����U:6.�m ��K B�d�mB���,&�-��A�9^��;���o�1?6����
k��:��_Y(It�!K�&��@�p���d��uÃф��Θ!e��H�	�G��ς�ZQsk�����%�C��N�˻�:$ѳ����
��w��F� �� @�F�R�<N�cF������Q}�,
<��w�@�$��SE��
H�F̃n?����ߚ7�0lp���c���-	��f��,�R���/A>״��������6�����0-�M
<���]��T<L��e}��s��4����俗�� ���a0굍q����u�e����)�+��/�� ��R� �+^��U�����ߥ��
��}_���(`8��e�`� A��t{�P�����f���!"�d$�z��#P�]EV��%�9H�EUz�pӁI3h4Ȓ�f�$jf􏏏?�J�A�b�Q�F�9�uG�\��.��"��H~�։# E���ws,�-����u���w~�	,�����1���l�-埥�}si�-�m�������0�-���A�h�%�P���h��;Y��#5�֣,��\��	`!��~��G!E_>K��O:� ��ew�nGW<�'"�t��Hdu�D�p2o ��F����]�.�� >(I2(��dl��j��Au�wVՈ^�Q�m ��������ʎ�:CZ�,�ͥ���\w�3����� ����9�@/�ZrabtDjU;���8G �{��$¼�4�;w$Q��0�K�oP{>!�!k������	���Q�M_o%Q�뭴�n�+nuY�@���-���Af�VEE�n� �TE"(,N����J��f�UR��;|e��!��bEÚܵ&�$�e���D�~4 ��dF��`��&jNd��1MT�6��:�!g�e�M�Z�f䡽ԅ�~��Wf�s�%KV�^��]��ݘ���+��9�_����ƹ�Y[�;Eod�d�-��e���q!=�	��ȷ���:/|�l����Q�`���D�MV����3��W�#�fe��D�g��S�h�`�N<F26}�yz����G)��dD��[9I�U}��%%%`є�H>�#`߆�VF �2x��൲ׯC�Z���yvDYE��"b���Z1��y3*��]T��n�Jj���qR����ZW��*�b�˪u��M��s�ٷ��6P��F���WA�Zn��1�7+Q��G�Y|���B��iI���Ew8�G<�.>T||n��g�?�>������J���y����H�Y?�˺��i:q5��k5�#ȆF�ז���}_������9�\�!!�0�k����Ю�HO6���g+{خ��F[���猪�#�������{�u��K��������QUo0�A�R��ؑݻw{��@t[��N���s��3�֡��w��2��2Լ\u����p\RtY��[W��F�M� ���nj1�ܔ��w�Fg�v�Ai�~�֚�#��h�)pzF��D��Y�t{�+��k/�j$}�%(Iw�[�~&qX�{�Jl:`�]IlW�ߞ�����@��̈�.?ᅗ��<&�#������>9ɮ!6	K���pT�)@�Ź)�����@��޺×���ȵ9���d�-�qj>ӄ�ϐ̬A ZK�����g��@��?��O�#N��3��neHt����}�K���׏B���$P<ӧ�{����,Ev�m�3a_�}���z��v���98{�w+���Ht���Zc��F�S��P�(@��0jT?Y��x�$M�����I)8��0�H�آ��Z���ĥ��>�X�Q~���ē U|�<��:��G�O����>A�������}�A�}���5��3�^��-�w�<]�bʜ��RZ/+�I���=�/�jż�V�*z$�v�G9��f@Q/]E�!�_9T�:1�[��=�U�g���-�3�M���ǟ�Aj}��G�����>$���?��,e,�L�� s)����$yb$��Z۴'�������"�J+�,w/�lb˩4h<�����4�3?�����A`�Q� ���*���9�\|"����\ 	!����Q�ɸ%op�M�>�X�]�ԛ)ZZ>���6�V�ҩ��[;��1��	�gAY`�h)���ڥ&0�ϣTY����܊
ڲ���]�O?׳�cIgh��s��>�vfa��,��c��yg��"I8��>['��T�~��T�.
�T��8�I��͇e�E��u z�Y��ݐ�ġ�m���|'�
�kbd�A�tz���$X;���_��@�:���;���ӸUrx���"2�:��O>���# y]��{�
�f��\�}DMf|�&~���z,`���u9�����<j:!�5��K���9 �X$�����⑕���?������}�|z�j���\ZÈ�6�$H���g�P�qv���'^N�K�~"A��(�ϑke.;|�����C�#�������d�Ê�! ��.�����~�W�]�d��	:{�[Q_��Z���b��+U�Ϟ.6��.c�
Q��7ܬ�>r�jއ��ˉL}�g��,�7�p��*�ɀ#�[8�xH��}IFyon��M޴+�zk廍w���ξ���_�,J�BK %���섾�`�q���lɆS��YXu^�I�kL��'vd_e�1���GC��Qr&��@���o���̓�a��$&P��L���0���LNN������}V��5c����/��ڋ%�2��6���G��Րj�.x�G�c/�ս�8��0��_��8"񘌚�x��k��6QD�z�qR�����Ꚛ���oQ+�a�:[��40��6��a�>�u}i�}��`�(�\q+1I}8 #��j�NuA^��ێ���݇�?�]w�Դ���֧����Iޟ۸�d;$�2�%?n��Ã�@����;�ۻ�W�f\8�&���k�&T�1@�j�D��c���k�$�O�8�'������	C �H]#���ߍċP���D&��� [gk��m�ȈNa!ǝ�T+����h���^�٢�F���\)_�zw��:O � �jx���<�niI��OL\Zٟk#g��:E@��Ja*$�s���H��2'@�	m�-����%�Di�c.DV�y��L��f,²���X�f2��0����K�Ǐ���2�������ك�+/�?Ǧ�3��*�-H�1�,�-X�(oB��1���0v����u���`��j����kpDxxڅ�Ja��N�W��|.^�s�U��ԙ�I��dm�Z`[�����ط��U��"ӻ���']UrU�ML8��n��7ͧ�����]0��?�V�WGf��g��͝�ԒY�ل�!�����b ��D��L�K���!�n~�C�}�8�l�8�gΎ#d��ޅ# M()+�����˫}���r*nu��p�U ��z��g��Y�Y����Ӌ�)bEe�":�
uk�=$�=�Hd3~��W� ��4��P��GN�ED�NW��7�ǩ�U<	�������#���u�;�Gq�j���l8�^��n���4a�7�;�~k9I���F�h6u�pp�i]��u�y�39lƄ{�H���nؗ��"���ܟ����`�1D~��G��#q�HksI�}]��3PAX�C�ѡ굆4�ӟ1.�)�W���<�i��NN职:�*M�����3��+��.ɍ�9�w/<���S��6�U��"�����u@;}�	/�������	p&��{����]���2���[��G����bP�G���2�{[�����/3����?��ӃhSki�ㅬ�[��ܼ���>�Wk���V�?D:V�u��s���ݸ�� �V��5.�a�q�j����'�p*NL�dG`�9��0D�s#�u׌k��^�_l��Pd��UL�ƛ33a��ᣥ���3���{{��Ig��&/�zEi��]�7k����"�1õl�f7{��O#r<T�rz��ʕ�����0�z*ֶ�*�'�-BM���u�q}�����ټ�0�@�-)�LV|�a����	L�X�s����oe����4[��s����Aov�S#M{b��c����v)���:��0̞y��[\wM�$�5!\���<�QK�b *�2�%�3f��¶�f�z������bj`]�%�E�\$�n�����#�R��n1��� Ѯ���mq��9#��z �<R���V�a"�\�;_�ߔ�-	!]�j��!��ԫ�}���{��'L5��?�1���Ev��VF^8�^�2��+�\a�	C7�ٗl�cT��\Yk���6?B	�2cц|nf��["�
�u�!�c����c��M�%h���OR0����2�hJn���]sA*�﮹QT9����J�.�rF����o��B�7�n��VDTe��Yԕ�]3	\���	+���CSʠS�����g�p�Z`�k.�&�c&����>��D�s�R�ʹ�U���\x�!|J�Yr���{��"�s]3T[��{W��G��;Iv�n�-�Z0���BVe,�ZA�g��K儚��!L��U��'���l"U�Q�`�$7 /k��m��:\�Q�a\_	c��[�2��,���
��{~sl'	�NĪ|�n�$��"R���R�YفT96y�1��L��c\�O^�f`�a�{t'Zź���w�W=�B�������0"Ùb��W)����NDF:�&�Y9�{j&�8���:��j3i��O��g�h�W��:��R�Y-��T�e�
�j�Y_�5yY6�z�j�����<����h�F��Gp�uj�pMÏ�����ܑ�D�� ��hka�B�l&��b��]L����V���Ϥ`+3{G��]��-{yxhTd
Er����"\\�[��b�z&x�Ӏ��%� �d����׌���6�������P,o��Bp�7����n�ָͤ=i����X�Ǽ��1~(zt�(�SƈL��B��:��6��[�g#Xmq���DI�T��Iʈ^%�Y�}l�cH
 �񳙰�����g;�J�L�-�^"�����Ԏ]ų�=�T\G��wAQe��!O!8�
�S`��������ͷO(W�M0��Rnogg�p��t 6�'$�8w�=6� M 8�ʁ:j�ʪ44����(]F������Ʊy8�q��f�<I�-jD�&Q����俟4iT�|��~���������X*�D��W���N=&�T8��čj����Ij��$�I.�\&�Lr��2�e��$��/�.�C N�f��_&�Lr��2�e��WI
ٍ�N���;�qC�Fn���7��8�j*´��ҏ���T�?�~���������#���	.\&�Lp���gs�%S?�V!���I��<��Ҏ��Do�C�?�]r�r���'�k�Z��&�~4F�+��ѫ=��:��BM�L��4ū�P����$�0�Q��7K�:أ�-��#y����/>_�����rI�:�����j��Uc���e��UI�?U,����;�(��Q�=���÷셛=��D#,l�|a~��� PK   AaX�34�� �� /   images/4ae31398-47d6-4d15-8d33-5c428753ae4a.pngT�4\m��=��D��5��.��Q�����w��� Z�=��D�-���{������]�d%fɜ���{���]�LR�..!PT�Հ@����	6&��3k4#��U�4�|��� Q����4�n��՜�oUM?./�%��� �SV6��-�5���kȌ��v7Ys�L��6�`�3��+��LJ��#���u�V����e��w�eN��Z�c���fH��1/��I̋{�b^A�Q�|�-�e�|P��Jƫ��"3H���qC�կ�U��yUĘ^����Ոy�IA�\NP�9��R;k��t��~���?Y������`��@��\(Dh�]�H��].�1y��DAHHˀm�P�Qz�������{���UF�?fo옛k:$��Z}�SaD�������o�,S5����}za���;���Ң?����Sxx�3뉢���yߍLǋ�sMa]�����(C%%�f�g��&����60)^A������;I4u���*���t�`���GD�GW�������ѭ�"���B������#;w/2�>���9��̝yU[n.����h���:-���Ȅ�_�O���ۛot�>�3HM����E�]���T��qa�oaj �iS�����b�ה�$l	|*~k���2��������ϟco�;	[wn����+)���O�ӥ6�ڜ���2�|���Sd�V�Ok���,�߾�)5{����N�W�(%%%��Yt�^0KMA��mkJ�q�\�d`"����t3N�V����49П³wqu5�RMm�
������P��۱
��R���WM577�<~Ksw�C��P�Uj��3~�+W�]Rf��o˗>X(~s<!�}����uO��'�&۰�].������t�=�����xm��dk�^�Ҥ�������d�do�-�pԚo���*3���WS�_^Zb``�J����7^[[��ߩ_�_��3FX���v�K��}I�<ƭ���eZ�KB���]�֛b��xN�yV	���OZ���k��r��E���`7�-�NH���,Wϓ�"##S=>8��Bu�Ň��H�y�ϥ��2���������)�������'�ؙ�oc��ɓ��<[�M��6�Vc�����<��:o��,!u��5�Mp�9ݾ`dg/�RT���=���}�W�|��Y����<n00hl�'�:!...����_s��R��DFE�8�T����h�X����O���/1��:\��Zȣ=���v5����ίڊ]p"^!�iIII�]]]�w7�333��sߜ�����-�b��};�_��Rq5��455��.7����#k�~)x�;;���rր�-]�2~��Q��aYg?{H��Add${�A��M�aSh�U���t�F@-o�༌GOOolN����!:\���۸x8�&�"nчb����of��j�%��Z�ո�_���ߩ�����O���#Q5R8�`{�D��=�㡾m����p�	Z�,�����І>��<gf�0hr���[���"����N��ܮ�`��Aˣ���q��|�b�;����1�#���ߑ+I���on[}�d��[�Ywvn��n#݄)#C���,��w�4��OOO���J+*��F�&s5{��LN�^/u�d���HUᓆ���}�ֺ�7�)2ǭ_cmރ�sc8��|)�p�[S���\w�P�--W��T��x�Cʩ|�9f=�U�{�[�>~�X ꔉ!5B����ӧ/666Զ0,���
��}̀��L����;X�S*8,�z]�|���a�ٚ��-*�r �Ξ�Ϳ������և�>���y����F�b��|=���(U�����)�<+�!G0:UWH�����J��Ȇ��\l�V����?�7(�����HN����e���$N㋦+M8��T��8���°��aL���7Ҍ*k��2�>Mkjk����]��oK��P���q�Jެv�QRR����I��;D��ymJj���e�,�<ʶ_�&py��otF!����� #
T�m�cӖ�{�;[?h�׉L������f���KHh�v> �iHU/�}�@^�R����������\�7�/*����>�GA���2�;3U��[��.$�_*l��v��+���~;y}��yBʇ�������6���E�x��h�)��*�p���.�Q&fff���H��(�����>�J�_z�"�>11a�݁I'��y�'I���_�ƹ_�N�v�05����@�\������\��XRS3���N?h�+4�q�d�.��/5��QM{�t��W@sz<MLK�1wsuM��*p�%�T25]�-"&ⶹ��铑��qX{�������m��b#�"{{S�((��nz�����H��uGT����zb�=622r�.�x ܄�NT�]���j/�vM�T&$���Ta�?�3��%�ƍ�}�˝:�WW
ꨰU!q�Z�*�6�^�k����6�R��_\<�t���C{�' C�)�.��k=�ew&�>Ua,1ۋ\K8\,�k"��ww?�5���P-k�E���B�D��B��H��/_����b�i�wZ�GC�
?!Ac����E0JHH� ����w:����:���_-###�G2�B��'����(`9��A�� Fp��x}�.���Ĭq>���WMA0�����@�3�8����B��=>c����B�f�y&)):���|-tŎK�ʧ{-��ǁ��w�|������n��۠��q�[<�J!s��b듬����Ԫ\��|,Mc��x5!w�HZUU��@�2�P)���ȷ�9�G�0�ʎ��®�bW�ۮv�� y�a�kb}���R1�&凍 �Q ea����Vș�(�Ss,�:�j���1��?� ��{�ݜ�R*�n z�g(��J5�yJ��*�)���6h	}�����X����ï�9�!A$2�/_��&n\m��f|���cR�4j���Q���o9����7{�I(����"��1�������}�'|)�PH�s2���p�M%���}��^�ծv�ڑ��e72	�s�+`|\v�jl����0�Dk;���"S.��?��lp�`�z�X�)�������"�?�̠�q`CN6'Kkjj�������w��byyYM�XW�\�bz8��[�8
�����xs�-��"MO�V�+��Wu�뷋:4��ӝ�܀{���t���&���#�Q��sL�����Z�2��L`#� �N�� .0!>�k.�u�N���E���������y�eZ�;F�%��I���є��8�M�T>]]]5)"^�ۈ����W�K�\�����mj���]� �V�rZ�9.<�X\���p�!�r�cYP!���Y�<R$i�9�k�3�t^��f4�H6a�V�v<f��<�J�v�j�-��>����T>���E_��R�d�UR�U�75	9y}����IJ�\�W<�P�\O�1��EnA�P�@5�t˴�sss_���?MHH0W����L_���#��܏����������@|����3��=C���)� �S�'({Ldd1i�����<�GsQo �������1���M�G�<�����:W.Ow�7�?�r:Z!8&l��l%��� �c��m<-����իW�vS�b�@�./?ObfdIب����y���RC#��!��6�<��N<�:pd%gk��43�R��=�tbi�tt��6N>��1{Cݣ�{��MUv�ʤsY& ���.%�\B�����+��W �8MϨc�RR|���8]<<�ʴ�>m�5��pX}���DX���ਡ1V��Ç��ff渖�;佪�JH���|5�RK����E����;�.l� z��/����8�D�x�\h{��d4(���cވh��J��!9�0�	����E�|�?� ̉��z�^Sjhj�{�C
źrqqu���$���nd�Z�VY�S��A���=~�qqqA�߃���o�}�ߕ�q�3�6  ����._������ο1<B��[e�(Y,g#��1�i{��;�X�� �/8)A�B��-f&���x�9�|�S6a[�e�OE�uB���p}�?�?�ߕZ����~��|��5jh�X�ˍ�mm���+���L������JF ca���,e�98V�̸���%}@�eK��]��p,iGG��	�_J0�@ԁ&�<��!����ġ�����3I�]F�Z�������D��.�+>>���W�9}}JY_�z>?s��\π]��I�kt���^�e<�� �с�'�����<�z���0���b<����������r��ݐ����$/+��rCVk+iTf$}���3� �t�Z�Z����f*7�'�a.��WYU�}�Z�lCr��c�j*�VVVr��*���oXi"�褼O����} �1��3��������ͽK-<'-�;0�q�^P�Nw׻�����n|�_7��I�7M���1䵏$!%G[�^�2�&�F��X8*�9ޜ,цX �+/���D�������=E�m��]X�jT�/%فP���l���O<�?}����a��yyn����,f�?�Q���T~T�him��`z�T��ާ���
�}�K��� =껻~��OHI�h�:}x�Fj��(�+�l>w�7�O�C�純TR��e���>Ѭ�t{sU�GO5$���n��3�����?���ٽ!g92�Ѩ�5@����6c���i'�������7-�'�q4�.�!/���^H�}5� �C@%��RuU���{��me���~���H#�o�8��/8���������A�4���>2�--�^鉥�z��h�Pk45���X��L�/�a�e�I�z�7`Y��w4�8K���Q�Hum�;]-b���dQ����ޗ3`��+
<*��G}����pŧ3��4���V�W�0���`��1��5��V���ͱ,���_�'�Hl�7�к��˴4ٗw�f��S>��7�u
���,}Ę]�.
��޽{�o� g���es{xk(�VD�t�c�,f�gd۩��M[I)�����膩����f��@P� ��y\PP����}Ī�Ѡ�;�M��QY�y���V�vc�G~nw�/��<��.���׮���Iʡ-�uh^	r�M��^���gf�g{���V~D!�E9�����<�,�L��b�m
�e�ɤ�󍉤 �ρ��v��(���=��3?�0��V����-�EV0m	�Q���411q|5��,�
d3 ����4�k�Ō[|<��f������U�^���0b���܆���)F����
s�}G�$��0b�e�7���!�]h�  ��]��L��qtb��K�������`���������~g�L"(2<�տ������ߋ���R�Sq��U�;@g��m����~���; �����*!�s�3��mo�D��E����.<\�22��'���Vqq�x��~��K��d�t��q�%У�)�z�,j�-�˙YY�6Ֆl����[iC�w��4�ڌ1O$� z������4�Lp������x���x������w@��w'��Rfx���|��5O5R��H��U^�H���3�/B i�шy�&�R����S�P�(���77�B��O_o��R2hD�K�r墒�/�Z�Ѷ� �����H|����#羾������L}��r���N�ݪ�����5Z��@6�_����h����m+�}gK;�������ps��R������/��4�0C�j�ܻ�i�:���`�֟��a1[[!��1e$`�����~�՘g�XTL"�ׇ�<�O���A篧0�z�`��q��{RPPDx4�_��&7�%o�9	/??0��.a����%��b �9�\\��[%4l^�|���6@���(0r�3MN}@�|-;lB�M�C-�o��d�^0~`#@r�������B��a�/��J<�Y���X��)�������z� ���؏I@��{�%�ܿ�ۀ]E����'��^xi���ҡ����Q"���A���FMCs�I>o�����[C�@LLL�X_5��e������S�����l�p/��삁���%���}Zh�&%��ud9�کE���ӧr�$�k�L�gs�^�gggc�t00�)�|u_z��͏�d�&鳍/Oܘ9hS��9{[���/!��{NNΉo��ci9�1d��h���������:[p���L�6�&s��������ۄ��EX0�0`���㬻�q�k�^�kv`,ɨ��"u$M�w���gt1b���$NJJ�F�'$&��q��)�	�],�,��.�\���O����s�W��jY�V^��rP����1�p�T:o�ҝ *6� �,�'���2�]Ű�����Ys���I|q��fKd�t�oǧ<~��tg���X>�����q�����?����K�


*���?�;Z퉋��%�
lؽ@�B��bcab�u�"�)TI��eg/&�y��j�����g��u��1 tQb�� d&^��.�݇����)��"���F� �#)�,����K����u�ݜ�R����'N�����〛� _��:N <�H����>T���6tO[kjj���<.�A�����75#�9��?���u�e?�C��x�!��g�>����ZXX��\_���x"�X�Y4���L^�y����m 9�S��@#C�N�4hS�z��"7e��d��.�'��ym�՛[`�m����,%%��I��K��|c��06"���(f�ܙ&�0f���i�=�hr��'�Y�r(C��J�`m;P����||$j�v@\��}�6�L�����Y���O��ށ��l�W-y�N�j��G���ۡ^$M1�Ʒ��� �[��]�p���ɖ,<|>����E@<{w+�$���nz�l�V闭 6����L�}�f凡~٩�2��0��!n�J�r�D�*� ̐ Sӕ���=��{����u����=���W���OH�2����?)VA�&��A�����J<���n6z�$O>&!3'{�4��= �7`eF�����Rn�+�ڞ&g�.կ��D�F�J����k���5�^�?���ò�!,,�16>���1շܮWmi����'<F�(�}��ᇠ���K�A��N��.w��\ȹ���_�^����t��� �����8Q*8+�P�K�ve�B�s��e_��򹿍�����+��_�v��B��:�I7-��﯉M�����^�;�<1�3�4<�t�o���uB���}I�5��ǖ$b��'9M�:���,,LL�'o������?��t�@	�[���Lo�S%հ�쪛g�_ �?�ީ��bݜ|0���'Ҷ�m���}
e
�sߞ�|��������u	 �
i�W���F����u W�BY�gV���tc�?���x���a�}�2W�X�=zD�5&�]/�����ϼv>��p��Ĺa���� Z��9�V��֌*�/e�5?8t���D�ҁD�YPh��fV�����"6���u���������v�S+�U�!����Pf�����7��Z��fMQe���=��o�	a��[��%����e����ZL�ؿ�`;B��������dei�o�,}����&��g��T@� �w��R�lw��>�؄+Hx���i�ɲ��4i�Y �������=<���ue�(|���&5s�y�1� ``�"���k>�*[r`��C�`���K*Z�)���=��H;A��e���
ϰ{�-C�U���}���@���I t��#�)$����<vO��~�jq0�s���Y����27����	�����P:1��uc(T*s�*;�^����g�� �p9��~WG�QO��UY��4�X||R�0W�@�-��v���� ���~��'�mM K������e>ת�����Q%�Ck�-@�k����EX뗯ɞ�A�GW�C��)���a��N�V�{���3�\�`h4��iMyឈ�Yu/��m��9�ZWXp�~gs�����3<F�B��g� B��=PVTL]�sx��u���gO]A�����}�@���>�AP�YлT��mm���\q ��a�S0\�����rF2&&$TI� }�\GOO�|��a�s���qH)�E�
U?�:P�cWX�2s�}O&u��/���~�9ޙ�0h��B|��2CY��XD�'��b'������&��}]M ��O[�����+�/�ͱP���������iļ'j|�v��п�	Ï�q������rz�vju2���}��0++kO�aGՆ��^��Bpv6������C���4<��b��,àڠ�s���ݸ:ۓ��A�E�d��t�К�
	`����N!a
�G<<<t"����H���88�Ԡ=,S)q�.��M�iu�F |�btm^�Lx,��w��1����W��g313/���a#9฻�� �����:�U�Ym�������t˴I�}�[|�G�G�W���3}��\���a/�Cp
<W�?�M�����=_|�,,�OͣW��
�hbF�(%��8���י���ƽ�� ������������rg0NQ�'�?f�⟃��]͑��ū����L�.{�{[����k����m��`�r^j�h���WPP�����b۹v�N��8��tЖ�"��t�(���Q�����k�)��u�������---����"��������1)�>�[���@Y4��~����<��j�	V��@���h��y�����X���kS4<�llj:���C4��j(��K�~g7e����Óh(���=�g�}�D,Η�ݷ�+���L9Gu����>����_���<o�uggg$�ۄW���e�,9,,��K�U���R]]��)����& ;�t��\[M1oRW�ڏ6���>~�ݻ<��_�X|$A�o=��Au��&�`�w��ᖯ��Ⲑj٨5r$���7�ih��\=� Q�uҶ/���~�H��y�{��DJKK'B�Sa=/N<�x�*�����Hܤ=�����"��OU��1���=�)#%�A�����E�����"( �'O�i�d.k
����b�o3�G��p�{~:��G#|�DEK�s?���UUc>�+?�ܮ���\��d�y+vk�k^�(�U��j��B7��v�F-7`y� fl�V|=[��~��?=���O��j2}>\_ld��Y�K��SVq�d�f��	�r���S��Qڝ����{ݧ]��R�D�-4�	11��*+�Qa���5��vcؑ��l�n����}����,1�������۽2v�Zc������sNt�I��q�����dQ,hy�%2f��xw��������ۻ�4�|�n�WM��8[��n��ʮ�����Z��Q�fe�x읱���
�o�e�/e������t��T\̾|C�b9��2"ȧq���l��h�tXx���ۛ�E2���?6|�{��ҽ�����hJ9M��-�럀]DH)kͿ������K4>��������2�F]#ų����<]q��#e����IK�U�+������ig	d��@�<�[�,�Xr)ܷ����fF���ӔYV{�o����E�fђL8��l���OsQqs�A��j����s���Y?ABz��Ե[��H�m��+P����FQ�1|�ɘ.�r.��X��h�I��}�J>D.+'_�������u�~G�A7k��;cnu�E�gl�/�ɰ4��Pe��.��� WnV�����Π���SO�?Y�M;m�'�>-��y��, ��ރl��p����J��e�X����~�~]�>fH`8��@j�H��찬��9/v�5�U!����_i��#��Lyݿ�����er)%��u�5�ڣ���9�*Y�brCD�~�%����G��*��������R�R(��o^[��jXL _��.�^�l�͵�v	;��jZj�9::�k��S�
4#�v�;�K����7OM����������Z����7���|g:�q{�����*smcڐ�:]Ε�9���qNӪ�� 1;|�<X�1y�\�Iك��3�!����1�b��q� �T��b���Q�oDiU�Q˥ݸ�+���!��g$��;�A]]g�3��R����74����q�Ç�禲�dy�b�Wu `��}�a�~G�<���&��_�ܟ���?��}ZJ�E]�ݶ���P�5��:a}��G���VW����IԜ�9��G)�e���L7�}����xOγ�Py��?�4��O�i��5''Oaƪ��+��[�S�c�'0cͯț���A�������:h:�������s۶gr�D�l�����r��T��H8�V���%$$hS㇝%)���'�o[~���������M���	�|������1q��k�7��٧|�P��ڣ�9��q�,_lx�u��m���ݧ�%Ȩ����"88Ƌ'7Sx�wUTT^�U�=��[n<3<�[��uk�������pӷ����"�s�SaY��z�Y1�w��w����,�L)��|("�(�a�Ǫ���ISK󒌔�2�φ�o�V�]�J˙a��o��D�.[���
��_�
��nt�"�&�۱���<;�x~\��L��C~:"�t�|}-&&�.�굓��R̈́�u���a���~�4'YTa�9�@:��ϟ?�_a��~�����_خ���ѥ��Z�c��h{	lت'��<S�$ʥ�hr��餐��+����'Қ��1�/(vb�5��e�����`�\�:����ݶ�_�B9ri��s��)r��>ׇ��lR'�>�w�v�j��v��i�P�����y��N���P�!)����ь_Mg�K�y�L���2���ɍj�����l$輄�#���E���<� ��R���A� ����e�e�޹��:���{��PW�N���:�a@�5P����z=:�w>���|�o��i[/��A<PЀ˱_�ܯ�����5�y�50
ț�!��t�n��,zy}���u�Q����e�t�*iիd�u��.!��6��?z]]]��bb��4]�����J��� ����j�]Q�<�B��5rZ�zWKCR�/��q��āxBLp�����N�H��$P��{��3L#��㺜d�^z�@�GB*<��%�Ԉ��.��е7!�����p>�s:���:z�i԰�F�k4��Հ���\�yTQF�1oUQ�w���gN�1֣��ck�r.Wvk�2܄��Q�o���0g{�?҈�$,_���4%M�zT�T�IJ ��h�m¨M"����@	�E�PK]*�<��\���gv����=�%���)O�1�q`y#x�9�_����;��k?�&���m�7빒���K����f��Κ7܍�����,���+B"�H�]���4HD{mNl�sF��q4�[�5���ݞ|�)ϘT�&�~-���e���!L|�g�����m��	e�h?��S����&1��������[)H��l���6�y�;o&�:�7�l�<��E��~-"����.����|6%7�@*G�M��H�\�q�0��(����n�֟W�\���dBК�I�r�z]�ʏ�pxiC��<���zn%$0++|�k2Ɍ��=���k�F1�5��%��^�ɱ���T�ы���S��	C����Jo����R��<V������I)����;~P�J��H����ewql���kD�!���E��˜��_{�)��n�H��p}��wAa!���峔�,�m'<�]�*śx�8�4OH��aV['���{�?��+م>�m�{�2{4]]T(����oꊠ���R�Ü�-�dx]��[C��Z�Y��O7jRP'c��	V��T���\���@�_Ka�:NĄ�DgT<6��E�&X*���`���*��%�I���lN�S#��s�lqPKw�����`Ŧ��?��g�[������>72ߚYbƟN�щ`K���ݥU8ac��=M�=W�H�f�N.;�?4�L#���!�y���#�|%''�$�AA���>"�RH��ɝ�RV�Չ#*!�+\��%0�Z����q�DS�jjjC��Ƿ:'IY�8�ؼL��\	0e�(���j��H/	Ų�E����jTh}�H����[�s(�*n���3a�W��ϋN�hi�3�ʗi��F�*��Q��6���924/�:8�E�j��"#�xj�{Jj��"s�bk�u�Ox�X!�G49�v�X���I[����ᅯ�U��QB�a8�+���#�8�/K��o1�r��F�%��!�m1��Է�91��Qmէ|$[Wy�5��}���3/#��h��|�׾�J��]��p8\?�(������9z�T+���s\�C��%������w==y"!%"/���1L&�q���]�P��kм�3�,�b�%`�˚?Ĩ+�v���!K&%��g?QG���P�����Z�&�CZm>�s���ӕCY�ْ��O�/�8+ e�I���X�ظ�Ҷ�m=�!�[������2��$%t~�`���� FkޏŁD�H��:>6&�&�i�$�(#�E
'm{W�����J�R�z�ɜY�AlIM(#!_=l����W�`B���L�l�Ei��Wj'w�B�ԃg�aS?�m�(v{�����^�:�	�KB��p8nRrz�����$Ci)v|�/8�tÂ��D��6�&8�������U�"Kj��w�X�04m�|Q��+��ޙQrp9���f�/�$C!,�i�n�� X?��ů�D#f�ؗ�-�兛	V�F2Z����u�H&���EX�X/ %<)���މ��U#�Pg��ƅ���8��-�=,�����*z��\���&�G	��p��U���	z�`r�%\!*l:�`V��UE�l�OVp%���7dK�����������|�#���&�h��l�љc?���4���:�����⍵,�Hd���J��t���Ha�f/l������4��>�+�����eVYb�-Ŝ�z�Ѵ��h���P�	<��T�z�G���&a�3�SY�*A��P�&p���������cɖ�L�9��X�I��B�"u!�_Y�5ܲ���kC!a;��9�x���$#�u��$������1�'hK��@`�2%(�Ӌ<&���>E�;Nt4LRݜl�@&g��mr�����q큫���4�aЫt�f-(g��W�J�&�\�d}��W�ͧ�sn=�$T��#)v�Hя����N�mߌ��K'a���Ǜ�c��p��!�;����Pj񸓼`�6�*t�����"�K��>�Mv��-�#�Um ��Z?R7G*����/���]"G�s�~q(@=�=�%��@�+�/28۳T� �ۇ�����C4 Krճ�G�`����D�H!�LV��B��'Wǖ�s��[;���Y��=��4��ja]%���C0�j�o���?�EM����>��ɑ��8���0Z����/����P�V�N
�ڵg�l�8�#�#^t�-
�31
,�M*MUň����ŋچjx��ݸ6|p>X�����9j��˼4�xL���⤚�[\����q^Gk6#UtҘ*�;���4��y9*ʰڎ1��e@T�1�N�eh�^�m�`����@��TC쁒��r2�H���ȐY��"�R
�F7���#"�>p-�G����s@xC�i��a�M� 1q�Q$1���뜎�gnc%���`�\S�*�I��@�M���=VV�mq)��b
7zK��eӨ&3Z�|	�z�i2T�G�L�;P�=����L�����[!2ή�.����挪�R����-b2���J鎃��{%ߴ���~weS[����}|~�Z�:A*[Y[��DS2�XkP"���#9�_�^\J%���H�Y�!v����RV�['�utDϞhY�]��#����I��ڜZ:�.RK俅 �d��M�rlW·��d��h�M�e�%{��:a�A"$Sh]�ƶ	#Z�aB��dZ����]��=�U�b^��{�;or�Jl�A�}J����n����f���Fq۝P���,D�����(f���?��{jH��1�
���z�pNN�)��J�`O4�je77�m�G$�̠hcp�W'����H�΢# l��B�2�}hF��爵~�{B'��Db�%
���7{j�$�`gg�ȥ)	(V)�$h�t���VU��Pbt]U��K���	��4Գ� >��GU"Y1������T��>|]�@���3j�q�/,�Z#�)s��aP��=$[)��}���ˏV��G�"��;�k�A��Y"��au���X!Cd{D0Lh�($k�$��;A�����*v�ע���:b�GG}�1mo�s����֡�n]���t?+������ք|�]��pnVy��%��Z�i��M�w��n����)�;J!�a)�3���+.9+:k�w���N�$����@��u�������e\S�u�˂�`�2hu9D�{C�H�Zu��;$� ��$s�ӄR��#�Q�
���>o;[���v$4SK)f�Р�[�E�V	�y����fك�!������G_�ǣ&��J����V�92f�OM�X���f��&���n�h&����t��I�z8<h)]�(x#6��f�n¯���j�I�8I)�`I(ɶ6�R�4�)PR������yH�������>}��ː�T�XZ?����~�����c��E�	�X��SL���0G:�1�*�4�s�\��Ϝ��?�=��Id�.������a�S�P��.SL����;�lJ��7��8O?����{0��h�[�c�\��XNX��C &js��;�l���1[�Q�ٳ���g���_�V�_�[�K sIJ=du[�I6����fC�ݕĂ��GW�R�n�L�X��o���-�����G�ܤ����H�0r�QS������$�p�Q�=I!߾ ����P���y������,�&*$J����D0�KC� ݚsV�<]]�?�`�<�#B[�3
I��c�S�1�yt��/�;���bQ0��ҥ!����f�긶���z̒�?)��Rܽ�Ц��KП����� q�Qu�oP���rt���pّ\����pB��Dw��GA�P6v���F�@V��цh�fP�)�*�xp�}S� }�wK �����i�����~�6I:]�rd9F�C����D���}湮'$I�!^o�WS��]0U�bE�;<��oˌ�A	χh�$�L&
���}J�Щ�1I��+�c`S>���ž�M���!��V��@��#��3���j���x�\3��c�4wA���L$��G��<I�W��#���0��7O�.)`(#��yi7S����������w;:��&�&�4�}�IR���,+g�#�O�6����^	�����Bnl���� L�\���U��Y��ώ|DږB��3�6p�I�������ʝ�=��#�5�q=��k��ܰ�t��@���C��dc�O�v�������pb{|�Ah~B%�?�����M';a���"�!881Z4p����	v\\cq��>i/�К1_ߠ.�Rm��Qt���#JK����U�����
9¿�0�Ua����P.����D��$��ƿ��c+�ָ}}}�8����>Z9]+I�	3\&X��^��2���ڇ�)A�P֯��	�uビ��!F����]l&�y�Q��]wDN^;{�� #���T���"�m[��Pi��`#9�e��L���WI�!YC�1'Gh�c,�q�[�U2�ݣv�_*�M�B����I83 J��D�����u�b҇K�UE��ݕ����%āe	��gZ+��|�
��ځI�&U�Je!�xX�C��		���MhX/��)��L59�T�vԠjc���E�Yev�{E��hOs]��Fٸ���C�e,6���){tXj�}�_��7CE�|:�c4lEw��A�I�O�"H�T9�Z��s6K���/���I#�@vb���U���pA�O��3S�'5���o�n�� ����~:�?��ݣ�*�+Bf�z������eD	_Pz�ҳ�z�-D癌A��P����L��R_�D3��]�v`����V���Xh������L���#;Gzy7�+-��C�a(y��r�:�^3x� �iWP��&�d�!j�7&�3�-Vp�fPE89S�s���d��u��e�,2�Զ��w������.�t3b���Uh�1����u\�R�="��pO�6 �VT�'�߭+�Wp�1�◬6D�/�'_����3Ʉ����_9�Q=�ٮ��Ř�f1#�eMe�0�1|�jd"HT��9���Z�
/*�e���,QR4����x���\EF�R�	|t*y�$�`��T?���i����h��
�%^�����������Dh\����N"40��D�����#QΖ+������α.��i�m-��H��v]#|9��G�s��-�����T�&�Ry�h<DH�..fru�g6���	�^r����8��M��m��cHy(LF!!�!��h�+�JRZ��J������r^!RS�(^�S7d���ƤFW2��{ =�l��de����*t���ُ~�������ڠ?��P�T���������n���#޼�R��ݎ��da)wc��RÂ���8���k�rR�_�\w�&�8��Zj�]{�{�������.�R������\%	��-{VX~��Ʈ�R��f"�tO�|H<� ������Ժ��B6B8X�p���`C$LB�/1��6��1Q����/�@�ާ���3*�I�g�:E:ψ���q�y�';,Bs4_�~�`�o͟&09d�V)!��Ù�=gmy��dP+��M���t''��o`�Z~Q���-�Fm ���$���^�ZJ��?j�B��^��2<�����I��̡j�h�T�O��ͥ%���?@���� z��6f��y�
nn.���&+��K��� �R#��Bǣ��\�ϲ�!d'II�8�C%��RA����ٽ�0f�P�:u2��Ç���ɓԨt}�;���p��
,H`�uq��Jf�D�_��;I���G�x���C�K�p�@��Q�$�d�99W�%��k4zл{���?��|	�(22+�
[>��Q'�Al�[�W��0Y��np�O���u������|���]����O`��a�]��Jp�	 �`$�X�Ձ���?Ȝq��������W�H�mNm�AI}�O����j���VՓث�Kf�`1@_���9��������i��w�ß
(�DQ�f׉V۾?�\�Qd7O7W��-+`����%*�_��cc$Fa��`��p"�
�`�D�"R��IĝPM���V顨��w���m����0n?� 3� �@���������&��TD�F�T2wD�L�@	�d�����������f�A��*��PQV���O!�I�8un޾*�(�L�"0���(�mQآ?R�����R�	hU
�VU@e�Kh�2�gCP`�0�B���IRF%� &���?���ЌV2�'i�ߠC�y5��J;Wu�p���3QK;���+xy�@���<�)�ӳ'����oBDd+�s� �,)��+�N�e��[x������}RhFJl�*12��Q`�TUmZ���E��T(���3p��]�����n���Z�2���C�N����,�|0�˞+��m6�`���S)�e��k1bD�~��4ik�"j^�nRԧ��,���Q��ę,���!�[̬�Ȓ��;�ꈓԎ}N%�"�I�*i�*-W�
̛ݺ�Ί;�=QY��@֮=' u�|к���*��#1\�͸f�M��B@��JY���/��q�s�>~�Nm�G
��h(//WwOi<���Z�*�vU�O�^����sgZ��oZ5tT���
&�%m���S���T>�;Wq*sIT杂Y	àg�6p�ԯ���.�P��$��
��KK������C(-.��D�9�A��&*+�ು�C��0�^Ⴡ�PhV��R�wc):d��3��E���Y 5C���X
o ��e��6�%4�� �e��,�1��j�}A�SIQ#W70Yx(,*��s�������+���0DD��9.�h��If�`-�OE�f�\Q�.�v�R�o�r���g$R��F��Sef�qH$
��O�3Y�b���5.����=���� ��R���E
�R���UeЭsG?.�\PQi�����F^ԭ��:Wx^P�n�J���gAr�J�b�?��r�	И�B�i�altO����M��_�C?�w�A``pss�R�x	���бSg�>;6m�:O/�^^i���C�����������%g1�w�rh�2f�M����P^Re�����*e���z���J8��������Dv�"{�9���p����$Ю.Ɂ*�S+$S'��ضy���kP^ZkV�����W�����-"@��
���M�!�к{O0�"yLV�W%�L1�-�*���n��}cR�� ��$�� ����A�9�Dօ����Z��|���.j
�$'��ʛEO�����ꭶ���+P�S �(�7�=���ӗ�@��T�*M 
K9<��C��-��o7��� WO	4Pp����17P:�CJ������>@���qUJ^y��z�+0�*��.�f�`�)@V����%��h�@U�s`3p�rhX�z����ʓv���&�Rx ��ݡ���K�1{�<+�'O�ʵ���]��?��Z��z~Ι9g��z�bH� 	N�Pܵx��\�/'�"���=�C�ۍ\���r��̼��g.M��߻���ܵX��������ޏm�Z�Wj�� ���z��ѫj�{�{���H��je���N?��|3?�^�X�7���=�0n����h#��o���wp��WbȰ1<��щvV���a��K�z!������%�PC� �At�����g�k�B8@��*��n)��^}���D{G�l�N4�lS���hQ�V���ipH+�C�1S�1�pݕ�a���X�����Atuuq�w�]0�2ƌ���~X����6�]:��v'l�I,	]�cn}�ڍ-pP[1�+E�'q���a�M�#���g��l2�����.�ɡ���;�lx^�8�.���B44��3G�F-��Dz4J�)�-��bw�9���wDB�{�=x��'q��"�+ �-�p�w`���X�e<��2e�L��wE�sWR��ay̡.��9����o/�B�g�aVgL��?^�_:XB;*�4:R����N������O4�l�����.����_>�Q]�����
��������|��V$����(*:�B�՟��9W��#���^Ջ�0��u|�;l�lL �͒��Z�PQ�����H�!������3.A
AE�*�y4/�M�d��˸�&���e���d;��P6�8�c�s֬�	>�>�;�o�].c�����ð~��^�3���?�G��|��%-S�<�R;`�&I��#�t����"�~J&�;�܌s�8[�lŷ�|�X��K��i�}�ƠaC`�]p�|�|ɗ����!�](58\^�
u(,�����ob���MU��*PW�P.��1�U˗b�{���A]] �Fl��G�=�W��&\� r�"J��OJ`�b)V�a��}yԴ �njօ��✳fa�}�EwG'��D�654��V)����]�z-�y���N�2|��;ٝ&�e��Q��T�k*|.'�k��!������T�!�J �r�I�x,у�8���]r9N=�<��k����0z�8ĒI>����Q,A	kc$1;,�r�+�uD>,[�-R==x뭷�u�V�5y.�cƌ��݄�s碩y ���y]�^�`wP��*���-���K׉���f�)��ˈD?	#	��Q�W
���M�����Y��j�`�D@�{a���3�ePS��z��E�v��ؽ��W
��_]r�����D��e��C�Z6����Kh��<|�58��y&̤R(tTEd���2�a$;�b�#������탒��E��W��u���������-U�f�������`�����X�b���N�R!�=��������f�d��U��hm݊�O<�N=�;��+V�+��)�㭷����}��a�� ڠQ����&*�$�,�"�����#�Yل,�8e�LL�v�܎Q#��X,�'����&ې/@��q&���7�x.Z�
)n� ����r�T*r�@؂aV,�0�r~���P�3O�C)��o��	&�2�s��7���[�	M�hꊥ �Q�yi,���N�[#Ӗ��iO�>�&0;y�$�ڵ?�^���D�up���a�
\z��x��W��BS�~���"Y�,Q[/��{�Z���k ��t�OS=����GOw���S���0����z�OO���ӏ<
~�9n�u6F��T.��`��=���L�������EC4�Q*���C*��ŋ�H��������Ǥ�#��WD��͸�������X���DZ*K�#J2S��!���Y����B�$g&�Dtr��P���[H���2a1\�T�S�}.u*���TA؁�|G�s��S��3�א�O����P1y��Ϗ]�#uzQ�(��L�l�R�TQ������Gx���q���cGk7n��F��i�=u���݁VHa@����<HW_w3�rlN�e��T�ے�i�S���{n�b��6�jM�4�����y�F��a���5�y\��
�m���Gq̑���X�XW'Z�l�%[�]���_��;p�=w��?�g��ѣ�"�Hc��/�Ϣ�����A�7�=*,�����G��`g����9��ϳ�m��{��~5jN�5�x��y3=�>���1l�|��gȤsX���'ҬQq�n��ɣ��"уc�{�H�*J���� "}����4�1�����`�K8���sg~�I�}�!��%4461�C��'}@"�^o	�7��ԕ�v�\N����E�\x�^' >� �s�Yx��w��3�`Ѐ�:���k�+Zw�c�i�qA!@��+�D��������&�4���X������fbؐA�����l�i�{�iL�ko�=
媀������.���tǓh���Ln�y���[R-eo/�Ly
������>
�V.ǁ�I{�+���'L��A��hl����1f�|��'\t��px�� �F�\�6�B�*�Z�Qy7u-�
T ��n���$.�\Pz����C�ob��<^��Dj_�p:��δ���q�A�^z��_)(dڛ�諃�\�v��i���Yݡ��l�Z�MS Eص,ZW~���	G<jA�1'���c�#'ӯ4gg�Z����HdJ8��Y@��:'Hj�T�)�m|��W�%>����3U��C#�4)RI�b�(C��+p������.�%r�n$�v��.ǵ�������5r̟�,Z�m��7]�ÆC����C����)�/]�+��&M�˗����[[���{ـFs?�_d>����EBa����l�.��a�q��p��ә}�v��K.�ҥK��܈|�'��8�,Kx��p�ɳ0z�q�숡��	��s+K-1iM�K2�)�z=�eR���=GB��X7&O��������?C��eV���+����7�|3����(Z*(JIE;H��{��%x�N���1�L4�a�L��)h�؎	������A��'���r����������K/���֮Ô���ٷ�� C���-�%5]���`0\��a���`77�㬳�@��@ѱcq��wᥗ^���0���sϻ G{�+:馛��p#��I呜�*Vl���6��F"4�?�e�X7�=
����8k�,�x�)���O�@_��c���B|���1jl�ց`]�}�<��0h�8.(Dի�첽�.�2U���汆�&�-V���WP�1�ᖊ��&+�ɺ���`���jp&Z��B�Zzm�����C[���_)(����ȿ|��j��1'gm�P,S��S!�9�F)��)��*�X�W_t6f5��>^\��}��F��<v�έhK��o���=��{���A$R�E�����a�s�gN=�v�H訸|(��,��_�`�c2�V��`�u�O��Y��������w�0a�d�X��l�~7?���\u�"sF���s��K/���lA[[�菧���eW\�-[����.Y"�B��M��
�mh���w�N��=�ဃ��@]D2��S���-�ۘ	�e����C,��e�p��g�PP������J&2\h| a�D�'�4�-��0��w!��O��������Ϡ�!��=#Gc9>�,]t	��n�����5��2�0z�X3�,��Q��
y6Z���p�I'`��Q�}�m�o�)��l���5W^����y�=�D"�-�6s7��'�`޼?�7��A��`˶�hhjƚ�롒�]��h[Tio΋5�0�*��ж};�>/���7��w_�13��Kλ�|���1|�pBA�?w.RY�| �-[�o�	�j��Câ����>/��0��x��h'�_U@,օ�?]�X��*\w�U������~�Z<�������G�c��pȡ�p����cO�M������+�c�]�#�UQ2�ձC���̊Ɍ��l4��295�}z�,�Uj^��|B�-���^����
���,W��6��z6b7^~މL5�_R��񂲸Z�?~����}�^�������f"#كJ&��3U�p�رn5���wc�}2
۲Ym᳗�޹C���<fs&qTPB-|;5 %f9�{#.:�d������?��y(���J��Ph�%�EK�L42����p�@�,aۆ�3��5_/�S���`0�-�[��х��\w�}g��<u�0�M���<4��s�98��s1t�p���8p���ں�6Y�F�M��A��_&�&�+/��x'��{3�=
���?�L:�ٷ�a*����o��N;���U?aW�|����Ǐ�G��x������BRnR��].c�~{c�q�7o�>���iL¢E��s{+.>�<6�hP�����1q�DVV�x��rx���[ǻ�}����.qQ����2����ݬS1��p�a�{`��'bԘ���t[^I�ү��Nrú�����g�}����lg����7�]vr�&�qV��e�����>���C���=w3��/
E����H���ӯ?�����Gc�QG��'��ƍ��J$1j�(�9�;�L�²�c#,�u�t������Y���ݍ>-ذ�'��N�p�U8��S�ò�����a�����#��i���3�矏h}3���Zh�_~��������dI���@o�$�0ȽL�XM���� ?�tO�I�q�ݔ�����wb����� Y�¼L^���IG��K����4�똃�xA�dcO�C���2��}.ؒVXTV("�e#��x�&�N7�G���ҾGL���>��9��\!�E�����Q.@�܄=�\x��C"k`�IgM#�9���z=�+e�z��6tm[�R^CS��>��Me�2��GU4��sK�%âU�<be%��m?�T�h��1�C0nω��,��=}�>+H��v�}��|�ɸ}�<���|��:�<��8���1�C�K mDQ3 ���pd�s�!�*��S�    IDAT���g��1|���1tF���������Nd�%��Z[[�՗���5[q�}sp�%"�N`�Q3pꩿCgWFY�R"6�ai֧��P���OcӴ%�56a��!��9�M�Cg�!����{��ڵkq�7�7��{�á��@{W���	:ʽ93U�d�N;�7oB0EE70x� �{�6v̭[���m'�]��7_��܋;_�D*�T<}�Θ�� :�\��˒t���Ib�B�� �P^�5�m	3�aS;~��زnc9�\-�8��sp�U�ǝwމ����֛o��+������p���u��lQ���:r)�{��R���k1e�Df��w@-�����f�����Xz������w݊���m؈t���o��y���tĉp�`w�����>�DsƝ���ez�����Ҋ��Bd}X����𰖂J�EX�v���4� 1Ll��V��ȥBv���f_}�����d�y���1�-^v]�;:+/�]�|B�m�x�yr�U�"�Ѷ�}<��=�>c�ْ�	g_��c�F�d�E�*b��aB_7^}q�yw:��Q�G�2�O��R:����N<��������;њ4��~*e�99�|�V��<N�lٞN��d��4mѷ)��ATh�>X�IQ���w��
N4��T��9�^4Z�-H:��c�Ġa��ڛ�]r"iD:W��������5.��l�W]r><6�6.[�e��G�@]�k�o£�>�7�541�h���8���m��/�0���8��'����"�8�CH��io�bɬ�
�O�\�������b��<JR77t�@�=n��lE!�Aߦz�Z�#F��)'τh/c�^{a���"���݃
?�D�Zipd>t�H��r�����.'����Jt�׆$�F�D�>}��7�p�7i�$̞=�R	=�F:�Q� ���!�pP�R�Ff���7$�3�YL�A*T{�5�U�k֭��s��pwu�1%�N�0�C�j�J[���ş-ƒ/��+�.ļ��F}s첄�jv�9���r3FޘP�Ǆ�`�h������q�E�aÚ�y�z̘1�uDDw��hnnƲV0�e�s���¸��'�E!{�\�y������#N��N����q����a+�Wת	�걢�Q&B�s-�<krQa�`y���f�a3�{�����\?w�@o�oRP��11��O��)_?���h�f�
�mY�Z��Ԫe��Ǚ�_��O?��ӧb��n��«n
O����_��Ӻ#Z<x���ѓ)��S.��a8w�կe�@�� �$D����
p�5���<��J$s�7�(8��������褌�����5C�s+��:���@/�X��x��'R�V5�E�H�$�����d��I���Q,�%'��DQ3ѓ���AvJ0�<䲊mkWb@c o/|]�Z��9�u��!�޺��l�Y�c%I�mwa����cɗ�cێ-xq����u���;x4�Du\�ˊP ϐM���D��A_�FB&	�Ӊp�>�d
*e�P��,YL���()|XdɆ��cɗ��ǟ~ƅg\����C�|0�y�%�N�NP.���\2����Jદ!�I��O3�{�l_ ��>R��R+� �d�I��y� 2l���I�ѧ� V9�0���H ���*hF1��I�1@}[�2�Do����1u���	G���lc��+C���<������U��Kq��`����(|�0�+$
ƢP/2_�D���P���e�ا��2�ʻ�ܳ�[�gD�����eH��G�0~�>�L$љ�C)��롓�X� �2����O<�0o��~�{�w�!��N~o�S�����^�x��M�̈́�P�oՄ�!�UQ��w�����58,���}��G�WV�����~���8�X���̤��t�R�Y��*yme�?�^}�a�^ظ���8���7��*�ݻ0m�>x�ȕ�8�虈�K�]~�1�
K�]���^xf��f�s+�K2J� w(Ԛ�*� ����d��Ө�S��HU(��=	�M^ UK(TD�]���Q~�^�$[���/����&�X��gB+*�\���׏�)�8<^$ rU!�itm^��A�'1��1p�`<��C����u�\~�,�Z�|n�s�N:�d��q�l��#E��b�%��J����� �tB�V�����e�@Q���S,c��R�Un��Yk������eі�������,x,����X���?RS@N\�'D���P畠�E|��G���q�wbȰ�(�L��!d3	���(����t4UZ�aGQ���y0?�(��hGw*�8�vIKCm�Q��4A�6S����&9���vKS3(��:��x�T(+�s�A�s��X��{�;x�
�b)�·a��o���PPx�A�0B� ��ZYD������*�L����F[��0rI<�ԓ�����espW ��I{cۮ.�./��zr%6vg�$7$��}@J9��Hǣ�կ�b��5~����_�ZJ���~6�R ��o�r*L��g�n�3zv��������'���|�A��x�Z?|F�RF�P��KAO�x�c�ae~Q��oa��q���6^��wH��Ӎ�WP̧��܈�3�@N^{c��A7��[h	�7�	�ƍ�V��KnÆ���7
�V�b�ح�B��J�!�+E��
$
�Q4��"��<$���흲IU功��D���,�͆���D���Mi�!O���y4#��?� G��h�B:���` �!�)���=��\�B� ���j�r�,,��k̙3���r��~6b9]�4K�s��]��sr9ې����l.��q�p��Y;���TTx�Y.�P�
�����<���[�E�g����e�KFV��i��94�;���P�k׹���!�<PH5�UQ��}��s	�	Ɉ2|(�>�8<��S���U�?hb�I��=	�b(�d�<b� :����j@s߁P49UE���(��}�٤V��iCۮ����PJlm
�	�q�`�/q����]�Q>�Z��D�����N��}�BWJ��bD���0�°e7czd��=H�:�+h
yѵs2��h�p�Y�c����xn[{7��}4�M�yz%ʻ�����qL�5�=�����{?v�&�!'�t�i���`�tm'�w4Yy2�B���)S���5��n�g���~��Oh���&���[���?�#O�U��/�� �E�ᲈ��b�7��W�a��0�tj����B�ȯ��!YvxJ��4H2Hq2��R4�l�v���Ǐ�.�#����hvzY��|#`�D0�����:d�%���e��ʅ,�F����(P���^�2yM��F-)l��:�Q������CĢ�!�AI�YR.9=��x��`P..	�L.���D����Λ|�n��G���-|��l?�#�j%���"l��H�LVS�u��P�u'�i��4�D����u��b�
ѓ�!�HB�eAK<��͓��k-8
��-/	������A�1
���n��!�+	-��ϴ��_s=l>/Ҋ��uV.zϽ�O�E_�-6llŀAC���I $f��3�?��6��Z)�6���`�U;��d����\L�g���8�x�jXX���ddQ�\�I�7
�c���u%�N��$�Ul2�}�!],@��M�/��������p�̨F��s);�Y"J9p��6CE:މ��<��b�q���Wغ���쁼JN� lN7�8�R�fo7b�����=Z�U�q����G������C!� y���Z�=e�H�-ڙ�ڶ*����ui=;���~���l��KV��l9-�U�4�ih�.�W��W�*$S@PT�s��x��8t�^�e�sɯ D��������L$�&�7u#�N��d���S=(����y��X��(�F���B�H�^%���5K3$U~�K�Z8�2�-�UȆ =���$�J���싂�D~#�Y��B��݉��Bx���ꔒqd��@i�e���Hs3<u(�ZK���'\��O0a�0i�����{�܂�:V,[�s�^{M��߬������/�Zx�w��h���b�$3�&--
��t�F�"�Jv���l��&{�M� �J8$P�aY#�Լ@�na�
$�7ExC>x�~��m�N�ٮbm�P�}3����� ���Z7E%�*�����7��fμ�\�w�(�^59���s.�ϼ��n݂��Cml�t�"�hl�� ;���x�Lf��"Z˨���ØI��M& ����	���_�����@.W`׭h�CrS'��#�ip#����>.H�u�m�ƣ Y(�3PWǯO�T��&�9ǖ��
��.'�=���hCI�P�2�p#�I[��neR���y�gC�Ro�1�t�1R|A��q�C��{���
c0��e��S�B�DK�OݢS0�K]F|ׂ����I�&�?����l۴���c4�<0Q��\,Y%�E-+6�z嗂Ҷ�<��l}聐�vu%����Arژb��2��;2t�T}v�Jn�fY�$�v ���wS���(���ǚn�PJU�VP��Er�R�`��x�)A�9Wuk��hF3E'��
CK�P���S��
��"c�.J��e[�)�������ٲ�7F�Q$�A�;�Ԥ�UɆ��} 8$h*����{�,�<�BOvn�������8p�}0z�p�|^��z�C���oP��E�i��r{9"2����a=�9�#C�4�%ԡ�Y����J�J��Oa���R.5�潧.;�M��f���#!!6(Y��Khl�G�.�xA�����b	
��+ZRtZE�,�R�� �+�G�mZ7m�ߛ2P(��K�W��w�N1@K�A��ɻ��3u�d�TQ$�� n6%�H�(k�������A���x����m`F�'��(8�r�9X:����#�܀�Á��4��[�8d�	�t�d�I^U8������<c��q�$rwF#6���n�u�1�|^�8�r�ر7��w3�*�鹳(ߚ�|�����h�v�����c��ն<���sƱ�h�+j]f�}�S������n=x��w�#H� �P�N�l�04+�['���h`�����1}�x|���8���7E(Fo>'��ۙ�#��y�#Μ�8ղ�;�"D#�{n��yw����i|��e_�@>�)��RRd_��sk�	�"
�@��`	2�ɬi��:*:E%��T(�K�/�<W�6�,#��!W�P��P�pG���6x=f��d
J.��N9�eT�64�k���q.��xE|>�%�a];9�iǎMLkRG�r��o���{r���u�������?��b��o��)���lt��p(g�S����I����X���B ���Y�rI��D�)C�PL��������S�R� ��F�l�B1��QR���ۮ���#h��]�er���h�������j����C B���ki���15���zUC��m���B�ݰ�Z�ӆܴe8~.(r�b*�r)���p��0X~׭��鯇X��{]�2I��^��8	��[�I�H�UT솊�?���p�kG�F���<r&s
do�)t���h���埢��"�M�9�e����tZƶ�Yl��kQ5�w�|�[D�}A�-8��f�8���n ^g��ƽ
�>U.(zO������߬Cy~�ƃ_�|�F���� �P���ٺ��tЏN�J!{=���O���e+V����E��1�d'WQKG��EH�Q����	��I5Y��z��~!����p�����h���#W��6�����
��~�^<h�$�(+��%�}�am�azP������B�h�%�w�BjNA.�C�X���q�t�t��
��-@KQX�S�9����M;�ac�YO"���2�~�DxZ:%Br;�S ڔ4%t�]�ѐ"s5��.�+t�
�q@?dMΐ�M|ɶn��%�%�8�	z�l�Y�"m=I�gJE��6B���C�M�� �G&���O]Ð�Q��H��*� �I�9�ɑ\.���X��m^��Őڔ�!O�NN@8� "�P���c66��!��������zr:�0%�M��B��J�V��H��*��E8er`�����C=����wb�ڟz��
����C`H2���
�6�U��Xd�صc�H�i��("���ۃ�b�Nqdu{P��x��ւ5¸ȏ���c��oԓɐ��^g3���vO���&��.��jvi{�z�bv/(Dimx��\Pj{jQ�<NAq��D�[O�\����>��a(�����\u��4�@*(eE��8ϮVA1!@��
~X������2x�#[q1O�Ӹx�'$WY�E"1Ԯ�k8ꕀRZ|=�Շ���Lk���F��:$U��S�!s�u-�u�p�>��aJY�$��(��kN]k֤��6Ɖ��@7��%a��T��4�bT]�R)!��?�E����݆d,�!�DZ���`C��Kf@�aB$�*�*Ҋ
7њ"�V1���B
���eH�Jq	.$��MPD�lH�����R�`7P�� �B�j�FV�2=L6��[R��P�;x,Ht�X_By���2Y�Z'�t"����C���4Q�Ԍ@CIS�FIr�c��U��Y���+IV�hc��ZAj1�����"b�*V�6�<U	롬���*�B���G�J"�T���U#��Ą`���4���[7�s�v��hes;�� h�aI�q��N�^�ߏl���V.�t�S�o�P��4�f/Rwf����1�ԭ�=�B t��:rE����a��8h�(4�Ml���ׇR�jO�������^T؅L%���!߼e��B?�FI$�<j��Ӷ��'�yh�F߿�0��P�g�ڃ�\���a�=J���KCM����2`m� �w���p�՗a��C�]��(bJU��.^�Y�X��L>|B�)��

1@nрd��k[���������ܖD��}�0�I5���F�>m�(��'t �@��tKZK�8b��bst+�^`RPRf��ԫܢ�fBU�h��a+���ʰ{��Bt��~t�@U�y�$SV(4�V�����.d�>|��A��g��S�K&-����.@����2f�BQdz�ѱu<��9��#�5D���
�䅑Ӱk�fH�
S��h3��$�uN�YCy"e�[n�X���a��Ayi�i@�砤�y��@}��Z�9�o0 Y��튣O*�J�j���.��켲�����厏�v�q��L@��؊v�Ѝ�Wt�d3M�h�X*~��\M�0�#�et�P�qFWs(*YƜz��b��Mz��./�\���d�O]N���Ǚ�u����v �*�~?���;Z���L$���k���G^Ӹ�"�\+kܩq1ի�ő

I�j*)w����C�0���b(�_Jo��-(������G+�Pȝn��T%x5^Mw���w>8�����<���C��Æ۵��ŕ
*�(�����W+(A[����?� N:j��j=θ�21R���Xa����ȗP��TMikUm�ih�܂o5����:R�2��3��^�)�$�&a$im�movn��P�H:4��A�cIW9��*8��'j%;�R��G�O��%��C��> {�O�J$XU2J+������%{�4x(��n�Z�a�/2����a����*����E�$��k9E9_5���tIcA��Ϣ�Msk^Њ�kiA��EE�����☂T��#C��X6���g�p�	�ոC�Cz}��$�l����f%ލR2C������mA*��D0/Yﻒ�t�-��턫.�,X,�f���'�9�"t��jpA��_t�N J���,�wQ��ݣ%+�Բ���B�fG>WD8a6�Է�����`-�8OG��Ќ:Y�P7�� ��.�[l ��o��\	���8�����SB6փ�;	�y=�7@���|H��#G]1r5�1LT�H�L]-u%���>@`s͋é��Y�R�H���g�N�L=.    IDAT�_�<����>�$UY�/G��xP��3]�?���I�B���^�_����?��ٚ��\���~�X����e���9���t�ng
�e���}|�֋�:�_�
7ιjՆ�N.J	nZ=Am)6i�#T�n�ZQ�~��������C'�;�����/�k�J���)"��#�mZ�6������Y�]�M�@�:���sC}#��=NF�)v���.�bQ?+�l%���F^6���I��&��Vez��Vx(��0��!۪�n]�T�V�����i
p;����4�^��5��~%ry��ݜW��w "�}ѓ�C����ȵ#����Dd$a��(Q\D8���Q0��U6��;;��耍R�+U��5"�P�"�����2r�"�~��x��(�j�]��%�e�(��6z�A�8 �X�M
�.t�lcun�:SS���#ʽ�;,J6`��A�cZ�U�d�D_P��p��-�a�X���â�ʽ���K�qE�y�$?�\U
y�9��+srs7j���I�5Qa��Աl��MT�9������pC���VBO!_��љ�-��Je�w��Z�~#�z~�h�!)�It�Ҋ�*����p;�K��9@�6J�H���a_c)���WPz��_�<�>��u�s�R����՚ِ|CN��h�@��n��G��oUP�������b�ZtؾTPh䡂�gb��)-
�.������X���8�=�a���o �l��逩Pf�E����r'�FK���՜T�+F>��`0��&��KnC��A��f
)-톅�32Ϋ�=�D/�ڕZj�-��P���8�-i�L�o&��v�l�ݼ�����MkWa��=p���q�}�~2R<B�;�T���c�� ��dry<t�HwlA�����?ގ��8�� Z�@�:���}3���Ô}���x�J�v%�k@���`�8��a����i.r�����P��^�"TEd�c�ĺx|��6U�}�xs^N38o���Sw$I~�`�R�]Df��b����'�,`���9e�D�ڐ��9Q�����e��w�״Δ�L�t��M�@�g��lG��G�~�O!��JU�F|�����0+{�1��0O~Rh����r��OcS:OQ���K�[�J�������(�n�ѵy+���%(#<�D���0d
e�Pv���>���вi�o��l���f��x*͗mŌ44��#��3�$TS�J� ��2��>��J������ '@ؿ���:�}z;�׾����X���"�bs�����
Z�RU�\炅��o��7�P�g�O���l��Zݰ}�&*E���D���/��TP���u_��J�i����N�k���5j�D\���b\�M��K�C�mm���0��`��p�%�`KND��Fs�M�B���TMG�/����(��R0��ގk.?�:?��x�oh�?��.�P�:�;��pc�gc��{੧@�r�Bud/|�lɮ.�F��������[��A�)"�c#R������#cޠ���YrO�?M#��H뉑��7���c��5h:p�X�R����!����+S�.&ҧ	��z��mU�����P�Pp4�4��[W��$�t�PM}��ΈߋlO)ZA�A�>�PH��H��8/�Ă$���'A�
5Q҅2�]pVu�h�q��`��ٹ\�T�ã"aL��7=�0���n�x��=A�6'r�u�)���YI]t�Qʬ8��y�PB&�aQ���Tt#�49� Tz��QĪ�-[�Y9�f>w��M�WE����I![�3�J
�PS3�%�́&%���(��:�Q@l�&$ڷ�TL�z��G��Ç#�h����7?����V�J��Q�C�h�ᾡV48ݿF���f�_����D���cu:��;�m����q����l�j)Q�t.x�����$�6��ǿX}��˶RA�L��h(�0Җ��i?��>��]�����n����B-*|��CBf�������:jSE��D�Cb�pTY-�01�
�J	�;�3����"�����䶥�Z{��G�.�{�F*��Q��6���gx��'p�!�`��x>:#�폪��F� �YĮu�qԁ��y��ڌL=�B�uM0�^T�6�E	�L�;��)��.�e�T.���2��i�W�\�=\a/�l�s�
���0����@��
���J�|�:�Y���ƌ�V��p�!h&������MK�(��!�e� ��/k(fHv��\�2[�-}8$��F�����[���Kqґ�c�ɓp��O@tx� �)�6{Xz�w��s����O����^Ɏ��G�m`Z�L>��R��f��N;	3�;���M��=L?�R��M��0��4j�j�h,��<�8N� s#��Q�/�C�5b���X�Sf��(ʎʮ(^9�B�*6��7_{�;f|��r����!�Գ�WUu�n��C�R��!#����=KnY���aHS�~�u�wƌ
'��D������O�|���|p��	7ð�P"����w�΁��/�����5�W��������pr�n�6"=h䡂BTPdҡ@MV�]�<�����f,�c��:��+�ܦ��ؕ7 jԥd��J�����!�K��;��ȩ�p�Ga�ؾQ�Ȗt4���Z$�b�7%����("�j;e
�'��sJj'�<�ݼ'�3z�a�D���*�~� <��)[�(q���r�h]�.���t�)�FDS����-x�Ex�ax�()�[�⬓��-W^C�����[qڕ7�~�X�=U�bE�u9�EE)��\��D�?�ɴ=�v����΍kгk+ҝ;�f��PDCc�H G5Ǟx��4��o�;«Ywā���~��E��e���V�Yh�L%�:A"%o�E�(�8�&b;��Tu�l$��pA���e%�d/s�&�^���S��'���<�2FN�I�V`c05��V�0���<�o�ø��fhӚ�0�
��~�)8���1v��m����i�<��@g�p�F<��˰�)�
(Q�&$�IM�(�,ֲq�j�\�Q��H�o����6�\v�X�a\}s�O$�$�r�o�8�8����}�?��G���0T�n��{b�������Mrqf�+fMSI�!�Ѷq���~�E�|iX;�H�L� -?ZA�]����L9 �D�"A%0�n�e���_[���R3.*�K�����!�*j�inVA��<�Z�� Q#t2�&�T���̽���D�?N?������b�5:t�2"�9yhE�w�q 3��J�DJ�8v�~8���1�O3��|�o�؊�^��}�X:�T�r�R�gU�`DmI�Q�u�V������(��I�܄�BV�Q" �T0U�CC�*j	�do*N��3�C��P�����S��Zex�p�܇P߯?vnۄ+�=��w&|Nb[���U����`��`�#�U%��K]Y�D�鄙ˢ{g�J�e�cF�嵐d$��ډB�U%��c�b�~�p��S����UD������Jl ��ܼ#���-#ơhs2[C�R[�D�)A65��|�o6��}���s!��AC8��xw4��P*��~����0�$#bX��eP��?/�}O>�Ƒ�$�:�GUE>ޅrNa<���1t� (�$r�NL?t
6E�xp�	���&�9�IMM&D��<^|�=��ՃE�/C��D[�RTf�d��̤|��b%����αQ�	�{3�E�x{�<~߷�UL?�R Ԃr���O����TF��8p�<��md?���9L�~�M=��	�<F�ٞ��_����`�i����vmDsH��݋'{��M��ȗ4d�MM�Ҩp~��z�~���A��"H*V�e��V�iu,2���c�n��2��
��ï��除�B�Iz﷕SFrׂ���и���ǧ������]ykv��G���TT�g�X'*Z��<$�! O(W5Чj��7�#�!S'��c��aNE�_��\*U���՘������o`��8谣���7��ܾ���y�߂�
\����3_EvnI�D�0K�k-�l�$��	�uK6��~�b�P��ᜓ�����5��Q�W_}���=��ē8񨃡�h�-aG<�iǜ_�`���T�|��(�w>����l(D����n�����A�@!�Č���I�0n�`������\�<�����NЙ�cSk;��`1�_�C�L���#�@������	V�d	.���]�H%h'3�	�2��h�，I���8[(�DVvɆ��A��.������|6<������E��	\PD�fEynI��iiP�)8m�~;�=v��5��A�y�M�5݆F��K���f�:~��:� ���D{^EF3�%�A׬
��]*�j����1K�t���}����q߭W�r�م��G^E���!��d�U��J���?b�o�_c���']�V�gc_�����Ew�vtmi���e�$�=�aDv���#<��8zھ���#(_{�}�o��r���ࢳ��u���9W,c��'C���;
Y���BYy���,*�0(������Vj���Ձ����Ķ�:��{��l�ZS��'���/�RŮ���7�}�F���2��+g~�v��B��8*(U�&�
�.TT���ݼjD�E�������_B��F���Ba/.=�Lz�hJ�����5�hѻx����o�>CG!\׈����Ts�K��B��`�Y���t�z �o�R�iT�	*[�`Z��Fu7|z;~��3w�~���P+!ՙG]����(��U�pޕ�B7#�4�{4�e8j����bOk{H��.(�4�0���b�w_G4
��L�PAٵe+75�m1,Y�;�Y$�%��l�3���P�2Ҵ:��]6��XV �ND���l"�B&��
�ۉH��Ӄ,$8������J�-_� V0jX�H#ߎ��~>����{�<��N=�*b'h#�R|Q���ܺn9f�4���#�%���M@��Le��+���k�x����8��0��#��$��&���e8H�H�Wm閍�
u8V+i1X��������־��%�w#� �@�a���	�aH� ��:0�����q��t�Ӯ�]����T�;w�w}�}����-�������H���m+���KN��sO$O3c֍,kJ�8��LH�~{��)Hw�2n:�.:�TbI�q��j�s��x�,lv�Z۴���J:e����-�����C�("Ms�Mw���1{���O�/�"��Mg�&n�u��=I�Z�ճ�d�d��Znt�w�����7 �a���fT��?E 	����-�����L����H˶ן������(�������?���s��tD�ZD~_P�]c#��X���+�jJS`3S`�Z'�D��m[�u�Hf]8��&O�'��t�vx��oy��/�e�V�%:���Z����=�KF�����aP��6y:��0O�
��ޥ!W0X�A��cNRf��I��m��a�Nc��gS]QH�O��	��U��X�q��r,;��D�>2v?ᄬ��C1Z���"��< �l���&����#��u���T4��5��%��ױf�fVm����*@kr8qz+�z�t]�09U���ۋ�#.�9�4J֛B�/�h�����z4�ĒNQVQ���B��\&N�7H���T"A&���(Y �E����'���;y�����3i&�7�C��3��Y(�Y�j���f5��/�|f.Y�f������՛�Rװ�3fp�W+�����=���#᫤;n"���rz1�$�@��1��S�'�v��F�8�Q��&����R�O�q-� 	O%	[���wO�6�U:ؾ�.;�H���B�Y+�]s;�nm�Y=��d䈱VRp�,�N��Ǆ�b��!�m��ӏ�K��U��k�~�exK�+(�]^��e�l[�5�+�}�nl3v���s�����/$�7�V�GW��EjA��;G���g���+g1y�S��C�@u�P���H�"�$	ó��g�tE�j�?u�m��a�������s~y�"Q�P�[���S�0R#����V�Z�����2A$:�P���PQT�٧�՗���h19��5�켷y�T�E"P5����>���ٱs
U�j��1!f:*2t:UR.��L<���-�7�w���i�j�s�1Gp�u�0i�p2i�����SNg��TF��'e�p�8�僈
%�&�|�LV�)M�7Q�@L�ݝ�ŉ?�Js�2N8�@n�}êi�.ΌN����/��U�Y�v5�D���6-��Z���� �� ��G�l��%�s�ΎY����J6&��N����T�>�9��U�t�"�}B��S��2e��<��#jt�S����_�Kn�RP�(&�~&�O�bRmN�n$�Y���fh�S�@�n���nl�mXOww7Gv����-]�)����#Ock{����\	}�p�_h����w>X��Υ����Ԯ��C��9��f�̘u%?o�f�}��Q��I�p;���b�O���7s��{)w��YR�D��	����T��(�}"�H�i�^�Ӕ���K�g�y�_x�v�K^���e������W=��r{¤[�R������JO>�R�e#�NY�ZDoX���E}nTN�K�*(��%F��}A1V�b������c��Q��	�S]����/?~۽��A#�C�<��u�sBE�&��ڡHAE���EFu�6���VB�^i�XG!�8L9k�ue��dC�88��C9�ģ�.�QuPg�|��g|��D-^���=i&mr�&B���k�4��n5�~�y˂�8�GqdcL1�s�<�";��i��n�b}XɄqc��"k�j�Z�|~09��-$�>N��jeB|r���++���Y�6C�$�>�p��ƭ�b�7�c@�����R�/������8�=w���l%dC��Q��%�juO�0�W�Q2hጕp:�M47��̦��G88��*t�pdB4�_��sn�琭C��Bلl�ļ�a�lvu[�;Mx]V�������>^L��ɴ�M$lc��l"�%�#�tbMEu�X�l1{�ʩG�A���A%�0��,)�2���&�W�-ᬙ�c.(�x�$\��h�Jb���|H�:43�l�9��2�Y��f�-�}����7�K��~����⫠d����?�)Ζ_�΅����T���cμ����KH
gE�?�`�b�)��L�ښ�8�Y��z��y��\~ѹx�6���;N9�\�V�n���9�d�Ă�ziݺ�����	�L$����:W�h�`vH�E�F�W�6ْ�C1�
����b��ϖq㗢`���c�b(�!.w�q�u�����ܻ�O���<��c?YS7'T8`gA�9\:��%�V�AM��w�xJ#pU��d�ج:Yb�T��8��>�pSwŃ�_�.�NR�XiD[���W܌�x0qa7ٵx��6�#��l� 0�P����	+P�-�ky��ٜ��Q8�	$�D6#iqvK޲1q�MFz{Rx�6�L}���,n��bR�R�ݠ���ȯ�1C0���o�����0�۱墤"}*�nom��(��'�)��Z:�PN<�DY�k����	�|��s0���'1�1٭��B�B"4n��3xl9ݍL�0�'�\N�����c
�◫D`a"إ޾R�(���������G�cЄ�1�6IJ�z��-x,+ު~'�X�q�:�׬`®c9���?n�q^'�7Xm&���%���l}�#��^��d���l�kT�d$�nU���d���p{\�0��o>�b����y���o���`g�$G�yo.9�,��k���jB{�����&���Ռ�Q��M�
n�n�* �i���f֌�5r�O��������P��Ǝ�nU��sQ����3O��{j��ӵ�$�>]KA�e5�3��2t��
�	���T�a���nu�,�s��d׎�^~��{w)7�1���?Yy��k���+��t(2�HA���荨�g���*[�H���ٌ    IDAT=���r���-�j���WaJQ]�uW^ʨ��,3e?mQV���ĀSg�C}GDgVAɍ�b�9���NA�r�%�@�l�$��[���s��Խ1���p��$^����9��B� ����_6�r�COa-D���Է���S�&Y9�`��kă=���iÓ�{�F�k�۩*-ՠ����9�	۞���@�a�"cCj����A����d�L�#��+-�xg���#.��^�s�O=@����E�5�1�n8�iG'�ᲡK��R���|~�o�0BY3&��XZ���x\��1g*�Â5&�0��R�a�`�>Lݗ}�ܓI��p��Sq�B����?�2�۩9���$fΆ�_���&E6h�`��Flf�rԭ��3�>��n�
�]���R���?Q�c���*�g��%+L[�Pn��i���G��}�4q��4mR�:M82��u�����(�����g��5����z:Q���b��)	��lk�n��n�T�K(-�����8�Fқ���+�/"��g�qy��wH�v�;1��l�_z�����Ŝ1F��B�-�D�dg����y/���{Y��A
ʮRP�+Ʉ�ZPLb	�"�[i�ɔ��v�O�C�qb�V4H���t���#rŅ3���1�g��O�+�$����O��ec=��a�$��&_~ -��(�-�l�jS��]�	Ρտ��tO��.
�&R���QlC�Z�|x^Rva�Z(�8�jj���~f{g��]���љ�NĮQ"N���X���M��pgL8�1��[V2��Õ���'R]^B.�% ��DZ�\&]��m�ӲV����՛Gvn����9gCBý崉EķŢx�����`NP �UR�5�W«�)�t����+%U1�ف��/e��/ɮN�\@\��L
��zIn��t��Y��+"�l�L��EEĺ[p��h��Jgs���w=RC��䰣g�]�e�%S�t4C'L&���AFd2����X���~��0��oO����?��=����t)�~8÷X`"�j��P��������'O�[¼D)kYզ�ʱ*0'���$Gy/�nn[�+/<�ӏ�W�'���B�'�!�O+ݥa�&H�u{�>�tJF�FO̤�Iu�W��ls��0��ߏ<��E���{�'J��<����7�h��[
�#�0�:^}����7u�!#�ܷ�?�����%�'�		-'��G����M��GbC�
K0�Q�1�8�e�yX�s�մ����QYR�i'͉����C���Ep��f�ޝ�>���k����6z6�X:IX�GDl������w"�y�[��y�NR {wA�#!�����JƔ%�c�ڙ0|�&؅s	�ʊiݸ����I��q�z�#ƒ�4ۈf�I��qr$�΢v�������Ɩ���g޳3�ܭ�t?�BUp^\&Ͱy{��D}RW�X���I"�]V����P})�ZL��KKo04�P7r�e���\K6D�-C�v�t<v���V��.��2z��X\��F{��,�3O#J��������e2V�?�\R�`�ۡ��WM�����Q�ⶈ��Y�5X��'t�#���r8(��t���nՀ���<����O�6���/1`�Dʆ%m�hO�l����I�i&˩r\���d"	X�eC,�t�^s�\x�j�TD(#�g��4�v��˹�ֻ>� �J���)G2�Qlے���dA.�ݔ�~�6UI�(Q3������ �Do/�LJY�R��.A�Tĝ/kq��pF7ro/���{��Q�ӓ�h�ىH�@?M�m�|�~�����w$�V���yu��{5ӑ�q�Y�pV򦅐�5[E�Й��x����{�UP�z����-T4p�~P����Ց�((.�dS
69�f]!:�I:wl#������r����۸Q�3���������о�i5߭�������������f�[1�־�n;7�� w�e�U_�A�d�L�L.���Ô�R�#��ZAe��1F*� Iq�6leӲ�9��ǒLĨ]��;��/�η�j��ο�6����H�E�b)�7�l5\�%JU��;nK�doo��(#(.�
eIF��o�NC[��~���[�;����H	������>.o�H�w�E���7�a�e�R�z	��?�͹Z�NZ2L�y	��y	�⚝lʄ�6q8��q5�(��l#ǜ5w� �*=�l�D*�I��G��ep�O��[[�m����&r�I�Q(SƯXT�C����xm�<���b�1/�[\/�lN}l�bQơP"KJ�l.-��z\E,3�U*��\�捿�۰*�p�X��0��e�5��+ꥧ�M]�%���,"���,H��N;D�RF)(N�5�U��ٱ}d�������@/�ti�4�p��yģ��bb��Tq���8D���U>�����X'�2�o��<�$/���)�<��RPD��DVƲy4~c���dh��8��b�ZG��e�+��}���?(�􎷗��m]��P�Z
�v(��6�JV�x��űd�ym�����P�Qޟ�<��Ǎ��g������Bi�>+����F����e&�� �Mړ���o\AYQ!�=�P�G�әTn���fPr��5&���.%�%C"SM���d�xK�
�*�7�B�O���(���?����/{�7?}��k.�ŅIW�:b&����D����D�d6Zuc��-�1,�"i�fBu��k���Ś�d�B�>l�%W0i�i���J����6���MG[3v��j*#�X;q��&�bN��g�9�%խa���.�M�*�{���~F�V@_8�]�Y�զ8~s/>� {��P�ξ�,�׷�����>�*�h�����P$���'�)i�ԝcۚ_R����O����P)2�K�$��mJ^%���y�Ͼ�������9�FM��G�����Di��s6�a�,�� ��0NS�ҳe9O��f_���CyCtE%��=D�=����sOSVbX]v���o%[XJ�� ,V���9���\D�a��P^���26�XA������sI������*���aw�'��u�؇f�,�J�գp�%�������Iڏ�F�ü���2��v���οtU����Z��72�-(F��N@V��ʢř�u�ڷ���c��;yPi�2��y�S�4���竚�_P�}��Ű�J��lK����M��T�<�8��s<~� Y"�}�*9%d���y�ݏ�e�:�;��$յ�ńka������n^|�n꛲\~����~ѩ[ec��I��I��d%�X̋m9
,�;�1�e��2y|�ް���/=pf�v{W�>���&"�-<r�}~�T�B��f���`+�"��j~��3ߊJy�䒆�0T�2��m[�K��X�1*�
�{�=�y����L8!���Z{����8Iì����N݋[�����|ʂ�?��z�E���,vY��/��M��z�����w�ߛP�$��C����%imm�l �5I���#ܛ'|H�B<����vV�&�Ȓs8)P��cbJe�w*K4��c"ӻK��w_z�1��x�X��s���@���F4>�~�=C�Ob���*�p�E�h���s�GW��'#�ӥo����h��j�$��g�<�o������|�3U#&��U��-C�k;�x�FTx�t��'�p�Mw0t�}��J\:;v�sB>>$�z�Q���b/>��`[3g�����NN�I&�D�$�pQP����L"�aZR�77�����H��Uફ6]��v*�&E�!4��_���~SP���V����q�vC0+����)�P��!#�ǔ숴����;�8�������)tK�_5V����Ps��w����_��71�������5�FR���p��Ml�k��W����AKw���IQy��|�XD/���aG�&�s-�]<�p
μ�N�fb&��x��\(�Yen4�z"�q���k��˹�ӹ��c��Fc|��W��eC�'�YX���[o���>��o�^��	�h�����a o��,���J��B6R�n�����M%)�������<A;�=��.��&����Ӯ��H(˖�&67����7ɤ���SPhf���9�$&p���h�N����^\�e�#�G�e3���տ߬�귫�2�[��b�7����mk�ԕ"ں�=��w�ч���^��7>��.�7�&���6JFD'�0��x\6�K����^}�^��g��f��߯d����X����*��o��u��,�rC�7�^|]�,^_%6�ǌ��Q\U��<�m'���q*�6`�жi�8���	�\���æ_L��I�~l�P�ilW�*F���|�S���t$�r�1��'q���IFU��[��'��Fl�ـ��E^b�.�{�1v�X.9gZ�c�fe��bd8-(�~�V��L��۬�������POz-��6���)�����oAٝ]��PPv�}�H
�F	[q����-Z'[�#��0����@-�M�|~�/���|U��z/��C�-�o�/�G˲������u�e�K^��T���|��7|��w�n���X�`�%q��*�:���l�����gｉ�L�u�����H
v o�vu���ÔN���SG�X҉>��$�K�b�KOq�$C������s��,�s�gp��R�5N�e+W0k�L��׿rđ�N[�v�i�<�X|U�e���LNh��S�P�˥CI'3xL9��6�6�bx��?��"��:/�Uf�4I�\59���5y��X�b9�~^�7�`�� �Oُa����C�2�ǲ�1[L��q��5��P^|�5;���x�ͅ��/���=����mJj�L��o�{ב��UN�y|����F�JCk7�;�L(6���5C5�L�X��R���������kT�v᏾�w��0��bJ*�hin��Ir�S�}������/���G�k�#ر����#�-U|�����I4�Q&qF@D��%E��՜}����,}Vn���<��ה�ލ�٥��c���XC�o��7�~������O�I�ŋ�|٪d-J���R:�x����Z<v~��\,���s8`�h��N�t\	�b��M	K�{N�Š'�M� t��>`�C��V:�>]7�0�M�QPd�Q2��@�]��߬�w����_֮D#GLObIt��
�t(�L��=��h�������u(׿����1)(#[P�]�!����Hk�cA���o����d�����3A,��0n�ø ����L�B@�R~��2� V��dRl�֦&�� ���>��]����uYb�3ֆ�vt ��%M��b����y/0i`�~M��|�ҥ-� �6�c�)�����28�Ŝ��*u;��[�KÞ����b$iW1����2[ V�X9��s�풭�����:2=�|�ޛ9M8�$:C)���s�
4YP�%+*�α����s���y��L����:�zБ�J����WJP�פs�~J���ě�1m� ^{l��$_y�3�y�e��O&�q���V��đ�h�YF���^��7�Sps���䋯���?���F{k���j$��Fi�`�E��a���&�~�Y<Yض��?�~)��a��&)��x��5_�)G�C��%i�����+oT��]L(���Y�XE��nNQ��b%x��������-�˵�!�)g\xM�""� ]1a�zu5+ĶBs�`�j.:�0n����p�9W�5ށ��d?�k<�<!5J�Ŏ�[��0��SJ���.���$CY��qZ�i&��{Lc��3�k�ij��;��̼�x���0���f�:�j��&D�-�����c����L~����;���U�#�n@��gc�/|��t��������店]��+y]��rDg$�)�R��xg�����Cb� f����y�9y�a��Ԣ��錄0Iʪ�a$U�^q#��$vB֮��r��EoWnS�B���o&�5�z���
���l���D�T�UH�]�����*��	���9^x�ç���5��^I0g�d�h�*֬\ʞc���]�T�$(���5L�<��P�Î?�����Bi�I�U���3y�ҭX�:~a�g��m�b���N��4�eyg�"^y{���U�(+��2Y�u�&��1�RM���3�ǎ����L���c�U��������buI�n\-1�n+=�63���R�egN8�b��2f�}I'%�4�5��ob�;/r���y��;���/�ْ��J�X)��۶)�&p8�8��Bo[�9>}�ixc�"����8���N�n�xC�֮��k�y/!�ʚ���r�Cw!av�r{Յ�e����\N�L�IKtЧa�Y�������d��p�r>�?�*�Ӆ��tJ����fn{o.D_�z&U�y����48�șt���+iQڀ-�VҚt(�t��m��&c�3^-5{�$�:E�i!���֍?c7%8�8��s�e�n��E��ʳ�D����B���,�j����6�w(��X�s�_1�Y�W�'#�����{G7�0�w(�b줕V��Au��X�Ա�:���}��{O���\��'���N]��)��hA1G#�:�5|[[2q�S%�i٧����L�<�����o6�`�==�M̔��d9�Tߦ�	y�j1v����f_u	W\~	��[8��٤|�1y�ԱC^b�d�CC�ǥAq"a��/��>k��?-⥇n��C�ӑ�o~�-�>��I�h�1d� ��G�;��﹉b��)�$��^ġ�_@��'�)&iu��"h�p2�-�e�$��fs
s,�;&մYS �J/��)�_3�	�n��)��b�ve�>}��3y����D�����\}�\�� �����۾Ӆ��3g�ZLtlZ�+�͟��c�g߯�����'��[HV�V�L�^��>�97_ϸQ�y�E��廵5�u�Fg"�؎u��;ܚ��qY)-q5s��	<v�,�,>��ގ�r$�-�ʬ5gS�Lq,�&�Dx�紓�m���G3|��HɃO�m:�G��:,11��ރ���l���|�B6r�!�p�_/P��9���g+k4n
!9��Nb�>�$-���S���>�h�18�Yl�d�A_V�W�X�(�H�����Zjp�m��SYRA��M6��v��q��s��39���t�e����8|�d3�����|5����J(f&����"��noRHd����q9r'C� ��{�W�kQ)��v3��� �md$7��Y���ZsZA�h{��O�7��?���>�lMo��Wٰ�XK<�%%�n��H�ܠRP<���~Ģ�o1aR.Z�����I�U�� ��y��7Nwc>�"��\ÖHS�v�W�~�!�������Ͼ����^����ehj4�$�]l܅���G�cY��g�q�,����n�f��jk��p�i3)�v_��0��to]�%���N�!�p4����c�"b��+����Ӭ9LyQƜ&e����:Y�z���y��q[�,]���7�E��=��J�O��m��(�P�n)�����2nwa���\�TK8#�g]��:p�̔z)����m'�JRRॳv���ɿ�V���c��+�W?�LXb8L|e�^ƌ��r�?�l9g]z�A#�NN�=��c~��+V떮���n�Ѳm�>|g�r�bO�4�۞�G��#v���:�t�ldp��ן}��vݝ_��s��g�<	g� �**h�hU���n��f�P�ۯ�q�*q��K�iڴ��؃'�J�����;��3ΤI������\.�ƕ�2���e�, %Y��|���*�(3;ɚ�Sf���D��̦-�I��L�s_J�ٴf]��Z��sN㈃��n��rZ4:�|�[���-�**���]\EcG��ɭ�|"0,D�����.ř/4��۶Ka�w~��/(�vF����|w"�f�,9�d���Ɨ�w4��;������W��I_)�]r]�_�F�kA�kA��0e�ɶ�9��C��a�Vں��m�5p)�<!F�Ⱆg�����(����:�N��7���<t�M�[��EW݀�r8qkq�(X��jpq����of&    IDAT�4�.�2i֍��)R=�Ʌ��z�t�o�մp�u�1t�>�����Έ�RL]�l_���.?��g��'��MQN�yު�d
��"��������)��0� P�%�J��Ku�������>������Ϡ��B(.�3�:��	��1u����y��|��
n���[��C�{�	IjbP�zH{q��JJȕҗ�iNP�����+��3���S�5l)��NIn]�P�����岰�:fϽ�5�vh���<� E�Ej;)�f��oo"��e�y�J���;� �~'?�X��� ��̙I�������;�I��p$�Ǐgk];�'O�j�ބ�.ʆ���J��c�=t�6!�Yf�G�_����"�Vǰ+�<��c�|�|����}�L���9�Ù崓����c��!Z|��x+]w+�c&�+1��:�4=��'R��3�n�zl�,����eG�eE�:�l�8��>
�V�K��j��/�ᣏ�a��Zzbi\�b�G'�p����)"���U�vYZ0���^d�+�^��������:'ߗ���w(���c�e�QX4L�5	~7�r�eu��Lt6����w������r9ӵ/z����U=������6��cc�%�3�,�v�-��^3E%��(|1�O1�w���Γ&��3HҜ8���й��C��Ԣ^�A��
��i����7+T7i�2�-9���Hގ�-z�y,1��nvl\��}�6_���h(������8�q6�]���FgWLר#w�]RC|.��LqՕ��?
ATwB�J����D��)��������aCm=�_t���+6u`u�JDT�SRh����@6�go��ۋ�~X����C��_<���O0�"#���4}���Q�6y�$f�)�v@q 8��O���ӎ��[���x	��5���s�X��L,[���w=ǆ�V
*��)I*n��#G��Ֆ�n
JJ�°��z�	ծc�U0���!	~��z
<�`O�B!�I�rѾl�i�Î#�Б'm�1b�n�r� �Hě=�57��'gׂ2���3��q����[o4L��u>7���������
?C��)�@�~��?�.jZz����RLĈJ��a��ȌIG������j� �v���?69��IB�.�}�M�]��;��Ta��+��+�7����`J�J'�_No2�h#����+֏������}A1 c4�%���TD*/��P@���⳦���o?u��{���r͋�\�*��2�)ׂ����H~�Q�U�)+E +@ԿNR\�n�:ۇ"Q�-&��֯�Qk�<Y��ϕ�bRg6�*d��J�T"N��G}\�+��U�t�0'ׂbTd)(<����f����E:��#9NO�&:�')��� @ye�x�FN�Ɏ�̅�-��!l�b��$�1iO��l������mc#BR�tJwΙ�)Y�Ȍfl�|���38N����\����x�L���T���M˹~�f�8���z9ǟp'M!�uQ6x&�G0Ys�z�D:���i#���8	���jg 9�-;h�[G���9���'QQXL4��֭���#|��>�r)���<��46���M_g�P�m�T����h�F��5����Ŏe?0m�`/zi<��]�SBl����Hg$��>�C����8k��'����#��U#(,*"�T�?�r���I�,�0H��ЁE��S�X�9W]0�3N>������(�e8h쌷���_��/�z�X�I��GbB-$Hω�JaֆYL��Vi�`��K����x�������ӡcssK#n�auHĭ�ln�P	'�E7��������)��YMj����p�NC���������J�����z���,��E�����Pi�{A��,�)(YZ3]��<���{�^����������̕ݮ�a��+�"b_�F.WO�L��"�)����E|:�������jn4K�8�0ZP���84����
�
GZn��u�
�Ihy�)J�߿�׹�$��8�2r�Z�x�iB�5���t�a�9�x"�ꍛy�yx�9.��|F��_�9QG�W_�����x�'hk�+'�5�I���RP�ҥ�SƣD���q��[�r��'q��S��i����>�w�E$"F���\��.8���:���>Z��3�Sg1i��e�ȱ��	]e
@���L(��l�L/�T��F�~�V�[�j����Oia!ɾ>wƏ��1�q�r]6��-B��q�bnkh&�%��]X@`p&�O-R�$.;��:�u�}�E�3LΆ�.�B#M$��� ��xJ�F�í����� _|��CF�ns-�t�Í������ڕ��L��Db�C	z�{)���fB�Z��eߑ����s���s/��P<NQ��P_�h2M��`���<�ڛ,Y���!��"Z���݅��t�ʥ�� m�mNSS����Bya!�Mu<��=�i�:���Q��ŖE�`w�K���*�q0]18���((��_������b�E+ʯ<-;������c���;�#M��c���`�J5:�+(�dw�����}��aU����r��^��7}U�]>��EFy�?PV�)���a��c2�f��O'��~�r�9��cIu}.�X�\.��qL>FN����?���e\�͇8yY0�I�|���͔���w��L�c���
$�>��b�����=y�������q�MljN�*B�b#)�Z} *U���G9�r�$�l�͍=�i�k��w^���Q;KaDwuǈ���5��@�.7��UG�m��̺�z"9�z�u�I��1RAmu�˚رy�nH�ƍ�]���Ѳm#�<���$�i}�1o����U�lX������3�8B��|��E�ɢ��r�C��GS6`4�t�����v�R �M����(�#��l��+Z6�Q�(����n̄	D����zz�؝."�� ����1aL�"L΀f oݼV]�e/@�#Td�q�
��t��a�%	u�Q�5q�Y'�����ߢ�;̄���,&��Jΰ�֮�Sa!��*,=��R�$��dp8]�o-cB�ӭ�[6.��ibPi9�P'g�z��?E�:u�ϙ�HIV�$���v�5n5��.,"l��蛟y�㯨�+!���J'.�])D�q�z*�x2��;]�7�Qz��}?e�����c��w4R���oʇ����C ����=������������C
ʕ�/�lm0}U���7J�X[�����(�/(�)�l(C�A1:��A<S/���D4��R($�!��]�'�7L�f��Z���k\�������F���CS.���bNG�����Ws�_&Ӵ���?��ȑÙ���312� O�氙��F-Q,�br���9��)>���G\@?�w��زV!m�9r�8����bv�Uz��H�fN9d
�wc�'����W-'�vy�,/6�Q����|��R�;�H�l�����8f����O���DӦ��4c����q��a�Z��JN=v������ٷ�Mow�r0��p�r�)�b�p�t�/��ഋoc؄���	Gu�+jfe%��x� <~9qM�;iٰ�]�f��!z|�b����>�E�%��bʔ=��5o��~��W��S1_����U�)�������b$Ƚ��Rş���v�4p�}�Vz��V��f_�������7Y�~5M�lkh��h ����V���.$�vѓN�;9�bL�Я�f31)2���Q6`˦;t(^�7l��y�x���Ē12$HK��ӏ)�S`��p��b�Q1r%�F�ܛ�����nMFAQ�ԝ�A�5��۰c�q����m�a�l]9��g$Ϩ��l������Dǎ����λ�SQ����_�ץ��ɫ���#:$@[��C���j�/����e��j(��/u�꯷�
΢����i��dF*k*�sx�,�ug3�$�EbÈF����E�Hm�lV��|N'���J�V�㥇g3�%]E������s�2��9���M	B�7�y�����+.=�3�<��M[(́G���x()���E��0�,�$/wV�-)��R�L"����R�2Ѳ�g��8w�s;�G��qPQ�#�I����lg��m|�t����mu�L�c_2k6�F5fu���Z@���룫�Q�G�*�>'��f�
�/S�0�tW]{������V>z���<��3��4��0lX���q��sox���m�b�hM0vt��&+���~�씕�)-/ n3�?x�r�"��o��˯���ie��r�u�*�U�V�<��7q�OS1j7�!��c^TEu�'�*]��r�
���/d:��V,���ƣs��, )��"C貵�<��k��POmC+��Jʪ�br��f3�ĔJ�˕�l�,ZQ�[\
��D6�KW[�X���3�Z?���0z�P�����_���#c�1h�@�*���s$�_��)��1��9����h��pF�qHFy�5HzN=%�:���CW#Y���{��ku�"U)("N5���o�S"ƕq�((����u��x-�`��a�#��y�TA���O/Yٓ��2RŁ�D���4�����qJ�+�i��%E�׸E�&��0��GU�(�Q��pIv�C�i�\��xG��(J�ڈ(#V����y���b禜�-���&�2�ɻ�f�_����dH�U�G��-��#�fؘq|��������8��k3f�ۗ��Cwr���ӕ�0��3I��1��HJ����RP�F�B)H^��
�	�����ׁ+�u�
�-�8=.mw�;�(F�B2$
���ɏ�,��3B:g爣O�K��U�ް�nY��5\�H����t���T:��¢"M(t���Oj����χ��YHq����=Ke�[�˻ﺟO}�����W�$��q�ߟg���5�X*��� �Q;=���))�(�UkO.�����niNr��q�F
�f���3(V'�X<��b֢"j�'�}�c�|��q��N��6+�d���m���8�6��"��l"	#�"��Ύ�+������s�m;]�dp����nX��׼��4�uS�����SPX�Nmm�>�bfp�$�m�P`͒��P�i^��%��hپ��x�]w�뢏�ᆛ��/��G�Ϯ�'���[�D"I[o/��A��>�����C�S�B�%nW8'�����]�k��J��|@����na'���a�t��e<w�,�9p�*�l��N
��,�l�7����S�c�5�~a�Ekz3W�x+-O8J��O�,n���zWԲ9==պO�;�pO�f�������OU=C��g�b�F�	�D��t*��"�����~�Wm"4�j:��}�`�Z�1�ҀS:�so$`M���ظv=��y��O>�,S�߅�~��QG��E^��^��3���믡���CO� s` Yw)�������:��I<Se�/����3x2!L�.f{� �h���z�ΞVz���\q�ETUU0`���$��_~������_ƚ[�p-��ac��$��g*����\&I�����h���޻�ੇn�e��k�q����<�Ѓ���Wja�b�����/�g�>|���6�聾<��|��ߋ�����ױ0�P}�i�Ci��x_+�}7_w�nv,��˯�M�7Ȟ��է�c�����������C((,`��N:�t*�M!����H�(���J�aOn�����q|$�I���u�F�/���c�q�I�0d`t�ƥW:�%d<]���%�.�o~d[K'ު!��j��p{�D�8�O���e��z�niTmOuQ�H/�x��'�������9�k>k�%K�����"_�1��Ŀ6��n᥷?����d踩�k%��H?�S6�yC$y ,y�|�~�{]���L�w�;���3�E�c�|&��%��u��e�%L��x����̝2���}�W.�3_��ǳ�������茥0Œd�=���4C�N�^4�i�V�|��g������5+�!���h�b�	CЬ'� �s���X�	����C:�ɻ?Z=]�����ȑ���&�h����ຫf�iy��R�PY(�w6}��yf�|+7Ͼ���������L��^�ҋ�s٬h鍳��N�h�x�/�e�$��R5��Mً2��[V�t��x9�7��تb�|�	�`t����JSK#�L�G�����i���GSp�O��8����a�2�6���CU�#xT&�}[���+�VQQ�n�
��;O�{3�t�'y�g���@%��y�\5]�1=}	ο�r:��,��9<�Η����?����1��-j]Y�u���Lws~[���u|��{��h�>�{�3����%�~��O��q��s���[8���0��%�/7��8�����������ŉĩ{m&r�0��f���f+�

4b��/�h��@ W.E��l߲s6Ο��ʱ����a����U�4}gD'�_X��O,���_c���WV�@����۔�cK�ؼz9~���Ճhi��M�\�y��6~�ѧ�~�Y5�`o_|�	���ᗟ~����i�	��Gg$�>>���qd�E�S&�RS0����QV���8o���&):�Չ��(,����	�M����c�t�FV���2���.��k������?��=w�3���}�q.���z�Kև���U:�;��*���N-(ҡ�G�zwgR�	����B�Jbʤ���'؈pOd[�c��b�,��jMn������y� �(T��A�g���+��p{�t�W2��8ƙ��瓏��N�i�k{.]�cO���7݆����AIf�g@e	�~Z�?_y�='���-Ɵ����jYO)�<P(EΈ�w�X#˟��n5�83��q݅gr����&`���̾�.�g/�u!W^z
��MN�J$�ö�,���w6��'����S� �*4*Dm���Q�]��C�(+��S��QՅ��
�m����v.��"�s�O?�h*�3/��/��\��"����J���<��{���Q�ۺX��A:�G6܍9�J�e���KƎ���ko��ʍ�����݌\�Z��^y�{�{D��v��;�0d�z�ߟ煅_1p�>4u����N���?wn��S�e7��4����WE� RE��+��tCH�PAD�=�@�I6���r���ܙ��?}_�|>�lvwv�ν��|��<�9'A�~���N�j��a$K״2��h���Z]�$�Z��Ԧ����L�`�-�kN������~;�3�y����x듇��'���f���M9SE���(O�#� ��]^��\}��mk����b	.��rl6!^_�"��ȃ�f�����k_>\hW,����/{}�@X�s�$;$�x%J�
�h��`��Pd����t#��k�6�<���C�"uit�U-_��sl2�o�Q?G@Y]AF���տ\��g�y�@�娫~w��Z�ۓ������LN��~P�Y��m�@̑X���̈��.B�>P��w��H�5	G�'�p]��cz3���'�)�����ud!�R��K�@@θ�A)Ob���!��$�:2���1>��^p�����%����n��9s������hó�<���N:���%yiE���1H�\Xm����J�A������ՀM��8��p��¯~�s�E�L�|�Xz�m0Sn���a�>h���5x��Ǳh���m߽DQ���>�s���DZ�S+�B�Pj4SM��&�St]sz�ўBP�F}|�s#�2�c�8�#a�)\��`Bh��z4^{s@\���k,��'��}����+�=1
u/@��{�H*Rd&�ǰ��Gq�-K��>;C��OƲ�W�h�]�Z��Ό�hO�ΉX�� &F�q�E�㠃?.�/7���:�B���X5L�H���j]h=J�E����:�{���ɤP�O
�����Uo"(O�1���$r�9�^8����u�=���P�(������1P��f��╣	̰U��$;p��u+_G����م��5��֫���9xs�[�ҡ_G��P��u�����9�t�n�|���*���Z���`��vF߂mE´�pY_4s�(@q��A!jP0����.�4"�f�Cql�*�%'qH6.D�T��9�ӂZ����{R7G&H��    IDAT� �2b��A�<��ڥW_p�3������^�bG_y�Q��w����L�
�̀��=j�:�X㱽ˏ�^��VB�^�g;��1%t�F]U�X<��މ�n�eΒ�edg��t�H�g4u4jw��\[�[�}|I�4n�6�^Co��\&���,2�G��$��ЎX�|Gu<�Z=���yp(���"�i���/�ʋO��?^y}�s�exs]I��L��T�a���0J�{*�R�� j|��n��,�nG�T��'|�GD!���܍�!7ә�\��/8��ez�Q�<����?�x$�]�Hӹ,�f��F�D�P���A�tϛ����p)��x�����(�7�~=�Ǽ�s$�����#��������{�����;�T�񙯝�u�ɞ~�a�0q��3�iܷѮ�X��S8���Ӿ'�W^��~�Y�{�q͵W ב���a���Dw�x��m)v�y'L4��/qկ��v��(f��k"W�EN�:v�jCk�E�� 3���.¬L�cl�8ӓ��S�����{<�l1�����Mi\�5x��Ǒ�=��5E�&+��B ݶ�����K��=3�y�s������}�Gq<6_�#�F�Q��q�=wb�X���q�)xꉿ�ƛ�����B��|��v��D9@�ʘ�LQ�uB��2��'�r&�Ӵ�u��EL�8�ϲF%ƨ
3Xa���V�m{�����S�6&�a@a��5�Rix�տ��s�7K��E��w������Rl����(C	=�к��8 �k��N�4hW�o����zXN'�Ťi�5#�W���R��U��~E7fk�>CQ���z�x
F�+�(�^������@?@T���6Smz�Vk%$�&:��Ж���ÌLF��w����o�D ��8"���~�����ŋ�^�d�F[���%]�lٖ�0��D�it�ǡ�,�l$�2�����݌�p�M��'?=���7M����R�&*8�c���r,��F���x�ɕ8��G��b!�ށ����殦��*�xk�X37�C���B����&p�e�b�̸@[,�ؽ%`yյ�་�D:���w��\�}qScu���:	y?#׎"�*NKu�;���R����A�0���Gf�֯�}�܇m����,����9������K�=�D2�gW��O�Ht,��0	_��W�nY҄*m]#�_Z��iT������G�&��w��v�ఃƢ�s0NLj�Ǚ�[����a<��K����#�=�l��6�`��4On����o�@2���3����c�Ugc�=v�d1���[x{
�}��ٳ��Ӄ�԰x�+S��I'��8L��mw> �އ25zb��N�#å��y��7OL�gkȜ\���, �N	޵(�2Ka����A3�iT�S�pl�L��̆l��:�0k ˔�P]s�mK��`����$���;��j�{�FnA����:���N�R��\�:�A����ǧ&׿�T�'��e������Ƿ|�v�N-gϚ�`��|�\�ƚ�+�^�<��+�^X���Ն�u���5<�'_w�P7��Ov���
pKi�j�M�6FE(9��hdΞ<��҉Һ����c�݀⺈l��ё!d;:�:@&�!6�t���ũ��H�4�2�%NsrB��V`�k!���e�4��0��o[�ޜ��]x~q�R$Sv������saj����8���?݈�o_
�����|CJ׬�ւ��*�P:���Y7"7d���Ь�`�M�B���ܷ0#����r�v<��#��۱x˭�f� �Ɨ�ͯ}Xʮ_��N��6$�����v� ��l�I��SN�c����q�m�cF�@.�C����	H�@|�mw�������M��������W�3_�:�o��k!�D'|���kNnG�N��boQGqt ��0wW���K0���tK���R����D	�=�4֬��+W�OO<�\�,df��&S��_�s�N�Mn*储���
bn�����w�p�'g��k��3f�E��[:{�b3��HE,���0��`�X�̡0r�pb�5�n���O���xL�]�@���E��-�+E1?4�v�e�nTі��n(���9~�+z\UH��t؞�QO�Z��{0��T��<	�+�i(�$�RqdՅמw�%;m�7Q@���7+���Ͷ4*�lv�����~V�ϰ�'׮|[������;p���Wx��������g{����z��/xA�Cf�mn�'��J��^8�&A��YR�m�j7�Q����9b��O� �d��$b^�F���RGat��H��y���ÿ���n�v�O�e��-h����l=�t+LXp�&K���?���"��H,��c���Zi��ۗ^��m���Q|�o�N����~p7�|�_~=����z��at�Y�p��h������C�8��>��q��r�ݚ���
k��1�͟/F�����`(!֮|�c�Z΋�*]9�=o���i�\�F���t Ɔ����B��]$�"���C�_i��7�Q�ېr`�ܙx����v��?=m4�n�c<;Ko�]x)�X�%��y\��*����Z�;\}����/�TM��gE�SgY�t�d�'����m�t[Tjx�ɇ����.;��(H:e@�����'�ƫ+V�;����5P�$z��b΢Ţ�FU:�U�Q�E(%��|��!N����uC���;#Kw�Ӹ�WKљNcx�0�t�7��[��tb΂Eh>֭Z�6��K.�)>q���^�|`�Ob�f;��b�^�֑L��jD�y�k��xf�Xfitx�T-MN%-}2c�S����4���>�/d��zT��6#�'rJ�=1�B�3Fq�\4-�z�E°�#�yj��-%_X��ۖ\z�]JyS�ȫ~�[u�y���X݆S,�69��� k�MS+W��ٌ�m����>�����������n��w�~���'��ǌ�����%s��I1�nxdD�}g�;R
ov���7$hT=&
n���#l���G��U+�5���������	P?>�T����x���YLK���K�$R撘"��f@!H˶�n
�<I�(����/��ހ-�����_a�� ��c�ʦ�U}�EW�_���8v�i>���g��|豕��Q�GG�\�2g/^��g�H��L�1�fHv���6C,�F	1��5O�Aڤ�s�a`j��\[�Œ��q�@�5�~� R��ں�dj�*v��V��X�&Z�D�@xi�3S�Y:����/
y�LV�Iv��=K$@�|c�(�m��b<��q�-�U��̹�����T��D�#�3o��s��YD�I�W��O�����M�x��7P.�008��_~Ͻ�2RVZ:!�25{t��f/�U?���b/�MR;+�9�K-��!X���\�9/=��})��ykxN��U�p�]w�e��\A<������ဏ�%Y˝3λw��:�t���̖�Td�:��P+�ᔋ�i���c�G���7w�v���{���f���s��TJ�����[#��=���o|��jN�x�P����8�>�X�b�A��$um<$��8L#DҊ���<{�UW/ٶG��)���^����W������t�}A�Ƽ��\���Fu$ՆS_���dj��?�������h��+��~�̸�ƻ>��[���?wq��$'P9�W�]��Ed�6�'G����%R�W�K��u�u��O�:�ZC
w�E��W��o��T:Cӱ�n���K��LIi-����P!N��U�h#K�VP��L�^n�0�i*X��S�����ڋ$�e~`L$^Ss|������D!?�%����?��hw<�p���C12�/@M$0{��p�0e�<����z	���Ge��H����vӒ�0[�i,ZE��h�ў!����U���$���<�0��o��.�T)S����Bte�.O�c�+/�S�͘%C}�nC��T����:d�)��!ҋ���U��n�:kf����$<�����*�B�������>�!�q�mX��?Iw0�щ�����[A�T�!�Z�F����63�E4��$�rf�T���(�P|�d6�Ǜ�_@oW7]{5fv&DT��j��A�ts
�s��q��%w��9� �j?%��RW��K�4���0��-����ꋯ͛=�o|��|��/.���?y�+��˻}�]�?���?��1�s.Z8]+��0����C��8"G<�F*�_�l2�~j�򳯹��v�w�&(G\~�ѫ���d�f�PШ��Z-�3 V�X[��o{�����]5��`�z���z�g�қ.��h�--_���(y��5�l�EW�؀�A*v�iHg(n�P`ۈ9F� �(X8.�������#�y�}p�W����9G�e��37����!�w�<�(��EQ�7�p�EQ�K���U��'�C���cutv%$h�u����T	���!�@N�q�͸��rZ��M	�Y=��ē��1�pwe@Q�i7\����{l��B�8�]$�I��e9$ב͠V-��'P�9��*Lga G��M�J֓1�r3:sp�(A)-�+j�T%)M�&���'���+�+�|~J0�	fW�"t#!t�T�MT��D$��%-�:;|�#2��V�|�zYg|?�=���=��qdr����0t]4Tׯ_���[7�j"���"��� q�T,D�,�BAĜs�ftw�aW�r��X�?W\tvX4K����A�9���U���~#���+̚�P���dV:�q�9�U�z ��]����^t�����6s�+H����F�~��Y>���A�_�q��:�������ko��M��ko�i�t�\3>��Y�\y�/��)f�(���q����I|�`u͛�;�k%vz��N�1�����ݷ?���>��8���ϻ��ͮ��7'�}� 7fu��lN�Vtc۶9���6�)[д%`�ϝV#RN���I
�:��Itv��7^E}z
�m�Es7ó�<�0�@fF�\��?	��u�ފ�`fQ��EWj�H�s�]z�֐�=x�	���u�'�V��mƦ�xc�[x~�k蟷 ��������W��%7b���a|�>1cҾ%�B��T�颔<��}��AI�$C��31�z���L� ,V�0Y4D,�$2E�[��2�4�%��vE�����%X2��%մ~Uc����3B�91v"�s�Ԫ��]!-R����%H||r�bI��	���)-y<�DRΚP"�e6xvm�xD��}��u8o�h�j�ʹ�̒�˶Ṏ���&PE���r�e	�K�6�a�Hr��\���zi��u��fɗ�L��[�Qƶ�1wf'��{7�������y�����[�X�vm�3�ʶ���$v�Ō�.L�� ��얥�26�ꉙ]�%��z�C����k�񯬯?<�z������>������w$2����]���C��B�Z�nX�윁D\CO6�rl튳n���[�TD����x�K�[K<������x��)�h�
:TFqJa��\X���}���������w�s�1������-;��d;��'RM�@"6����l�E����$u�pc҆!���ȗ���قy��P���2�_�X"	���D
�U4S�"ٚk=Z�Q^�eb��''іj�Bq(����4԰���5����OC�2H��0{��x��X����XV+.,�]3���U8ͧ��?5��3	T����I��3�dR4g� ���䯘�K�b��J�g���O��5��^d��$Yj�6d萟�$E����2�{2�54\��B#/�^�xҠ���%�Bd��uy�)S ���]:"\�|�_�F�K���Ys��-8��ҕ!$��<�e��JVI�!m�ā]-��TP,U�'3���-�fdkL�\��q�>G%b0�8��4S��D猥�.نW��j����s��3�Sl��%�@��u�>���B�F�=����MO�}Fzz�\vP��>3��GΡ)�Խ 1���d�f)�+��_�u��_n����u��c�ӌ����{���w��#����/v��08V���9]=݂�u��ߜX~ί�����z��1K>|EU�ᘞ�=�p��׊�JӮY�����?缣>��(���y�����'��j|���R���e��0qrmzŶ�'8+��#�ƹiMnH̳�MXZ�
�$���9��pjv	�Duj����Ő���uB7>�H�ϏNq4�1EyK�� �"��$%Սd}�*m��n]����g�1�+6�����Ky�!Gl�r���������ȶ�a�٨�u�S)��E��d4a漹�ݟ��R13av�Z�
 Q�U��)X�GÚr��x�0�PX��M�5i�ܲ�yneq��1:�1p��Z.	�ۯWОJJ��ҝ��i��-؋����]��R��-NO�85.�X#����[H��#��9KJM��|	=��R���������&�"���kH�-�V��bpe�T͗%Ȓ��HS.�@c�5ʂ,M�W�`rhPʒ��h��lf������q��0���FUfLqU��\��e���U9n	Z�R����
��4��#+���/����>}忺6����|�����?��vǝ>��������Fh��o��w&҉8f�'W��~��;��y
E�7A�r�5<��Bx�T�}V�s�e�q��09���_�#��c�玼'��_�Wֶ����50�?��33a���,l��7�����"��q�#@��+�Ci����C�rqg͙-R��a9��Wk���bܝ��j�$���#�K�*�����$�r:Ɏ<.�4Q�Mʃȋ%T<�=��Yfv�FG&߫�s�0U���̮$�t����֬���;�_0e��h���UC0�8��̒�Rv�QpAF����\�lpM��湑��f"|A�#ů��2���G�W�y�O�!����u���r�r�s-s�xrr��E�ae�0�������ׯ��� ںz`u� $޵E�Ѥ���ݿ֠eD/�n
���A�t�F��z�F�р�0�	�We�OD
�p�x)�'�Y������0�CL������5�����|б�<<��ZF�H �х��@-��)Nē
��M������C&n�:13hxa��zX�����}koo�������g���%Ǵu�����7��0]�B�'%{�X	$c���ၳo��7o�E?���y�G�V{_��D���]F{iz��Y�G?��W��G��s"��o=���,{c�슣-RSmp)�C�kY�-?X�=���h�h�D�Df)S���j$)
�g�	B.|>�-�dn%PU�;:$�8RckRsG���z�Ï��t�8��zԿU�+BP1�)�Ćc,�|�C*��]��+�F-?��կ#�M�J���KH���ud��ȶ��82J�$ �D��ڲ�D��^?.���^�)�Ը�8;ZA Jy4]�.�D7z�����#Tu�*���D/�"#��|��6#�R2ʚ�j� �9>�q�BJJ?�9�5m�Ȧ�H��&&096�d2�D�K2,�*��U��*j$:�N	�yu���u�����M*^]�W5iHP"�K����b]�y��%�$̸�x<.Cx~��m�"3�����D%E������2<,�_���H��z��؄"|�g�)s��C��pNh��y�J~Z�~w�g�;���O^�^���_�������n=o����\�~<��x�$�ő`y�W;�ι�+�n*E;���ye��ᔕ�Y`	�a֋�&_�{Aϱ}�_��������v���.����OODe�G��&~���B5� :�)$� ���056�Z�,�o�l�>�gM�9�S��J�X�wK$dD��l{���j<8~��S��<ߎ�d~D�̦�avc����J�+� �N���<�gg����)0��`4ɲ=�|��#�I�L'�{���kW�@�d
��ѼX�z5ʵ�,�l*-v��TRvu����D��1$-K4{xm�10��$y�@�d(����ɔ	����P(�ψ�p�g)�r|Z���J�}�$p    IDAT���*��x�p�3���o�V�S����n�">��O�f̊*v�5�'��7>��P�6<N,+�>�ש�ܨ��5^�dR���Od <��#%R�E31�d�tFD��
�F����1��i�҉)
(��.��J�ai��脧�%�%��I!�Gv6)��6��
7����ӉukW���g��܅�W�=}������	��:��?�苯wO�
�DF2ԸX��&̏���W,Qh�.��CQ����c^�r8e���yB��^��ز}�>�o}���,�݋�z��۟~�E����p8���PZ�c��eGVQj>��r^�*V�:�!?9&5�f���;KĒ�˰4�N��A�Q�@��Sl-�� gA���͜�G�((|}�Զ��*۟�j	�S�ׂ�Dz� m�Lj�k��v�٧�-d��fh�z:/&���h̢��G3��X+�����!�z.�e$C�4T�)�C�GY�A�'�%Qd;%"-2��<�C~���0���)�{�䄿��/����m���H��4"�=7�F#�L�o�s�Ү�'`�Ky���1����:~v���A�����Bg��-Ac.�Щ"EڬWGݱQ���� �n�Й������\�����m&�zK�J��P�!՞C��s[1"������-ݩt[;M�m��O�Ҍ<q,�E�:��Ď����0r	e�W���͗]���|�ag����/��>�z]��&H�SE�4���������y啛2�|��Ə&���"|x~mp�y~��gw��>����y������?>��K���:�%���5��9rɋN`�i��;]DX���Зa���D"��G�#�Y����I@�rH�%��f\nJ.>��|K�{n�ќ���&�qsC��F�g��,y�Py<<:Lp�1��0��e\t�	8d�}�����p�B�Vd��`K7@a�6�:���T�p��ȿAL)
4-e������"�.�h,\��H+ m|�xg�;z�,�f !�GZ���!�D/�&���ca��7����8d1+��,q��GD�����%��pb��?��C��6�/�	�b��nu�����KH�\(�Q���(�M��A%���L�`��	@�L���>b�R5���P$�HYM�~fqUEat
�̀�#����Rў�������}�C��A�E�%�~��E�zN������O�!�ޮ��O-X��7G��7\s��J�a�t��<{�U�+JK!�o��=�P�s�=G�<�<e��
위5��:���~h����P� =@¿��t�9��}W5݆�����[�`"2:���J'�P":j�S0��JBQ,L�R."���A��)s���}mr�rQJ�lG���4)�,H�Pg�^� l�n��e*TV'd�)��qJ!�D,I:RR�[��]G_��u+���g�?�C�OP,V�Բ7�nt\T�cz�Z�iX��&j�Q�U��mHx!�F����b����!��1���ni����XF����������wS1�Z��;"O�E�pj�O�����H�G��TŶ� �Cd@Ciۚ�V��^�k��<��~��V�Nƀ�L#��ڽ�0NY��)�s�=x��Wq�a���m>�z�#M�8gD܆S�1�8�A�>�P�u����F�D�J@3��*|�P�[![Њ]�{)TLi_��ٴ8�"(�S��$��STi���1#̌���p��]
5��C&t�w+�O��f'�v�5����r׽�����U�00����<�C�t�2�;��.|殫/�T%v���;�I��SV�o��'�ò��MO/�����?�?���|�ow��U7]�k��c4�&�\���Y����zְ��mӑM T�+��S�Q�(|��D*�\{�L�πR��D�Z�y�=͠~l��P8��1w19|tf�B������*��[�Dӳ)� �G2 99�L��uo=��/���>bu;]���/�_x���L2}�(���"M��_M�e�Zz�j�t\p���>h�oR����kA`�A�����u����!��6b�e�2�y�y����Zx!�C�V.��z�yRhV�9y�h-�ڬ��9C%Ezd���W�͚���5l@�m�ͯ�_����y�)|���`�v��J� 3�*��zg�á��L�}A�u7���0,C�C8���JNC=Ɉ���S�2�n�Ɵ�HP�Z��hL�MGbb��t�BL����)0g�"���%2<W}M26�Ζ�)�gb��Ȫ�����'ݺd��${���f��_x��﴾b#�'ST��w(̏^��]Wn���p���<�)�I�������y���躝fv�|�7�t��
������u�ϼ|^��)VV�Ι��uLј�F�Pt�������M�&ÒlV�@�,H��
���4�3D��qC��У]��0O��=�q<���6V�E�
��JP��/ ��`�f����(V�\f��/PL��*>�����p���a���:G���:J<�\.�BaZ���Ĥ��	.��t�11�˨NL��_��fҒ�)m%>%�D=��������73�0Iy~S���P2�)�I�D��Hq]�?ڬ����cƀ��]W,-���ݜ$;�^�l�kT��$���&��Q�"�c�U)5r�$�נ���7_�5W_��|����'�C��V;�"4"�.I��9u�qS�0�Vi�O<��h���ϐL'=Q-�{���T�Cq�p8��s ��4f]���	�3�LLQ7L>s*m1�Σ�lK7��4�7�V �P-!�ߘՙ9��{~�����a�sݍ�~j���O�X��`���`ɧ�|���c�>��+��$
?��v��2NOv�<a�����D~���W�<��_�����U���z������_��ɓe�k�ZГ��E��#>&�S->E�[�e�`�Q�*%!bڮ l��jN�[2����mH�&i��S48<6c�,����K�![г{g������t��1����W�'�rE���6�W��x.�*�|X����Wqީ��7>���:��v�~
V�̦�/���tP�1���c�bd�"?1!?'�;5?Q|��ȌS D�g���@"��fIؒ���7H���hB�{-�������~X�P��||o���,X*��6,Ӑ���8��f�Z�eۖ���1���z�\p�rء�M���/8���`���J �1r/p��΅�"bO"��%�U�I�4�wl�Z��������F�*�m�_�9�y�TZ�=|*
����1i�7K��=83%����!�>��#e{�"	Շ[���W׶��K�����͛��Ĳ����������o�;y���z�j�'�х�S�7��=���7(+��[�{���D�����'\?=������o�ԇ~����|O�xZ'�/Ϭ�wȗ�zaG���lX�@'kU��1[���2[�EZ��J��
�*R`�����h�H�$)�������7��Z�����u����XU%�gvsm��8�r��֭�7�̧19:�W^yEv5�/��d����̺�޾_G{B������N���i��`��E�S��ɶ)����꽽��Ά�t"زe@a�I����lv�d
;"��|E��#iIi�����a�L�[8C�;�������g�:�-���� X�"��R��+��HƔ�dex����~ыM[�~m�3�⒋�_�|B��_����f׽1]e��q�h�0���W����h���Ȝ9$��]��Z)@�C��
݊K�kd����2��2S� 3��	�s��d%l�a����I��ç���|��P��@Y�JMp�&��o&���Mw�r�9;���4��n�g�T�\rÝ�X3Q9��������d���N��Go����ˣ|��ێ{���`2��Wt��2��:r^f}�.����'}۞sr��t�y���9��}ϟ.Q�C#��fu_��"4��/�N@������sE�zU\����O	^�0e��HX)��U#����ժ�t�����GؑL�e���a���kXf�D\v�|����a���hT�agմ`�2��B��]�Zt�T���Z,��ؼ�/=�V�Ý?O�d0���,������K���F2�� N��/��xMG-���H˹Q~�.�YK�=�2��x�l���;%&�瑧5�V��T��a&�LPC��0i�y��J�`�u衃��\p��8����k=����羄���,TxJF��]��VRh���B��g�)�r�y��3�l�sfh�Q���I��JL�����4�S(ʰX�R"�N�C� �͜m��"\fJR
bu�Kj��Rmr�C?���?>��/������9o��s�ם�w�Ͼ�z(�k��-���Ž�Y��v�5�,�|�g�����p"���"�)t�v�1��C�ȩ'}�c�i���+k�<�������93�,8�l�Q�Tǚ�FbS*���/�V�$rիU4���y�;�}�.�h���q]xA-fSL�����i+l\�EqbBZ�qSGW{������p������4���`v/�+h
4����0���P��\㵗]���n��^h��,L)��ʐ�K��(���,��$Ca�@_�&�qObhir>��#��a$�o��/sl�UEYF+���?}D�O&r�###��-�F����+�T�G*i���aK6��eL��W��E���
���Ǟ�M��6�ph�J��fFʬ�à�G"O�!�R�uHuF�~��|~>��Pf'!�b�:ꅺpK�5�؄禔LBMDx���a����06��&���b�P�$|n��m��0 �16�npJ+z:R�<�����\��xy�˯�霊�}x8_3D�KL�s��.�I����|���H�\���m��%��֊�~�d����#����!�(�=�@�Jk4�p�����Ͼ��N���������q��'��W����{fo�Y��ilZ�qxb�-(�9n1:���юJ�ċ��ӯ"���
e�/����NO�6�l��Ԭ���� �����j����Tdw��$u�'�Cv],4�8�DZ��EC�Q�@�����&�펶xg��c�gsГmR��[��P����V�!�Q<�er�K60ۥQF",b��ld�$���:��o����أ ��n�e[`U3���@�q�իWK@!@��"����4�w�k��xD�EBC`$�:s)G�)!�����$�2T����ii��-�.n�iGs�S�AOgQ��0�6aC���O�	�P8@(����F���q�:����F�������)(�K<��He��Q^�i�q	ɓ/���PG
3����8HA~�ڕ��ẫO�ć�\�^���uM�v�����ۧLTܭ�ˎ�؊i�d��:�6�x䗗�����=(����G��'��;g1��\Jy`j�6A0�����:~}��_�������������ݼ�o~s�i���]�Δ�jh�5s�Y����ʯM�39�+;q���W��zL�9{�Z��X}���`OD|M艸0iPx�е�s�x�OKG�������ﺨ�*ѐ�i�Krٜne}ߙK��N�41�}�(��տ��G}C�,G�c�������ֿV0hOY�����w��6m�V�[��\P*2al�
E��o3���>
v[g���P��L�;r��a��\����ӡ� !��
d��x�$�H��2��{��J��©g�N!�5M�G�Peg�a�J=��d?�P���%�����X2�e�j�
��+�GO)v�X�	x�&�4A~4'G�6�4�l�j�V��u5�Z�,�����]
_k�SAB�0�N������;��__{�?��;k����~�}�����U�c�z'��d^��0P���Ve�������MP�~�o�^و�8��1{��C�4�L��C]��3k��>9���[-����9�׻/������]��ىy��{����{<��_k��~�f�b����~����u�G�^�h�� �cE�*QvAY�[4K�hg�$�x���+2��>�aH0�;^t�:�:��Mm���,�T2!�'���$b���1�ߩtZr(|�ߑ�똞F\��4�����T���Y�i�͝��@a�ej�8*�߷0�>����մ�sNBZ3���9P�xo~��6z^���2ϳQJ�Q�&)	�#����NnJ�9 �����fFI�D��K�Y]��x}������l��'VD�7_(��0�.BPt3��7��RqT��J�<<�\��t"j�*�RU&�Px�H���]Pt(�,��$���F��q�aNR6��yg�&OJ�75�q
%�AYj����G�r�!�����_�w�ǻ=���z/���/�?,_s����elf�0��N��\<��o���MPԯ\��cW��w�����T��xf�ݯ"Mɾ�n�02�&����3����?�r����W"���`�/O�:�gW-��++�~l��-�OJm�L�8���0RK#@����DP4�7V(�H�H&s�7	wL�z&͛Pnl7�(L[9ا�Q�L���yѣ�D<�K�����V��f��P�"����U�hh��L[.
w,K�r�\Qp�jObzli�!T��ɱ!ص2�z�rc��x[Z�2cPmN�����)6^��(+r�������-���Ll��F�56���w�͐�jrjBλ��H�ig�� �Z]�%B��;9��)���`�F�k�����'7�l?����fn3�l �Y��D��P��v#�yp��J�
"Ȃf���7�JXf��KK��=l��d)M�I���b<���@	ĭ� `l��E����$e�FRA:�!tkjG�G�>����ӓ���z�x���]u�V�=&_���iFqGWe��&w"aJ@��շ��)^��*�h���q#���k�*�����*�Hk��#��ڈ�.bve�V�^ۖμ���;߳�~{�[�p��NհM�s� 4��>1V�O�M%�x;y�}m��s��������>��\�Y�iz�Ȭ0q����]��E��Y�S����K�I(:!� dwo�41�p'&E�i��9V$��b�
N�� u4j�+��XVmm���bg�.��P��4�l�+2�C�Щc����s����w`bx޿�V�H���}��ߍє�M�l�����*YN���q@ia)�@�N��b��#�
��ͯ��I8Z�`����R酪��I��2��2􎑕�EY�p��j� ���I�S*7t��$aYɬ���H�\Tz�XT�FC���T�RFr���c�←b���A�u99,�s1�I ��;��d)@{G�F�r�� �A@%�I��5��Q)�2��H櫈U%��Qb#��~$�ZI�~�Zܒf�p�Z%O�UݫMU�f��.	���5���d�P������>w�g�u�WVl���at����w������{�f��A�Η�h�9Ś+���f\G֢�x�������7^���z蹿<aT˝0��zUj�{|���H�aO�*�x����b�]���G&���3:��ww��:����^|xd�oz����7T�nMK�ҝ]���*�<s��L��g��abyS7���d�)�ib���	(T\�Af{8ekG���Q�&���a�O�Z;
w�h!��/2��E!Q���d*2�E�i{���h%S��oP��ŋ�cn�<��? �a��Y(����ː�h<
���������Z�_�ш��c��QJ���j��B��v�Y�AW�"o��P����$6V-�������[�u��c$N��� �i`ɺ�4Q"� ���w��^����<���B�/�Le$�P\�?oaL�2��(z�F�3��H�y�5�s��L��Ff��T�#`[Xua�#i�8�
E� q����N�h"(�R�j���j%8|�aB�6���PZ]	&���T��o�EÂP����`�F�&�_���8������|a|���Y(C��G�u��W��ƪᏆZb��e��4#F8��U]Z�$fS&�
�ʨ�i�奷n��K�.�����15�5n�    IDAT;]�`������H��.K3�0�P�`�0ۣ�k۵R����74�u���[1�V;�o��f���D�ͤ��|����z�,Ės=gO<W8� ш��k�{�q�_i�I�"�Iڣ��gO8�����(�sQ���2�d�Y�䐝T(�!?:*A�ڷq�����`uB=������~�9�p$�H�Щ0<�����g���|Z�2��,:�hN�R\(bӶ$)%�f e��`�`N���꤃A1g��B}w8���V\x.䄴�Yԙ�^��F+�`"Q����}��&�Ͷ���q�ul��2e+$�Q�%�E�F�|�FU��x����N3��������N�DbԂ�p�sj�Q����5��B����zf�1Wh�b|��H��'��<̀Bk��a�4�iQ�ۨK@�PT�[Eè�.���p��Td�:5WDQl�ha�Jw�F�6R.V�����[/^��n���h�-�ɔ�fF)M�Ǧ�Xe�l���C�=�䓻���F�kaGW_W�XR�i3��z<���_A���gBͯ��Q�S�p��7��}���?��7��܊'`@Y; �đi�(/�et~�M��Rs(��3��қ�%	av���H0�ynɂ>AX^�wHXR���ftA�:�:<'R%��`L�Rp�2���ks2�F�/1�e(���$b�#Vk��YCR�y�n�NkH�������!=&f!��ȓ7���L�6
�P�j1��3N;�x|�+��{��N��x{�
��Ԟ�R�V��*5��NsaS��Y����)�	l6K�V9À�
PV� �
���,+!eJ���[�!Ï���u.[��*�Z�_cttT���.�)���
32{[�������Uy#a/��`��G6ۆ*3*ɅdSҁS���oQ�--e�2"��\پ9�����nN
���\�#l@��h3fJ@��5�Pd>ɲ�����&]�C�J��<k>3H򍚲�����EGٚ1�Fx�Pd����א�Zb�BשU*�J�T,۶�[�D�Q�k�j~�1��::ڳ�]3�1��؁�Sx����(�Ǻtw$�ST+i�3�����N+�i�|�-�,C��y7�8�掝Բ�S)z�����f5,���R�9v[ʥ�KI*\���OZ��yC1�Y�J �E��#��W�̝)�C*�;�Э�8ҙ�%B�܏zU�3���F!6�!Ő"e{�&�G�Xި�Br"����.^��;Qcc��Tq�'�)]��l���֫�ޫ�$�LN(��,�4ٮ"�x�i��a���#��7�]�V���_�@�{51.D>���i�@^���&�Z�|6e64�69��샋Pv{�4�H�L~�J
��X�H��.�9����7T�^�[�j��0����0��'����=�Ih�����cJ%,�?��j�I������l4�̊0nZ�?3�t:+�8����K�H�iTO/�M� %M���R��a��xʒ��V)��=���1E
3���&,�])l(��B@�3:�Q�h��:J�(�q��D�H@��k#&$GE�����)JXʕbdB�LR��3�Պdl��j5�J}M����@E�;q'`y�b���#���e�P�ʪ����_^�ix(χ�~����pDM5�fz�U��G}x��UP�^dҜ���E��'�v2B%��nF ߓ6�A�Q5]�5"�j���w�r�.�x��@Q�B��XL(G@�#�(hj��%ӡ�K.�!Y�$kI�C�b�ɑ�׎�	y�[%\PHrc��Dq�^f��"�2d
X�S/e�0�j�YI���[���h�Q��,�AƤ�#�q#C���s옩0uD�Kzr�9LON�L��p�|$](�#�:��a`�{��eG��p+�l�,)Z��G~E�0t��9>����D��Zx	���@>_ܰ�7�pb1UfvD�N]x"�5al�}����o��W"���j�r���A}<�GY@䯐?�C��	ɤ� �6[m�O�I�bɵ�W�����}���=X36-����b��P�*T詸41�TJe4J�P�	(dʶ
72��y1���Ӊ����"'��9����9�e����(�`4�-�Cn�$��{r5H���t��es�X�$�1H3�ӞE6H%��5�񍄁�t1��:�g���T���3ei�u����4����PӽSUmL'G�QX�d�v������� k�~��8G���g���?k|��ٍ�L|J�M��f7��j$6��4��� R�bN�(�Q/�";�l�����@B����	y�4��ӰZ��H�;�;��lF^\�ЍtE�"ex_>���HOt��^����z�G���:��vw�ҁh�m��͂�Vd@�^��>51&%�ϔW�E��j��j�컷|�l�|a����+\�~C ����J�"�#�r�Q�,�N��SS"�DY����̀djd�F|���Vf!�Z� ���q9i�`��n&Ƨ���a<�*Z��9l�h1>�����O��g����R������3�Ĭ�~�>^\����ʕo���/-{{�;V��kV�����=}}�u�=�vpP���r�	���5�+�#����`�ĩ�R�}�����P�T���,���U�0���a@��7�F9/�������f�+Sʄg[��9F�ؑH%"e��eJ4�-��l�"���9Z�I�&ט̴5��)z�JM>'���Ę@\k�S�� l�������6I@y+��w�ICZ��Z�w�b����
�ߖ� Ĳf@�	�vD�rglFi5F;I����Φ���G��n���7S��R�t�Pꥒ�ڸ�1��}��p��"�d55Q6gv"e����2*F��rL�x�Itl;�NH9��YE� Fbw�
Y�.��=�A-ZkR>�"�jP�GvdX/��+�����A:n`bd=��i����k�&��=���`|t[o�.\(��D�.����_����� }K����G�
N��8h��V[�P'�{{g��R�ԫx��e2�8s�Ly�U���c�I���h�]w�e�p�wb������l�2J�W�2�$��n;����J��/�ל;w.>���g���G�w��UV]��{�^�Lz5� J>ED��� "|����	
���bCAP$�$���;���?k������ʗ�>Lf�ι�{�����kϛ7O��m�݆_|QĀ�����ͷ���{�&����O�,� FM�!�h�� |����� �����;1m�]�������V�n��$��7�J��/�f�H'R(��roi
�5)�E��P
����HZ蔧�i��y���2nce�k��wR�)5�A�H
�b(�	L��e��iI�-�0DV@%6�U�G2!Rqi
�wH��;��
�0B�Wr�����_����(Wݲ�þ�s7V�]�l	�jɍ)K"�b1�<ؕ���ȇ��+w~]�oPXrW���j��#�cȂ*�1N����9RKG'rr|�*�hM���b.�bl�#���9�rTftd�y����dr���v��T���Y���-*�Ar3��a��h�@֟ ��PaI�e�����	d�vYq�i��{�B!���EY��x�P.��"������9��<o��p����3za��萾)�
��ۤ��A�_�^n<vE�L�$`���$�1�o�L���^yI���bՉU���'�����"�.�#F�XB�j���Bkk+R�4�y�u�l�u����3ϔ���������w�}�p,�<�&O�,?뭷jU'�U|�_���~�ӟ㤓O����VJ�l�f�gkVm@v��!؊VĆ��#a��OU�h����>Y�t������9�,�+�O���1d3)�P@�]�cҏ��z� ���իB�g�f�D��b�&Ls����U�;�UDd�+*6)(IL�$HJ��&��,�Vv�����{(���Oy6T��Koy������O'%P� �i=�����,E"�\�e�~��>Pj��)�k"�"�W�/��{��t+��{�3i)�zv4�w e��Ū2�2�o[���H/V]l�0q��\U֤m��s��9�l��$��!�"!�D1DR�:esEQ���d��&��S���0$qI$��bMB.;�C}��٧����܁U+W�x�^i�#pP�q�M7�o��,L~�,�j�<4>	U.t�N;��� ������\����t�R�\v�yg1�(0�y�������B&N�1�g���� V,�H�v�ĉ�������B�y0Riki������فe˖ᓕ+�v�Z<�� ]s��w�}q���@��f)x�ʕ��o�G ������k�\��G0gT3~\�{�9�t�	P�#b��݉L�OS+\����A8�n8�6$�cb����c�h��j��ƨZ���`����&W�˶,>3u%���c����D�"j1v��j�VR�?���_�݌�����7��ʪTg<6��=G(�Έ�X<�}.Ts�O��ݟ/��s�P��U߅7���h�묍Uo�[("�y� ��
�Q �|)�}1��Zdb� ��G=�e\�<�/a�ȇ�N%���v����:������hmE�jN���1�euB^@9�3���"�/�Th�,��g���^+ğBQ�!:���
�8k�M�]��1��p��T�	�Ry�UQ[��%�:s^z���89L)we����l�x�b��oJ��<E]7�!Qi&[�U�O��I̪���Z0�r�����cD�H���g�y<F��$����\ʱY����	�]%"��繜҄��D ���w��gH$����^R�ٳ�o�[ѩ|�s�)�}K�"�����< ���>s�����>�X4! ;oޕX�h��&���90`��`q�hSx�(Y�(�mlN��G@ɦ�ˣl!5�PO�`AEU	(6v�b7J}+P�`b�Z�z0�H���[KOƔ�JۢG	�(e���^+��v�D��ݦO����n��X���vӂ���xs4���^��9�+��^P|v�GC�����b�� �vAL�f�ҝ�
#��`�nkG� 7'ާ)���b��Q�)Ø$"� �� P�%b�,�Vs���"#+X^�Y��/��B�2���$�փvz����/�tGr��.Īsۜ��}N�,AgSR)�тw�x�`�ˢGqSo�'��^{
�x�bu	qjS�^i9T%LDj���E�A0�(I�(�)�3���d�֚���,]���3���^e9���{<?-���HH�2���
�Qc��'*M�2j�F"5����)�Yvvg	LnwM��(�`�d�i���?��K/��z�)�7^���q�,dջ"��	"�g�5 �рBPր��L]K9�����%_�%�DȔ�3B�\�$��O�Z�1�ӗ����([���&��[
_�1����<��K�s��'o����(�D��y�5��>[P ő���6��EnhP��74����x4��E��Eť%�sU�5@	��"͟3b`F��P84J�m�e��#E١\1���4Y�0���L�rEґ��F7�~�O�g�Q�̵Y��4��f(Ρ�A[�6M�4Znt4����G"%�
�)[��u�YB�2����H��k Q��1"&wu��u%_U�t���1�b�d6�sס����rT�Ŋ��MW{��#A��Fpm;�͊�}6��ô���̢���N���B�{�N�j����Ѻ��x�@ ;����7q�_�/�KL�4U��8��I��6� J��O�`0�%���D�V�H@��:�3�񪔧PJ��p(������eK���x�Ɵ��vu����4�0���"׶��?[9nG�V$��8�́6�"?<b�ݮ|��k����V×������q��قa�3��q(�P4�H�"!��4et�g��P_ȱ EĹUsR���,#�@s��0o;����D:B�:l(R�!�ȣ�P�9���;��w!3n=TH�R!oPi^�C<G20�`�!A��@�z��������X��,H��	(~�^'����uTD�F#�u�,�y�>�Qf6��ܹsP�}�]�^Ql��)����L0�"���X�Ҏ�a% � C�����B�m��M�JM����JfS�q�%�1Ը��&����72u RV7"'VDkDH�� ���Q
\��t6%��r@L�� �0�����MkS+�,� g�u6~��_���[��D�A���!���!d��-"Jb�~�TA�dIT�lvUz$
��²�6��WJ��eL�7�j�o��Hq��*cE(��"呢�Z96FT¡P�7��@&������e�ʺX��{�=�pj�5 ����PR���g�?����;fm���`����puNE!�D(4�fD�Г�hJNq����J�.�1ɡ� .1f�cU �ԅ�5��R':���P��+��ɫ�(�3w�6�V�*Vw�A���)JNj,l,%�W�S��Nda��T+�8j�����U��e��U@*.�����g�r��O�4���
.P�]��A�*����ԡ� �TQ�C�����hl��������Դde^�D4�,|�Q�b���L�Y D:����� c����F���Z�,�ρ*d�S��`H D+kYM��O�8��6�<�l��7�AG[�KE��"��	gK���{��*HDh_P��i7 �*�$���+�*��)O0 �PQ��x7%�'��<MR���� E�h�Чq(��.�
���[��u@a�c��rÉ�ρ|���f^�ĭ׎9�p���6.t>��e�?~G<8���X��c�t�6�<��z���
#SsP��I�R�F�S��E ��,�O����MI���8��������W�\,bؔ�ÆEDa6
�(rbJ㠋�>d�U	��D����kŢ��9�I��Hǆ�@^����X�|�p,$QE�Q(�Z��� A�E�����e��;�"!*񙄴r��͑t�J1�Bt�T��TF,�cr��KόT
��2���U5��YX�gD���D�Λ�����(:$w�1�Q_��E�l;�.dy}�Gc�V���P��C�"�4�N����~_������!Q$f�6��' ����*��Ooj$"�8,p����x�TN �[���H�RE���(U���%h�L�(��;ښQK̨�0��F@)����䫞��ߌ�L���l�P.��w�]_�l�u�BO�{y�zU��TO��a[^A�L���[�E�d���h���E2�*-�PX��)9.�"=]-6�Ph$̛���RQ*C�rj�-��j[�(旙Ȳ�#��*��$��$YBv��+����-=�=8*=b���WI�Je4�*�rd.��_z�Z��ȧ�(�R3d)e�ɲU9�z.*�앪IFt#$5I��R�6�	�Af����ԧ@ȩ�W�s��܊ԥ�!�o&��`dHv\���!Ĭ��נ��C΁@@�������R��X؟Ň���)S��ȱ���K?s}�]�2�>~%�Hc�?�ŋ��	'�$����	�R1բGM,���[�	9����>X�U�c	ia���}2���K��JN�P�+Gc��*�ٕr� ��=lq�P`׹�]�#}�c�����97��zZ��Q�1ꑊ�{S���3��</U6�����D!5�|��?}���P��\r��wE�����P<���T�(�QO]� h[u!ٿ36��ZZ�@)�ő����U�E<R)zK�?����8���?��X�Ot�/�%�a/3YvX}^�:\��"�K�ݪ�~����(ì�N9�l(����	�סR���"���Zʡ��I��＃pЋL>�$�eU�P�v�A�*Qu�h���C���r��M��=��mV�"��湳�7����X�ܐ2�S��3��o��L-�Kxy��W�T�%>���tVu�k�e4@��,?���ØX(�D1a��	��ꫯ��N����KY|��n�7r9��Л%��Ǐ,[9����a[��������nG2��GJ��&P(e�"��cu�(Z}���
(���ߎM�n�C1��P�)�H@�Ȉ
 �e    IDAT#X(�fL��'����N�3�P�C�ﱻ��]��� �P�2�p'���+)�ho�.�W�qY��(T�2|w�PI
o����鏑I.���g�����V��(-Y��ZPy9���ˆ�ˁ2�R�1(F�M�8���m���u�@��C{s��&��H$��vZd�Lk8��[t�v"����pa��
��4;:��I��(#*K�PD�k�3g�*���p���FA��UY!��";g#`")Z-j8ޫ��H@���������TK�T�dDJ�g�-��v�����Q�����[V>c�1�v_��cM�ntFϘ:/��2v�}7
�$r�dE7���&�6�~?��f�uZ��H4ō��e���������CP���1N��1��#�"�hZh���Ҙ��a�6��e���U��z1����Ŧ��,@R�ƴ���O�-�}�W���(��ؽ�`��V}~��XB�}'�֌Hy�P�b���Pt̀��F(Χq�`L%�k�($�D�OKU�|E�9���v��i���ClHЩ���'��aq;���m+�9P���`,(W2���2�=��m��G~mA}����,���?�ȃQ�U�{�w���/��ߋB� X��׋�r�HT@�,y�q��=�]�)�9B�M#���F}T%m.>�V�˴U�~�t.�R,p��{������� �Q�֋Aw�a��B^x�1��c�(���j��1����i���_��o��O?-�?�G�c,㱴(e�V$��V���Tnr�Nb]̝<���FB���<Lm�P4&r��r:!�6�$U����(3���"��h���(�|�玼[>˸� t�Sv���L�fb���ی����:U�������Ot(:B!���# !�b� ;���-y�
(Z�Ɣ���4)fؚI%U�!��q�,P�~�)J�)�$==ixcu!6u����^��lQÝ�P��j���@�2��I,��]��5a�}��7�=���ʿi�T-�W^�[o�-���+���ᜳΕ!�>?�f���2ա��f�o��T\�N4�uA�K�	�:Bi�P4���g�$�g8���:2��7�YJf��XmT����H�Fd��1�&����
OH�b^���$��/�UJ�����׾���6i2TQ�2���5��PZ&NE2��XBt(�1<4$�#ǐZ\��J�"zUq(Tʚ�JmU�ɘ(���@�K������՚1BMʎD���P�Ey�0�1Jrx����O�|� C@��Ǌ�>ӔgM��y��t�[�IٸPԧ\POtk c�P4�X?��)����V���vW[ �ղ�(���~%�L�f>�V��b/�*��QJ�Z�Y��>�R�N7{=��m�[�����|��yg��c�)��2����D7E���߰죏� �a�L׃c��#\��M��j-���B<�CD�B齖�7
�u�Cp'Y�ȡ�R��	�g����n�k�s�+z��p%̜9C���u$�19��"�� 2E��%��b��&@1Ƶ9@#R:�����zF��������1��x���#��ɔhiE����f� ��m(�KB��y-���ǥ���EP�� #�G�h�*<�qIF�N�%�#)[�yŲ��4F'�-��(�E�S<��l������rţ7]��v�K�z��a��>�G��:BQ���e4�>a}󌦔5�)]j����mz�JoF:)�m��@��zTJ��Ȍbs�Qs�2U�x�VD�dW�*hn�D�F��[(wpvr>v'"�_�J�E��s�?��8�ģ���яՆt<'���po��=������?��v�%��<p���ク��֖f��¨B9�B"..J
ۘ��ڠňq�*�^����t$����'�0B�8=�P�w�{�� e�	��bW���ͩ?�Q���f�Ұ�PİU�FFX��c�`�Z��֣Bo6-Μ9o��f�>J�%�*k+�N�dO[7�E �==�PL�%��f�Ɏv�G�w��hLR��;��D(f@qZ��S��an��ŭL�����9?vDa�fzn�x�l��OR���*�?���CIF�/�}���﫶'���q���U_(�+�]�)�E] ��|�(�E%�(|���65pZ�x�ec���fIy�C��D����U$����'Hg$<vx\4���R��\F�x��B���z!��.��S�졍k�ɉ3O�.��<L�<�.�9x�KH�GRx���?�T� �|�;�0i�cg|w;R����7U
e�b��� �"{�*+�aQ��FFmhLI<
�(�@"*cm �U)�9���¡P?"�х/r�+@���0̭U�X�+�Y;�JP%.{���^�����M�۴n���_S������&��hop�I'I*ȨE���sinjG2[��'�����K/���y�N�Y*�iI���W,ӤT<!�f�j�Q=e����L�	�K���8��Ai>,ˋ:���#�AG��(�N�z��0��9�2�VJYe_`�;�<�#5�a���늅���~)υ����Tp��!{8Id�]�����z`�`$줆n ��R�Q�X~$��#��#iZ�g�L��:����ɹ�a�a�n�:����&Y$�RP�Me�s�V�pY
�P����"	_YRm�쐔�Es�t��>D6b�e�ĉ���ԉ=�I��<Pq �,���{x��qDbi���dצ���  �1f^�b����}B�1"�:UΛ"ҌG�o�:�J�����gZ�Ҡ�ǌ��|� �����J�@��%��de�;[�Ϙo^~��	��� Ŵ�A�X���|L0������V>�c:��ԍ�ػ�~LQ�LӧO+�#�<R�ؐ����|��P3��{0~����,_�
��݋x���A,��Pk�� ��]d996,���Vr+��F�.'I�JE��N$��Pb
e���D�9�J}�X���a�~�"�2�.��b��6aV��1���U���n��HlX���v�b����Y���\������r�B�T�Ja����$��uh��ʖe�?��e��(�LZ�(%�uK)g�Iq ��(���ʈFE�As"�I�ߩ⢤�Z)a�iS� B%�����y_=���jk> �b	��������e+�+V0uǝ��edu,��A
�Z�.d����ݎW^�B
��@��� ����i@�S)XvOC�C a�,���HŅe�w�̵Y�!��rE��+dd�5�����Y��z���^$ua���($��D�nc��u@�6@���8]]�ӟ�$�l�dɝ�{�xk�E�c�ǤI���SO��w�������������w0�/(�����[��������B2���n�=���J�(��ɁjX��r�E&�b��)�O#gymؕ$-#V�[qP�&�bo������{'�C�ˎ�g���o�z��P.����pϜA{0��*�[������ȫ�E� ��@�,q�����͠.��F(l���'2Ѥ���!i��2,��N�K}I9�|&���\j�^p�8��1kg�]���xn�������;�-�����9a2BM�J�P��~���%`�5�K�P8��=���^�_��^�OhC�wz.FVV�Y6�_�9*����K�P|/hBm3F���cQ�E�Tt$D��Ze��i@�2i��u�9ˍ���\ԝȘcJ��CF�d�Zd��cD(��0e�4�GHj��)��i�T#;R���s��m���p�!���/��� .��W���~�+��_�P�b�tE6ǆ�X-�v�<`g0��x�2r|(�2����/�G�8N$0��޶ek)�ȣ��ǣ�@l��4@):�}��eE1:���=w�����n@٘�������M��C�D�{1������m��G
�^%�2�X?�e,@�j-I%GG(�` ebo*�<��TD�`K��!R �62ݑ�q.#fζb��~����Fp����˧|g�v��L��&���U����_��~�H4�7���%2����5�"��T4���.���!$��`+���s�9�����C9li.<F%�w���<��>e�o&�%K��F��q��j�ӑ��	�.o@jnJjv�Ẁ"c����� Tz_ke�� �;ѩ/S F$f͌��h�G�l�7�"%q#mc
��.;�/y�s,�{�=e��Nlr�"�:����o��'�|2v�q2���d��Y��,z���044,~'�m](�H*�6�#M�SE�Q�s�@��Fz���p0����J[���1H�� E���Fe�*�+B)����^E9Yz�.;]��]�P�r�C��&�C�By����;�m]����+�i���<��)�?H_
f2E��N��iQG�8;Ц��I3��<H��E���BA���6�^�r:��]?W\x����#[��7o �x�g/��E�`�oM&a����DQ$ ��J%DSa�Ȑmr=A��A�n��Z�]�ބ��kp�E�.%�u)SlC�ʊ����W�RjZca��<�OQג�a��ů�h�Sr~L��y(�O�2����A�x��B3�)@Q �g!�r�̧P>�^Q�"nu��u��g����xJ��9��^�<� �[��=n"����z7���E~s���ݭX�l�!?zz��/�+yh!^y�/ho_���螲�2t���f���T� �������_�j��=L<��Ѿ��#n�V%�܆�RS.78�Հe+��.�n�gS������G�����z�m9�m8m�F(g��������!�^9JY�P4)����
u(l�++%)9jMr쏱#
2�b���d
�|YJK�\�ł��+����4��0q<��P�%���~�v��g��c�<\��ѝ����7l��~	�~�+���r��3L{|�Q]ݾ02y5���H/Y��SUe�a����n�G�&�8��hk
��,�tXˆy�JY(+?�����矇ǫ�#���+djPTj��C���W2:� ���]2��T����ҩ�Z�u2V� �D�;�Bzi��m3H�SQ�A:�����=�p�%YK�P�l��/Uq��G[���ʟ
7�F�y���n\w�|}����� �ӦM�Tx�O���o�o6oU�x}���3彖P
�*�V�}g�	��+�̀b\����5��>�i��"����/{R��Ǯ�P��}{y�zÂ��]ӏ�W �U."�n�@�������"Z ��f,���Dů��|�үC@a�Q���ު;��4�Ly�v!_�T��.��f�hmMAx�N�ްJ̣�:�8\~��xȤ��{]X��/��:��ů������,$r��r6�Yj�W�Y![��Ux�lF�\�\m-��}��$�:ښ����qƩ�!:���)
������=���~'�}c��nB��X�T7��e�Rs^3w�jBWR�O2ƛJjQ���e����G�R��� >2�Q�Y-d#�h���!�3�L��#�L��������O<�3�8C�T��ɭPOb��Ej?s����9K?��ln�-�2�7oB&�N3����΁��Qs�-6���������^y6_:&NA�TVQ;��L9Q6���g/�y�:�f_Oy���v��J�s��������%ඡ������uŃ7]�3h����F(���3�-XX�~Lo�-�⩖�lވ��t٘�	������P�(�P���v���(>��PP�.��!7siF���&Y\�	jSdlh
�4��F��~{��`��&�*�x�ݕ���k�ޒO0~�L��ǣ/��ß�xT��$�����vPu��|���yX���e�h��j�24�|ؼ3�Lƺ5k�3��4&��ћ�ۗ���Thd�� EG zG7��Z�Z�20 Eƥ�@��Hc�vG�s����ٕ;���:��ī"_�r�8�).ik�2:`�s���"�2��׌�8O��!���P�z�`}�2E�����<
����N#�N�f)�����k_�*��cW)|.$SU�䧿����kף��-]��U�A7U��4�8\p��[�ț�:�h(���,[#e�n@��@.һd΁�\�� %^m>������4gs��g
�[��U�Qؼ	�.�FU�K�xm��(�c!`�����A���E�XK�t���c���jAS[+�T�:\D����"Z:Z$���Rho
a�������C���/��%45y�Md��U��p��O��/�ٲ=3�+[�+(��n)�|�JVz�PO��״��oX	�*�/%��v���erA���9��O�H��脑	��$bi��5�^�T}���5�J`S%gr.J_�t@{��\�Cq(
���k��.�.��Z���I���{��S�O�nq2|͈��w2E�Ԯ/� 56�
�~�:���P�ȟ�fp������q� 簡9R�hmn[:�y8���l.5w9�f���B"��n��'�/�2{�#�{���1س�=��~C�(v�a�����a����O�I�����4I�+1�����{��h��5���|�H��颞��v�)��e٘�Q�l\q[�C!)[ID���nW>x���'Ba����|�f���
Es9�Ȫ�QؼM��Y
E;�(,�q'�HE�����|�ll��@��@<�D�ǇB6�xd n�--!~����߰Û�a����ߺX��_)!��#��˯⾅O`��~L�u R%;
U���H�O��LMT?�p,���T�4���^-������\V82�R�`_�:b6N��)8���q:$���2��=*twg�G{���Hݑ�,?<wj�ϕ�+.t>��"7M��J.�8kXt&���6:�����)�����02�1�0��n�^�>�����.7S��ѭ*j�W7F`�=���c(.�*��N�/'h����-h?	��"�:8��/D?χ�c�ى���"�bAK&���q����N�����݉�����ş_yN��Ŋ��%�Φ6�2��Ƙ�{BG�25��K6F(��P�BU,�8��tC�HF(f@9r_
۶�RvE����>T�q�Ʋ+H�p��l���#�7ݡFPԂٲ�#&��oA@�G$b��HBR
�8߶PD&6�J>��ρ֖ ����._�;o��.9�Xn�v0��;��]�.��m\�v8���t"��	�ȩq�Ϯ&	�o-@(Rg�b�CA�!T��nl(!1< �g.���bp衇���/����&A���EG!�h��1<Z�D/<��� .=��˭
��?f��Bx2����e�z}(U]cR'H/��b<��x��7����̤� V����)��(��

�<9?ݔh�r���<V*����g[�>'q'+���P7v�k?����W��j�t�dB"�03�dG�IZ��)���_��~�K���T���?��p�}����z�-Ya���jC�lE�`��TW*�h���"�N��J���D(��,lP����$#�׬+�u;��о�ܛ���6u�Ʋ+@�]-`x�'(�nD�^�E���G��5�6]��N(
Yk��ec(�P�HD�Pt��f��f/���c��SL�����FL�Ѕ��+��}���gg��������-��o����@*N�i�Az�����|� A���P����4�Q��V%�[�T��	y�t�r>�K�&O�$��c�
�\݊��b͘Ɉ�'�x�w�q]�)�#�[.���������X#�6̭	(|�<�t2�}���FI����ߢ\�x��>��˨�� ���h0�)b��Hy���HNOԷ���m�TtJǟ1Bb� ���+��t�
�ۏ}8����T�<��]HRf�����#�ʈn�M~��0��"��he0}�T|�;���#ǪU�Ș�Y��7�x߻�6|��zL������-艞     IDATȊr�ީ��_">�@��(�5JY�UĢ������Pο�w�'��Pr8��Y�!�v� J�C�@Q�j��h`�@6�w��%N�)o�Pt�c��*�,Ǣ�@�����f��N�cCpU�l�y7�N���1sZ��9��I<���y��9ñ4*V��An랈�,��T8�P"��FET��0�B�2�*BVrj��p����3�@�EM0��d�-ô�+:L�s@vS~_>� (5��.���C���͌|�������f�k��E ��8Q���H������y<&�)��9�@�/������jɬ�;HD[��;�D&$��<�����kTUQ���(��kW���r8��Ӱ��e�f�篡�M��3�뽾�XTl޼	n��*��w�L�Ѓ�q.>� ��>�c�Y�c`��w�����c�A�a �E�Je�C��<����uI�q��=����J�X\|otg)�'�0�����ş�g�+�|��c^�mZ����%�j�����\�g#�-a@�P_�P*p0($��L�d,����ְ�����&���X��8d��q�K��~{
L��-��=����׈�Ҩz�����Ke������LD�%C�S`Ň�������iX�{9[%��d�CI&�gV�Y�K���%���n��КS���s��$؈Q�(�I=%P�w���f�bg
%�L�lcS�?�=��&���?z���}�H��Z�#	~�D*���k�S&����E)��T��C�F���O$<�\��(�)�W���<	DڱM�޳���DG{�m� Q�N�81u%���/����#��*ǘ(��X%�L�҃�W|��8T�[�����ˮ���� _ �6gP��:�Ӡ�A�1��O �1�����P�P"�)ϟ��\yۓwǃ�s7��|�*J����(�mB�HXT��f@�O8�%3B!G�J�$�̀����֌l���U��V,���,<t6�i�������������.�N��CQi.,g�2|�7G�6�� �Ȁ��UW�Mb$[��&��a�P*���\R!�SD�8�##���$���鹳�pM�S52V�n:rPтJ3̏$�a(#-^�����r\��L	Xvf/�p'Z�b�ʰ����}AĆ�5@1���(�YUq �5!��3�
hIҖ�SHT��@x.lT�48/G����涂�nr�b+�kv�<5�qĉ�"Cr(b(9&F6�γd��t��y��aE��RD6���(�<���=�+���K�ۘB:_0���/��&z�)���
����ߓ|�[1k� �-�Y:����P*6u��)#J�ɡ��T����ߞW<tӼ�(������~򞸷s�(��k$�!��[Dd�ҥ�&����1$�sb<�ܵ�]�}��2��SD2:�|L�6tu���R�!��{1}B7~��C�<��L��7Eq�7���^������`w"Y6za�ED������hmo�d6'a��J�����qH�V�5P)����J�#-�b*���vc8���7ހ����PPd+u-G=��?c���|�"r�)�]�Ӆ�kV�!wr���C^��C���,x#�7�D f��!<�Fƃ�&�LGN��
�v�j�δ+��k��f29L�<�@���Wi�c����i�X��^"=���_a$�xU��F#�~X�Y��.������G*��r`w�$�ȳO�j�?Єh$&v��4!����GK?�I'����r�cL�9Ms�p*b�*�0�n��d�8�P)-Fܣ�$�I	���g�@ё�����	(N�E�*����#��c�v
۾x�}�ۦ;`	�����"�"�y=\Y�����ޤ���#��ы<&)�2M�����+�b$٤GG6J!�B*:��׃�fN���E���_:�_v�Fg�R���_|?����� �QQ��ba�A�r�Υ
�Uʒ&�V5�Ǣsb%����p�Ω�������(�\-�`�z
ch�Nt�T���)'�u��	O�s��@Ue�0���{rW'@�k9��Čis�F\x�hn�s��Q�
Hho��Р{�w��n��rn�n�ӦI�C������ѫ�b*(���Dx��L>o@^��c���n�����I�Çr�S�L0��M�V�z� O�<�w�Q����R�*pҡ2���D6/��tl�da��%��(���E���1 ��e	6´�1ﲋ���;a���'h���o�X��p�[�>n*vD��-��{�^�k���(kG��8��\^�y�666r)F�A:��X������%M�,h	�QIF����+��s;y�*@y��r��c-?�ƞb���߼Q ���mC�f��k��P���;2�DG)F�X����Iw
���9m�q�h6�#��q.�����"X"�?��op˭w"����o{�X*��%�)1�L�*4�͂pK3�y��qH%�R.I���
xi��K�ܢ�*�X���b�(�ɴ�Gd~1��U�<[�M��xm�7�! ��#��A�������>}2V�X�fN�_CZJ�$%yT��S'�e�F�|&N_�"�ѡ�JY�_#kMD�L���^O�9�e�� �S�4w.3�ڰr�*<��#�7�E�	P������<G(f�S�[��
B��:�r*��r��T�]�I�+��QIK�3�L�������xL8)���%ｃ��|g��q�Is����s���xb�3���G�v�h���mK��G@�M�A�:��T�3;����X�@m�b��P�m����4q�Cr���fN���{o�>��7V�-�^���J��c�@q�s��_�B�����l"ßVB7uA$d��W�ymHģh	z�\
�J�Rk?^�I��x���p���Z�7׆Mq,x�1,z�ghj�D{W6�!�L�!NKG�^����
r�1�N&������%%c���)�3p���R>+�U3�dV�j��IL���ȃ:�|�a�y�����|S&��ԛ����ϖݗ�����ɓ'$�"k����jQ� ֬Y�5���.NH.:r5��*/� �{g/�N�x��7�A�8�ߓs�	Eu<�3����%�����x��G}�E����;�,�Ђ�����{�r��?-׾6���-�|!b��oEc�t
_�k$��r>�/�#�����1B�∤-�b�-kpX=v��#��m7߄/��%,_����#��W�{虱�pb��0��v�<�0@ TC�p�(��c�b�-���^�js�ֽl8���{�(�Bq�69�N�A��e��L��޺}��W�-�λ��R��㇬���P(:B�R�g�<f�}m{l�����G�!�Uh(��5w@��?�n��aMG�[�v��;�v�y��(�?�~{1�}�q��7/a�#��'�H#��@�	�]b�C`�"���f���K�q��d�2��ϯ���r	�|F�_�[����8�VOa�Q���A�B	��u�gs��$�&_�s..ZG��0a�\Z�Q�MzZ�ŝ�������3�֭Ú5����f;+1F�cܨ���*i�Jc4��!QAUq>�y:5�k�\%Z�C���1h���8\�,cww�ǜc�����~�3�A� ��_�r�T���k^;�n��4G�:%��QB:5!q����s����s2#R��"��(T,Bܒ��,&6�P������d<�ӎ#�8W^�-4�X��c��~x�����~�p&M�zc�,��2?�d''�]v���1B�|F��E��m��������o�J�z���5CR��\(Lyx��N�F���N�:��v[r(��x�8��e[x�M�N��L��B���{�d"�������F�^E�j�G+���3����$��;,/�I1&��G"�E���!FüiU�MVL��^����n�]����UF4���#��F��ߦZ-�P̋�c
lL���R�X�����՞\L�p��>oz.<F#.0�}&�������.���];&	;q�"�0]#KP�s�:*Q��^��*ߪ���0��1��S�_S��	��	�R*�Y͕�D�|x>}�����-����c�����c�" ��ǅ�Oazǿ#ϴj�F}]5��{P�܏F�̩��ɣ���y�o�B���Uh!A3g��BN����ln�P,�L6/`@]�����ɓq�-�Ì)��y`5&Ϙ���(���K�jC��SP���+�UD�b.-
_�AJ""�Z�7�M�y����7n�F	����]��x��v 5�lω�W>������y�3�e�K��VT����0B�\��q����3�z 3���9����r���\\ɖ	�.��/���objG�.��r�	R�-9\x�%������?Fs[,N/l.�Lx#�E��J%d��r&�T6��S�VM�i�Z2�l"��` _?�|�������<ˑ|�2f�>�T�Z(�r��P�TV>��B����S7�im�X?�mWG����k���<�� \T�s�1��`�<Ӛu���P������*�6��=ҎmFM
�w}m�+�3A��5�^m�*R���bA�~�B{��$�r��{�W�&S�n�AΗ�z���h*E�hW��� �c��s�*#f�E�U*�Ӝ���x��Z�~�H;���]N� �.�� lvz�LŞ�퇕�V��w����=^p|W�8�rW~�3{&�����}.�'v�q�*v�z�7�j]�'�B�hE�]�l�`�Q�$��g�e\OsJ���"�R��z������]�[3��Ml��هo�>�����w�}�v �x	(��a_�i����]��Pig�l	&u,���IW�\���f��v�n)�{���1��q���0k�)�s��]x�ݏp�ס ����˃t����$3I�9¢ʙ<TK�7 �͉xl �M.X�)�bQ|��/⫧�H\�?���ܔ�����,��"KE�L�Ŧ�s���h�wl�� 8��v%Qc|gQ	�t�Ν����2v�uךD��Y �$��֚��9�tA���N�"P�O_�F@��Z9+� ]�JUi��fH�ݍ�W�I�9�F@W39v��?%�c�r��b�wG4�������t�wȿ�L�"�2
�t���g�KFޣ���YLI-�ڵⵯ������Q#7M��?�Z,Ș�]ٝ��Rj��q���`S� ���C,^��bM-���|�+�E��9q��Wc睧�\a���߹�6���?1n�Lx�a�[�^>�:ћ�P�w���NM���#�z�B]��Q5]���p�9{����^��L|���[�?����iX��o��s4�ߍ��O�ն3��w�e��ㆬ�)��P4���_�-�D���T+\F�]���� x�%����,��MN�x����R|킫1�*a����F%��F�s\72��T:�n7�Ʉ��� �y�:@SЃD|^=v�1�>X�g~�����45K� �����ZTQ4R�L6���`˔>����~���Lxcsap'R
S.��j�*+;��|�v��������ߑ��"����k3t$�747J"�*5S #R2��B�:���M�N�S�*}3j�& ��2�c��X��!`\�w�ys�4�]s�58���qꩧʡ��ү�寧�鬥f��,�9 �5�V�:%@a��xl�7E@�n��k���*�s�{֭��ӉC���G�@<��tn�_&��͈�"����n�
'͝�+V`B�x�-���������;��p�H�G���$� �cl����/_w�B{�.��U<n
I���OP쇏�iF�B٢ʥ"}6�S=B{<���5�/��W����!�~{{����/~������}>�RvЁ_��n��AD�����(V
���pz���n�0�MJ�y�i�XRL�� ���}���o_�R!���Z��w����Dks���x�p�I���)y:Ǡ�Pm#�ׄ��69�P�)�j-��I�N���E0T�z!���5t�§�N�J�TT�\�t$�����o.z�=5� `c͡��u+:��z�1k�Q�Y��t��4-�'��
�GE(�G~򓧱~�F\����J�u@:��͑���{s�W�T��n�c�p�bQR]u��b�Et�Y�^.�:�k�L��\�y׹��e�I���7⮻������� ��Im.Q?�oZ�J>���{��9o��:v�mw��a|��_�����쉍����K�Ų���1�1>#�M�M�M���"��犊g����P�bNyX���촔�.e����r�v�P��s�w�}�>q����^7IYN^�1�C(v����Z�^���g�(u���(��ͥ)�i��1ܻ!6�X�f�;n�N��z��O����!�� ڻvҋ���M(T�?(�{\�����L®R��s\lUT��,U�|�\|�[��'+V��/����eU1�pJׯ2ufc`�Ȗ|J,+ҔE�N�P�^��3����ٹ#��եM��%��A����0�6��P���@	�T�SoH#��IV�T'��s�^�9��*���S�S���O���WTP�8T�HW���]� �?�'x����9�\���Ke���I=��U����|�x\I�"1I�tň���$-CQ���Z�c(�;�׏��v��@t����c8�p�����hk�´37ap(��C1d�@��0Z�aD{7�K���}f�>��6��so�r%���K�nS�qH��xH�<���sFO{��ʪ�SE�u@�)�X�Tb$)�(�]��$e��Ȓv�rŢ7n�ɁKS�ί^s�{�.���e�#�����B�s�"�B�Dy��[�Qѧ�m�@�@�"�N��^-cRW+���U�9t_<��]2�M�G\n|�p���s�L�Zz�+�O2�a(��Uu�6��Ĝ�N�v^�bi�J��v�%�8Gnȧ����D�2u�D�۰MM!�SI�as�xz�8M��9�(��,h'�8.]Fy��w.n����&(0��^Ե�@]���k�Q�rN��zD�z`�4+\E�͔J��k��R�J���2s3�w*���L##S�[Q��cƌR�"�J�%�2� Q�_�L��Tjd�A��U#>H��x)��0b�{~؞��4.)�:��T�:lbS��C��D>�O�����Ս��iY����hӠt�w4w�̕�+?Aϸ\v��8����i�:���M���o~�7E�3u�Gb��%��učA>]����>����*alY��ƬI٪�+���l|������[�zՔT���gʡPκ���;7h�{4�0�AdP EG(Ly�@i$m)ofM�&D\��>7V}�.�8pO,��f�(��hji�o_z_9�����#�6ْ]|d�G��%Qʧ��ũ����ۑND�q�)'��ӿ�b.��W^��_z�'MB�;S���%�P��8�.v�A_~�45��K�|��9ߑ�`9�%].>4hs����j��ݽ��:�g��m���"�g���V����������o��##�z+���t\7@��H�#�������4K�ʋ��y!]��E�g}l��N_���})���*�I �SM��A����oQ%5����b��-[�˴��S'# :4��f	�����U��`c�n�톳��~�ҫx�������D�����a�f����Á�+fP|$V�ė����"Z�����"�.w�x1 �fjp�5��[��\��l��kRV��m���'6�]|���.��v�e�jח��s��g�c�s@��ad�B@ɦbh	x9B��,��qm���1�;�M�z�b����%�D*WE���E�V�Ot�LE���#~����"n�-|�E�c��q��~�EO�@B������J�{h��"mvd)p���H-�R��AY��@0������&7����5�,���W 5�<#8
ZK@S��/2z�tʤ�'Q��Ob����Pt�S㍌� ]�֩PlT�nn�?7G��9:Z���j�R5    IDAT|�X��1����֌��|-�uR��U8*F?�HdP�ͯP��(��K�b2.�M��u�������f9��?�H@�T(���I�7�ɋ��ع'"��c��^l����!Bͨ��m������G�>������R|�ƛ�vS?&N�41�p8�C�EOVťl(���X1Mj ����R�[��؅�L���ण�l��s�Ly<��;s�3��6@���R��g/#=�M�*��'Oa��&������/���n�>b�BM��!������a��\{H��*�XKЇr.%sqZ��=�X̘6	�=�0^�54���Q����r�0�2t6�������dXX�瓨d�Y�F,x�x��U�#�3��E��y�WH6������7�>G�N�g�w�tI�͍fN�JF��I[/)����]ӔB���]�P�U-�i8u�c3�#�b�Ԏ?Ӣ8�XȈ����Y]"�E�$�T��(�bBmZl��}�5��1��i��g��������uw�ì����`�����P�����W�B)��7߄����/��틥���]��Cq4���^�����S���5T����E�C�Xflf�C7j�,����iE����>�[�4o��<g��=��_�H٘�ƟJʎɡ�(:G�7n�����&�{WÇ~��N�����lフp��bs$���n�����Y���]�PF�o���A���O���m+c���v��(��"�Z�j���L�ӓ����"��H��Iq%��D�@/T��s`���W��Z0��K����P��¢u$������(A��2�``��k��>��pF�k�P�ӎ��z)#`�A��R#��.�r��M��ԣ��",Q�;�8�����1������Z��٘�uJ�߇(�����m؊���k��}E�|�{z����Sr5���ۻY^�X�|)�H*F�[[O�S�FU��D��1��2Y���KEL�egx�ڱ!�D"[F&]D�@|��j���q��5�����8O�����4a&�����'�P�F̚^���U���DrY�����C�,u(�Mk����c.��;����5��3�PX�9��{�zv<���s	���Y��`/|tVߢl�����&��b>�h�S;�R�ҿAv��Ul(\8�����n��<���FGg3�����]�սC�v"�ʈ7��!h6-��LՊ�:�m��x,4\�W��ՌK/:O|-�_9K�.GSS'�9��VXvXd�90ʎ*�H�=K^�=,U+��Z��J8���!��ӥ"�j�[T}2Z��+��Cx�S�
5�'X��f#�$\�e,�`���~�4�h��� ?@��f�H��cN}��vj܌.\8\���^o��|�9�1�!:��
.H]��
��m�vy�y.�$Y�V}N:�Ӏi�V4�T�*���Ux�MLi���_ٴi��C��C�7(&Q�PN��)D-�Rɟ�i�L����UӪK�`�a�}�����6�o0	k�{�"���M�ĝwނ�I��ߏ��n�u�C��/��I�Wݓ6�T>9LN�#:�z��Z���4a�#�����U7G���w[0�~��O;��[����(B�ο}�g����f��.d����?=
e)�Q�GRV���e|�Q�?z�XD��t;���E��ġ\ֲ�l�[�x��Ɨ�87�x|~
~J��p�����%k��5A��yn:��Z���HJ�3Ix]N-��ъ�p?�wO̻�"���pϽw!�nu���o���r%�<X������ u���1n�x��3��U��j�3$�7$�J�v_}<Y 4�ӳ®�U�]�p���Y�AE� �X\�ʡL���܀��)bT�&@(�$\	QY�H.
�|.�_u�?__�?ˤsJ$��ˢ�@H�0�FK6�_Vs;<F"��n(��AҫT�.l�4����W@s�j�|� }��?<�ykpM�V���?PiU��{��I���1 D���x���{���c���$mr�=���'ϯV���1�`�d���s���o�F�L����^���뎸����͋�b��]�.X�#�8]���)����l��m�oQ���V�4U�I�يF�~�|��O�!� �y��<����?�D($eϺ�΅�)���Tr�Yv�_���M�S�`�_�vQ��R�
Q��J�,[������ʢݕC�@�h�d1`P�舠�""&��QPQ�Ŝ��(���ɡ��I���+W���~�������z�Z�Ewu��w����9�$p{jhD��b��ql���w�H�����/���	._�ͼo��O�|<��4z����X�nG9>���܊�`LZ�z��hŀ~�q��`��x���ػo7���+PΝd]�8<>�0m2���x�ށ���+NFӂ�b�/v�M�c��T_�y�4�,*�& �ea�d��ǀ�.�..>C�4�u��gj�;ik�	�l\ꃈXǸ/���&PU��FVPy��9a!#�!�ڥ�Lr�EЖ�̙��US��A�D���$+�XM�c�nޫt}��`|~Sۄ�1���J�A���R`3c�Z<��
#q�>���� vUU
�=�Mƭ�Ƌ��{�ܽ{w���oҖ4#h$��r��]�W؎;)6�Ď���];���(�?�]:aO�.u(�����O��ѵ� �o� ���Ǡ }�ha1j� �8��ȼ soI���b 6m@�Oͅ<?P�k�	�ϙ:��I/�3��G���t֮��G%�8PRф���B2�L�z��Z�H1��uHȮ��l��|$��|�V��/=�(r
�"�oI�q���c�;��g�#Pߘ�.�ܙ܈���~'��4�,�D[XN��V��Y8t`_���G�j=�����݉���*�-kv�X���!5+��jH����?��x�&�<@+�O-vrk�ѝZ�x���0n�8�ʬ��*�)8�T?b��d!�X�q�pA(�+��U�A �bd��������z�jIF,x,[U�zn�����2D��q�Q<��#���SOŰaG���[�;�]��&N��ill�	9�5�&����b�<'�Ru�x�LU'�J65cnxs�|�|�,�Iˬ��I���N۷o�����ΐ1ǁ�b�����d~�ypS�n��B��׏��Kѱ[wT7��
cמ�(.*���+1��0�IX�vz�囷c�̻��.���e����Z|��Yޖɿʐ���T�w1�37� �)���g1�R�k��/9���C�Iw�t�c����?g{�).ON��<[�]�qy�� ���+����b�X1}w�[
��r~Ḷ����,�K��]X��s�գ"��d�鿽�[��B�u����ݑ�3Ccm\l~%�L��s!7'��@ ��2Ï�W_y�s	:w� ��t�����ƉO2��9|i��;=sN$ڶA'�Nv5����.�]����f�i-	 <KF�T�D����t���kI�(r��դ��-d��:�!pТ�4i��y)�p�"S,�سg�L��"��Wk����|�����1˙�C$�p�=��#��������1�f���;_|1}t�,^���M����b�^Bp+�-5L�ȸI
޼���gq	
��}x<qG��������t턽{MQon4,K�v�j+O*�� �>x>�WC�<�S↺��L�^��4����K: �L�j��k)������q�-3���?�o�AX�a3&�0�dI鄖h-�<���M�P.Ҁ�� �e��`:7x��K��imP����xpe]]��������{Զ��G�}��!�<�^ ^LMO��j��pX�i���$�L�b0	-2��|��;Fþ�x�q�	�o�v���?����BvQ'8���'��$��Cq�����R��^\q�7�s��z8픓PWS�իVbS��s��S��)Q{H��\5ZI���E|mk�nUTߧkc�@`����hU��u��4*7����
Lv�A���@����	~�	'��O�W_!��i��+8�Se�,^�yy��p�Zŕx}\4�h���+�h�0�`@R���N��_�W_}ULz��z��2�ک���q���+���2�%$���D�X625�&�AY�|i�L��Zm��ݺɀ�U������l��#Y��������ɽ�w��!���Ӛ�{��KƤLr&|_,R1Oȁq#���HJ��KYo쯩�s���훶����q��Ѡ�}ǎ�������СKw�\�)D���M_J˥#_i�室&+���8N$�Y4]8�n��t}N4TnZ=�QS��8XJ]��ԇ��/�)��"�y�v�&i���v	�02��ߜ�zɭ��eǥG3&��46��p���G���㧸��p�k�Fm"��ʵ�1��	�+;��!/�B�z�@,T�HC��xid\�8�z�$�:g�L֏���Ln�����W��Hc�H-�'�*k1�����QS�n��d���KG�>��������ű����	�ڤ�*HS����e5��E������3O�<�1�yoi���;��|���܅�2����p蕱�b&����d1�}��Z���y�;����/���6�<�q+WC �;�~q%�͛'�L �˓)�H+��#��:��96t��%UE�rA^��ܳ�O�����Q�sY�|���%-:�.ŅOKeϞ*Q�ph����f�7ZS�,í�~L��)��`,�F � Gs�$��X�
55u�{�,�"��/��Rơ�z:7M��}�:��XڇH�m]��5�Z´Kd����P�-� �׃��U��9x��{]��-�0?֮ۨ���蘝�� J��#��QW@a�Jv�9c E7�^Hڸ9� �}D����B^V
/�����H��2��4����=H9W 	��"��(�X3��e�K9б8Æ��ǕƪU����_��d�ʲg'�LK���H���� �]a�L$�ժ�P�)���zU�DMq�8DbԖ�՚*`bE=4��a�[����r��9�^o4!��Q.mV���5P������3EYJ�Jmڨ��V[[#@ػwo!�?��S���f*�)��`�	�wʂz��'�8��.�;�C�P<&�0�O�z�Z���@��/�}ɒ��Ь�β�L!%{.vj}�w~��K�����"�Ks6�B�f�Dw��g4>R�Ǥ�3S��y����H���h�W��%n#�:֢]�~=�!S:�i���x���%C�}Đ�岱�$�id�c�Rt�^&��V�bъ�p�x�*a�������f
�q/|��Nys�.��R� ������5����{ZJ6��.���u��WnZ5�O�N�;}��!e�<??Z�mԎ���BW$Aݶ�H�: P��Ȃn(-�aiMj��Y+������e�L��d���"��Mv�Px��g��sC�����%���'Ĕ��KD�DW�N���r�cQ.�~����J���7���+V˄g:?#$a9)Xm����$$�0nX4�P����3�A].(�Ty�P�N��JX�(������H�W�A39c�[a^�.2�d
�q�{��`�G.n�8L��,N��˗���)���n��!�%�0��K/��H[�D<^�k��~��>��2^*N#�;e�L�0A��M0�[a�{�����3��׿��oˌ@,�(�	�"2w���Nk�u[o�u>��;�xmo��� faa��!��D���b�X\n��H�5�Ud�z3&R�k�}1�1''[@�֘ �N�[��Zv}d�|>��aą�^�|��Dȭ�h`��`����]J�~}9�Cr��vW�k�i�c��ur������f"����,�nĜ&4m���	]��M&B)�����
��\?��2zԴ{g^sp���퍔M�g�#��Ag�z}aO�0j�l���~)W`$l�Bq4;D$5܉�Y�������H�$7��~���z?.��T4�5K��ח|�����˟��0���d�����"������uAЙFi��5���_�Em]�$f�VlK�	;�����6�@Y�����׈��`1����q���\��ŉ�w>��(��X�����A-�!w������0��`��`\@���g��tg絰��Fࡇ��S��پ����@��sq�3$C9�x=�Q�y�nb�ȑ���H�
K2�d3~�`��:�\�s�Ε��^�°(]���ǋE�иѽL�6�|�X�$oǍ�RJ>�g��=�@���>�?��3��`�D�h�J�����t�<���ؽ{oF������'�IvΊ㫑+�i��Ka9
�4؅�����͠��5�V�E�o�~_q���X�p�Er��E_���
�1�i�ŖH!����C�"/�kV�����]��/x Ï��+V�ē��;����L���NŮ�Z
�����n/<�*��6��N�M�-��B�&V��&���ґ����7�΁P�x��sЙ;"�Z(v@aMYZ!���&j~ҙ@ґ��g
'[��jnFq��~�����$�y(�V�Ǹ�ӑ�械��#�!F�*Q6�#�M"��\�/�ҿww�v�}�>V�\&�sV�r�H��^(&�cn^a�D7J:� �!e[�x[@Q �Gw(��4ͩdWJ�0�a�j�e@hjj��O�!Y�|Rk��N��܆��TEJ0�>��ea�X�"����ra���bd�S_��M�VM���k5j~��Wi|E��FAtA*���2rD���B�EyF�F&�$Y��<9�c̘1��/� 5�ۢ�v��QղjŨEGKA�F[��*C�_~�%�}�],�}%�>�h̞���y䯲!hdH�[���K0�6l�dj)x+��pS���׆���J�~��N8^�s��M�6��8p�K;��)2jj�9��}�xv��i��JN�]��t�P�\^�z�蕪k�Уk	��˝()*ƶ��8���j�4�ڰy�;��D���1u}c-� z"��bwy(Y.Z(kǜ{�MϺ��4K'�L�����Ϧ��'D�B@q�mP� ��O
ф�9�V&��Rh���m娮*Ǌe?�� WB���^r%6T֢sY$�.�i�����
��4��
��zߣS	J;��ϑ�o?�7m!�V���EN1qKHڸ|q�u+�&Wâ�_k'�tr+_�����j:g>�0�H�u��ebxCZ�{���Շ}��7�{���ס �H��ӯ����ѭ[�w#.I:-&7]ZO<�!�<!W����T������"�:Gɿ�m���M�Bݲe�XI����M	Ǎ�]/^��2a��eb�ǡkF`Ꮎa����r//����r&iޭ[���O�i<�廘|�e��O�T�8��Y6q��5x�%�,Z��\�/�$�x0H沐���N�	�ՑP]W��X�e4F$h}ns
*={�I��ϟcK+��]���hn	I�P6��F����1=����s:��7Jv�ѳ���'�	�l(��N�6w�>Q�{ j"5�rI;	�����	����b7�RP�z��(�6\�˓����R_�y�sN��Н7|��u����4���2��'Pv��B�@)��n� �2�&��A	;�N���$<';�%""���͘7�N\z�(T�ك��p��/c�S/�{��Q��]ďTҁx"&�W��Hǚ�NDp$Qڱ=zti�!��_.�/?}#�R-AD9%;I��O�q�d�	ˉ�[`z��\�mZ�����t�$���%����"e�f� �c�\��y�����`�/nӼ�СC��+Ae�,�
���Ğ��4�v�;��w�#�D�����AHW���ά<�T��	'׍7�(����W�d�8�3��ʄM&�|����2�{����w�Y�`��~�!�o���-�/?��ٳg�W�>���-c�!��)<W$��6~��G�f�t��Cz"��O�$}��-ѡC8��������' ���[B�C�+x�G�,J�T)��JY��<N�E��	� �t�Rq�l��Ȏ�I)�=K�贤�-�$7�	0�ݻW_6t~_�R����||���9}ƌ���*p���Ꮋó/"��`    IDAT����h�&��O��R 譵�6@�P���]7v����Ϻ��Tl[�7�s�=��8�]qw ��8(�P����N��¦�+��B��r;Pt��b�q4�^4�xJ)��؎n��1�<���u���V@cM%
s���h���n;bȠ���%X��w��f� M�h<�S��������]��J�[N8���;�����
D����b�X�om�}E5i��<�GK���:c�+qG۱s��������o�d5�F[�?���.�H½kmDT�ɸ��.hZ�}�]��.Z.4��Y����p����@Q�++���Dl^���[��1g�q9ƌ�� C�ty(rw �*��0�|�lO��{�2+m�H�y^r&bM���M�<	g�qn��Vq���zIz?�曯�b��w��M�?|��-��{����Ͽ�p6�4�
�I��`U 3�Z"���$Vã1��nݹC�1��l݌p$"�4b����](����z���PX۷ߠ�R܉AMM-�m�*�]�q��ѷ� ���u�^�tF]s.�L�D-j�Q)��6����ݨ��XŹ�L�Λ>=(��U�n�>��_6��]q��P���c��
;���v0BN�l��X�J0iܷ�*��o�����w_=�)F�>���S�Qx�����H&bb�!фt�E�^��ӵz���'�����	8�������L]��Í��Iw��'�����ΉCС�����UKD�{h�������2�I�V�@v����4����7x�@YHt�ެD)	qiHnҝ���P)����;"���$`pQ�\�2�ِt�,�dg�u��m�@����(A�sZ$���{��f�������x�m�r���lJ�����ރ�Z��T(d�ݧ��>C�Ü9wa��r��k�I
��M	 ql���3�`��e���Xp�V�^'���?�[n��~�o�o���z2n��IP����圴���[�,�T���:�{QRU,7j8$��X�wf%�Q �����*.*ǒ|�O?�_]��\�[��-�y%��!�%��X��w>Z�-Qx�8d�@d��aٲ§��W��O�[o���+~�)����*p�W�C�ވ��H��h�%$>3I�v��]z�
(N�Un�0��S�ϟ5���6^Z.�����>kW��@��P��"��8SiK�f�#p���Ԍ�|v�K�Ϳ���k܉��r�1u<�L�5�hס#n�u���7(���s��R;����-���"7�BQ���t��G����@v��"�u��ł8��.I�3�sRbh��k,3p�	#$���I%	-�%L�O�TU�N�Z��B�6I�F�4;Yx$+߇��b��tY�?�X\z��X�p�(Z�-��ds�3��k#�G�I<�x������ "Ѡ��@�������?�]Oz�����DԬp�.\���%�u��Q�O�|��J���%��.���%��ڵklh�r�-BO�>S��I�
Pt�ŗ���0��+�
�D1�-���<��sX�f=��DH�^��0g�=ش�B������dC��p��C�?����(S_�3���Xo�*%�"�6m,5�\ֆ��c�b��EE����vlŒ�Gy�f�ci�ʟ��jj@Qa.b�0��Ћ&&)�Gi�L�C��8��  �ê5�
��T_�믿
�M�
֭ñ��k&ތoZOn;Ĝ^��&	5��J�hD}�Ɂ���C�ڼ�sO�1>q����'���6\z��O,d��]Qw�B�ݼ�����|�jRk"��.S?���Fc}���6a���8�x驇Y'��6�؃�nAc܁@a�X���C��jX�5� �3
�3��\��ꆞ�K�~�|��צ+��_���Z���皚�`j��d7�$�X����B��ݻO&��4��2�V\���[#
�@㆓���B+��U�WIMN(]8+�<\ �|���.-�v�/��EE�����p�����?` (�:?wPF9N;�4���	�CM����p�g��`����v��Xq����=�>y�3Mr�<6ǃ'.A��-ݸ��]t���z��6�+-6
9b�I�w��b]�r��]���V�^)�;��q�gbႧ�����gx�޽{b����=�xн��ʯ��>��_2�,�%Q�%u	I-1a�����'e֮�-�Ū���W �B�L �g�����e˖�"6$���8v�Ȍ4@J�`�.ӈ�Ғ�u���է?����֋���P��/�y�u��V�7'�.�t�7���o��ӝ��+Ȗ^ÓNJ.�Fy�ϒsP�*7��;�ͺ��(kkå��<���m�Ȫ����Gn"�jJ�>x����&�I�v8b�1���Ei<�W�p�����������!*2�Sn���[�/l��XDߑ�I�g���Tپ4�})�u��E�h����}�ɘ����+F�HK��tq��5�:u�,�n��52�if�	X�Z�3K�+[�,��ޘ��F�$<���5�#SOKG#
�,���xN%H�K^q�bAPG��U(�O^�c�N���vˈ��VIYñ&�؜��B>��ķ�5&�ՎA]Z!���ˁU�K��y��Z�yZ)F�f�ϋ���AU�.!�i}u�n�iS\y�z��O��	h��i�o��R�KW��#@z�*o�|��X �*6�qtg��IK��(AVS��T����7��>�F9-#\�
�K����p/���ܳ!g5y��d�����гWLZ�O�j䯲X�I,V*w�&���Rs�*� 66�O�1d�pd���eˑ����kq��0����Y_y�X�?�i�}`������7�p<�4�RId12n��x�r�`]�G��5��^~�9��xh֔�(�kZ�^}��������l����a��H5�75�K2��	��rx
�xA$�O�`϶���sq߽w Κ#��03n��7��E{P�w��h>���������7F��P����J,�u�LB���#����H��p��7����'I�����ƍ�d'c� %�4 !�f�`e8�I��,��ݚH�Q�~���U�Tq������Xǉ�Q�.vf������9��(��.˿|�L�9U��Y�H){7Y�d!��y�����]rݜȢϱ)J!I��Lz��`��3��
*���qkhjk�����w����!��+�2)�Ĭ]��p1K~UK.����|,fΜ�M���qYە磛(���Q�r�x߹�y��<�M�ω
T�H�=��p>�)p<�w޿��]�f��c.ç� �>^7�G��_�������/�ݟx�q�wʣх���R�d[���yf�h�p��b���WS�M[6JjHcC<<_��];�0��:�v|��2�wB�ᑶ�N���<YW���� R� \^��@�mW�:}Ƽ�&��X(B�>��o��g�N�|�H��(�o�@q���<��q:��/��?�;ڈ=;�㇯>Y<�@���cN�/�=
;vCC8����٧�����N���6�$χ#�@��ě�_�	��n*�%9QY��h�ނ;8�8.8>�7�|S����t��ג�+���4Gi�k�o+B�V�Bq2jj���2�L�&�q�S��،4p"�x�������C3��xcc�L�Ν��p���<	�^?�k8� ����kq�y�D3(�6\��1�MnCԲR��w�g�/H���)�`�������BqZ��%�q!J��4V?�^��t���@l�@%3]�?��������]:u��3��|��q̛3Q<!�Y�B�����r/T3�$&~�X��B�H����wfSij6cEU���:h�K\	�X7�ݨ�;H���O?]���h=���N�f�I����Ƨ���%�l�^ӗ��9���0��س�mۊ��zt��	�ͽ����I'���~�W\3	�z�E8�~���ÃdFb�Vԓ��/[Z�=I4�ٶ�N�>��(�=��w頳���p4��X� @I<Q\�p ��!/'�:���`���q�8�:�Zi:���D�������o㐁��N�9�q�����a)*=|h}��x���e�F��Ȅc�
�ÝF����)IH���ܵIjq����oE���--���D\&^/)߭r{١,`aȍ���5am~�ף�"��L=�DĢ�E��+-NbQ��M@��d_�j� w0���_/�.Mv.4������4����֮o�W��P��ciTJ�b(h���͎�/�0�T�\��&��{�5I��N�dᷘ\u+��\��ˌ����{q�����>0�]��*�Y�X�I��_�����ƭ���}{�t#y<�97�+;�>I48>|*lT���1��c� �܋�F���qsɩA����i��,���{K$�.����^܄噰h50.��#������޽ѣWO�]��5�ܾ]�=獺 +׮��#���i��ӯ�GnQ{�ON2��%s��ܖ������L@i�ڼ����L��������Br({�~w4�D j,�d�~)�H��C�N�d=�X�7B��,�,_���:���_DN�F���.	�+�nh�DI��g#�dA��1��c.:_|�^|�)�S�ި�01.`�]~��j\5�<���2Q�/p1�ٳ7� �;V$H�������hX~]h+��'+���e��H��*���*ܩ	�L����y}<'�D^(�ji˂�3�	��t��;w:NN�Hr������YSI`�xzbһ��k5������9�(�)8�\�k���N��I`�(U�B�k��v�r���}F��Ʉ�v��4٢e%"�xB�.#ǇI�$�)�װ=�KW�����Q����aZ���ѴM���@�Y:-#�cZFC���"�p�����(iE�H�;�ēp�I'��U��MQ�᳒��2D,�-�[���㗦_�i�8 E�ض}+�TU�����ɓ�}�.���Xډ�/���9�d����5/�1�./R^�� J펊�׏9��93�=8������|���@Z(�H4?��-P\̡���8$���6%�\g{�n�w߂+/;�-I4�b�q�=���/a����e���ۋ��lN^��K.	�3�ۦOC�98q��qMDbQ��Mh�Qv��ϻP�:�йp�۳J��g\5�Yf@�5�?ЂF,E�V�U��������]����e�r���7q[8A�z�-����$�M&�A��NTY,��)�[�.׈$2e�$�fD��.��".@�~$dM��4��x����C�k�P�݌�
�\�%R0�gy\�ϲ@�n������J\�w�Z	��]C�:>!�^`�#�C�*�D��7�hID+/_Ɛ⹫��JZ�paӂ�����f�>ZԈP�.�x)i�&����F��Աc{!����[}��|6��p.p!��������)�u�!iG}���8'��Y�z����hگ��A�u���o
!�� ��+����Ʀ�ھMz
Pƌ��M[q�����s���W�@q�~'X�ɨ�E%eE�T�}ٗ�޾n���o�{�UPDzߢ��n�ړ��H��To݈Dc-<���0u(�tB�
�q����W�b|��'Q�s�ڷ�S/��9�>���e�"��|$�	Y�	�N4�S�%yA=�?�J;�٧�έ���#J@��$��n�E�aذax�տ�S����1u9y6�9�ڰJ3�e�H] բ�w����5� x<.ZNz���ZE�Y���/����=�}Npr �@���駟��3r��P������������oo�X\pjA�3<'y}]� %ϩ�x��M�����ĺ���8���m,xl�M��b���5��b-��Y�
DTj
�6!x��K�c�T|CW��*� ��v:l�w�r8~�u����`�tqq�|W�.�/1����EEr��y�'�ִn$|�1w���#�SGC���k;�쳱j���r�y��5d��$qY�����*X�p��Tx�pK��8����>)�+��T~�y.n�_*���s��GAA>���a��e2_f�y��-���G +�]2IO��B�`P�CQ�;V9t0a���8>��ؿm�ƛƏ�鮃(+�G�0w�Þnϩ�{A@�G¨ٶ� �Ӕ�#��bi��{R-�q'Q��'<t����K$󲺱�]=MI�U���ɴv�7��"�KY�]Jr1�أ�ﯿ��_|�%%Bnќ4m܂�`��$�0���#���������5L��~����:���gTؖ�cJ	�"����E�JU+#2~�0�y^NFbtQq!h�Э����V��̩1;mk/[�.d�wu.� ���Y!m�x<�D,�+?���tS�¸l�6���V�WKG��k���j����/���T�����T����	�eu*�u�Z���Z����|�m�aժBb�R���_aD��[���X%%yZ.R'Ǫy�/-	SH��?��3�̼yI��W�&
��K���n^βڔ�fg�K�� �ҳ���==�X+�r\&��^dMp�?(5dCeQ1��СC$˹�j�訮�~�]u%�+6��sF�9��7>B^Iw�E�$��$$�F�2����m�7�<a�O��Ӄ���2rȍ?��!ԡ �Gv"�=��i��k~'JKA��p%k؋h�n|��(�V$�D�|����#��g��I��L��C2�w2�l���r=	t(���ׯ��퐆�,�LqQ�i��쯮�	�݃;C��m�ꅠ��	�;�N��$
(B,Z;���BhMBN )N�db�f�Yp3���������f���0��xZy^-���hU�;��E-&����u%��YU�u�+��J��(���J%
pX"����~^{
,zO��t��I\�D�|���b+o���oӷY�/���lmkWׄ���A�b����o����駟ữ�nE�O�V�'^�v$3稣���#���y���#�<���ffڴ�ܵZ�n��\	�.��Ɨ&m��%5*^p�T�{�����o��~�ĕ,)ɪ�f�bؗ@���,��ܥ�}.m�N�2�b���x��E���F�>��Ԓ�Q#�Aq������RXҔ`NIK&�?���{��K�vW��.�vۄ+�R����>7�}��gUŽ	[�k؇����R�8r}A�eI4"Z��ξg�v��bGU-�\5��!8��K`Lr	�R߄4cA��>]K��B�~kk��ǐ�z4�p3w䀸X͡��5������s���x1�n�,����(i��Z%v�@�jG4���F�9�ϴl�����dd�����pw5f��$�ʉ�nU�Z�TL%�;��<q"X���ZR2s-@��,B�A�����(m��ĬE��`k��a�R|���Z �R|�d.+_e�ټx|�1�(:�~���L�s���8����"������D��ff��Ȓr_	V��h����ҵ�,ڣ����b�P���J���ŋߐ��M�@�ڞ�~��ulә���2�v� Uٴ�h�Rx�k�}QuA+��f��v���@0y0��ȣ�I$����g��9��+s���'`�������F0����hl
!��k�.ti]�y��jvn��q��n�}�'9�]�>S�=�WO�A(�XZ�Ƶ�7"������f]^N�H��&\|��[28�p_|�=&�t;����H� I+ֺ�U�B��r8�t#Ұ�P��M��X�Dv���Q[W'��8H7L�s��&���ۯ���ߛ�.�\����?��;?��׾�ۣ
F���h����;���;w3r\h!�y�0\w�uBkbA��/Z7$Z�K1ǅ��4�o�o��}��k!0b���V��/�/^]�d��ֱ��FzT�+JR+1�Nv+�I)=����w�K�N�5Y��Vq��gu*:��Lx\rꮐL�s����qQ�ZD4����b��.�uY����ec���b��|�|��s"�JI?-NMj�e��["�ݦ���`,)��%�ya���    IDATA�D�X���|�
I����h��gG/���E"���]I�(+�.R�)L+y��$� ��;��1�ֻ��x���.��
���E �F��}y**�]3fꬉcN���y�?��~(�ɰ1�m�h�nxX����hnA�;�MK���o��;n�(u`W����i3��:�n}�.�@��>'b�&8�M(��)?-�h��D����q���&龗�����&T��-�N�N�:�w�V��;����?�bSyf+?��V��ݱ��j���d��% �������<�9Ѹ��JaR�`�?�d���D�5��	$5���Q�D��{<����.�|�B�Ij���m]�Gd����������z� ����_s�xO��is�T ƅ�����Y@E}Z ����21�ǦP� �c�!po.b=��Ғ�hE�4�N�W��ן���Q�2
w�i��^�r���s]�h!��A!��t�Rj��F�G��x�K�"K9
$�b� ��[�SaZ�u���������b!���a��dá�����P6`i��e�g���f�\������q�Ig�9���G� ��#b	FC���4.��E0�g �rS����t�A���"�������!gVƼ�H<��t�7�F��9��0l�Ҍ�@�D��;��o��c�Ԛ���0���P��0������k|�4\�0zt.B�3�\��֯F"ڈ�����%�C\	��T;o�������K/��c�B4ʪ��Q�d��s
%�����/}_w^�P� �3�ݵ�/�<�\�N���<�\h*���;��pe���!�N���y^r%zM�-���L����e�϶V��dVphˡ�AA�G|���xoj���6���\4�ZP�������\���VG��J��>~��u�&���IW�],�DF���7!x.>��,)��Ґ� ��
w����Y�f��s�U���u޼9X��I<�܋8����b��ɕ|ּg����DT4 RB�>���>�lD={�+���~��g,|l�D�RI�X2ڷ7e(D�� F�T�s@"T�ΤiY���>���s��/D����U�~�lw*CC(�$�p����	�xD�Q�k���+f?� ���g�x\,WW��co�ZDkv�]��HH �������Ǟ�ysf�%�4�0e�mX�n����
����]ꑟ���'�xS-j��P�f5~���	SC�$	�"�UY)���=���<�����:�~[&�#�V_\�Iu��a�~<�T�Ѕ�(	Ӈ��_��� 6}�t!�X�L����bi��gF8�iUiA$.@mT�	DW'C����A�d
@Q.��l�'�VE&�j�������Zp�(pi�W�Z*9R7����K��ss�ɏ�4
(
�T���v^翭)��l�ޙ��f<Y #@ܿ/m�,9<�K��ӂ��'L�M>���ܒ���ozA3ZG�D�qY��.��#�~]�|��/x?�prN��L���
�B���Z���
�EgB�'7/[@��7�~+�����~�e?:w�$�Y"���±����׍����_(�Φ��С��f݇O����@,�F��B��,G�
��TV�O�v���&�;8% i�Pr�y���q�Q�n�@�f'r�)8�1��@ �B�Ƶ��sFv�!�H�>��D��G!H�.�'�xh?��\�ߣ�nߌ��z��)>C���0������
���T��׎q���Ɗ�gA&6<���(٩䦚�v�ľ�}��|��?TX��I��P���xS^?'F�L�wܸq8�~��|��M+������JX흓A��.�]8�ā�2��b���tv�L�Λ�E���k��K`����w�@�jոiJ�R*�r
,	�d>���h35�u�Z�P���*��֊2�Q�rN����s�H���i�[th�����C�(!�wH��R�a۶-x���4�����������y.I:=�$���aH���|!ݙ-�:��z�R�v���5W���&���v�)�/,����3o�uu��ؾ���,����[�n�{f�ȳ'��Ӯ#���{�d�;�nu���6��eWOB�.e�:#I �`+R�c��Tn�0��1�n=X�J^����єv�D�s��g�j8���K�HV�oس����EC]=�� �\u�nۇ���R��M�*�3ـ�]
�E���!�
rJ��tn'U��E'���p3���w�W�x��/�,�DKsX����u�qa(�p�؅]�̈́e-�����8i`DQ3�04	؋.�@�j	����G]CJ��e11|L���D3�.Mb�G�������V:�.v�S0�E`%����G���֝˜úW;�*H�k�c(����
	U�F��qw/-�.�-���7�&�'Ý[D\	*�[%�b�He?J�b�K�;�qnR 켊�<�K(�
+�H�U���W/9c��z�ThԹ��!�pQs\�\�sp�5���c�K�Z)|�2
��� ��=3���ɢ1��ǟ�?��#�,7T@����
�B_q7��8^|�ݺwK�k��8��ťy����C�lv�$5rw�"iK�Ǹ���$���.���~����:\;�*�ߴ�2F���_~_�.=A}(�?xPX�vצӮ�l���Pv�{_���r{=kwS�Ar'�u`׆5p��";A�#��,'V����;�^y�L�/����]�Hʃp�	vI$�u��$ѣ$�zX�rb񰼞��0��98`\�J����"�D��؄�>�\v'�-æ	K;o�����᪛`W�jp����ԐP,ǤB���t�cC׆g���77��ϵ�^#���4����b��Y��ʭ����owm�s�{��."�s^�DG�,j٭�c�U���J�ݪ8%�R������0Y�/�X>r��-����d�h$"`+��D���� �4��dת�a���恱ׯ���v����+��62n�/3�w�8���E�r�9�����sΖh�n|n�8������ɲ��q~p�в���.��9f��`�kU�&C�W�2��w��o�I���ߖ�;g�:*YYr�B�K�8�v���^����:X��]�c���i��|�H�[�"���z��ˇ�h��<�/[(U�7m�<悛f�0���"l�}w���{z8�agU7�D
�X{�m�������Dkv⤣���#��1��W��E/��K�mF��%��W�lwY�(F�}2֭�M��P[�N�Wv*S�"�p$$>#��|w>� ��{�$_��Q%�����Q�r�0˴��n�sAHn��LK�/$b�d��aҤ��8�4R�2�$g�v����d�`y��|'�8B,��^~Y�ϐgF�`��-�Jv�_�}�5[�U�Ū �
>��bwuX�Awl;��P������kE-t��3O�`�{㋲rZn�αcǢkig{�9Q෻r�QKY��["�1��H@a#p�/�t�oY� �Jh��*�*�؟�|�F� 8�0�>�3�RMC��L���D����̈́s�Q�|��WKU�:,S���֋�p�j_-a������i�؝:w�rTҒ��X���+�������"��<��n�b�����Y^�f�Ι���;���`.=�@>�N?�� �N�԰��P����ڋF�|`�u�ע����FcYU���{{����g�o"q�mpb��rӊ4E�,���<8{�L#u(��؋��L@ԑ�������l4��;ш΅A\4�$|��-�����(�$�a=S=�,�0M�����=�kW֬Y'�yӶ���H�MF��m�Ƅ91���0���.C�uCc�Dc(B��"V�0�KK��Y��@B^���Fj���$�̈���t�����]��±���G�¿+�������85p�0o[����m#Y�.�K� ���vU,���b'�(_�)��6���FB����^���ٽ��З�4���z,�d���\g��ާ�����Z+m-��gW"W�5
��=�{q^0����`a��>�H�_Za�?XV	B�ڵ�g��FƵ6D2�)�9$� ��&r*�[�~X]��!�,\�մ^;t�|��ry]9�Y��dBs�n�R���)7L×?,��g_���,�ko-AV~	"l��	����l/�o����cF͘s�ă���*�wܽ�=��o�Y��ND�tL�аs��[���طy�Y8���� ���{�;��:�1'ܾl4�G���w#�P�a�z"ǓĪ����J��'1�Sq{��+)�����SOakd��.(}W)0��QY9,$�t��Ь���HN-�Gt�y�?���gA!9��N|>T������0A��
�$p�P>�F�����	�`�T�v�/l;$u22U��"�#�G�U]��� ����K�;�P$��bR �� �L�5-IxSK����c&ۘ���iK/CR�mV���=� � ��MZ+ƙ��%c�P�(Tq�R��r�T�oYk|f�O~��=���\��h��T�UBwV۰�6-_�?,Q9y�<����#q�i#u�V�M�/Eny`�7�߾��H�"��8��E����_��8�:�Q���f�0Z�bŌ��`����v/n�}��Aa�.X�v.>�"�r����;��TC�6�*����n?��<˪��.������8s��h�d3+���7:�.�͸���㖉���`��(f�>�,_���H:���5!/�F�7���ƺ�?�~�nd|��DX�Io��ޣT"�S.D.`�a�v��
I�g)Gɭ���+a�����TR���k'!�ggZ �:�)
N�'���}z��	C�<�KУ ���J'*��{3��q�t��W�� �����햗Y,�;���2��d�@�q#�(Q[��gIj��L��E���$`�3wf����u��Q��n�(fc���qL��pnl4��\����������e�q��X(�}�?�R�e��f9+����$��kf�5.nr)[�l�
7uy��,��j߱3�,y�׬�~&�b�cs���͵j�&PT\ ��ѣ�lD'�4B�4����/�*.$��r�۾m�D ���G
^[²��زyz����<��=�hW�	�F_"d�#�QO�^/��غnYŃw�<u��|~P8��wG�����G�?c/]�X�D#�n\��}��wa�_�헞��g�X"��>�
�����P�!�4��y���AgkW��hS�� 4509a�sP��)�N�R #F���Z|���yil���!�
�81�����T��ˎge�jԄ�IM�lS�H�2ҕ�b�)A��
5
R��E�s�M�k�ĉ�9i$�x]�x��^�����
�;��-@�{
(J���u�m�Ź[E�?�-}�����M 7�ʳ������χ
Zd�����z��iS��4!e��0-X�0�_���9ٹc���#E���/@�O�ū\���1�N�C�!��s����Ϣz���gn2t�	"�V�۹R����G��)�ù�񣊖��H]f��	.�٦�IZ�R8���k=s�-� ���ytӴb%Qp'��)=QҾ�TL��{�u���r:x(�e1^z�-�
Kvg��8Ϗ-k���wˍ�n������C@{�c�~ru�)��'Ռ��+�Ӵ��=p������``�R8��M��K����� �tH���/iF�߉c��-�P�u�a�J$��_ ���g�q��|P����:�g�yTHHί��6���ꧣ&>u.P�s�ݝ�Ъ[Z�Xu+�8�[I��>+w`��k"�0Ap��u�ف�<+*̐�ʇ�:O��]�Im%�)�j@�d�e�
0jy�Y_��ïVE-,��
(vkG�'�1�5ʣ�zu����鎒�&�p�<�\��#�C�w(b1YLN���0�â|�E�G�����B�#N��~�Zl�n���t<�5׌׃E����ؽ1-37v&�a4��~8&�˽h
��� �sO�sg�.�*���i���X��.-�*������z�l^�=�Hڭ0���<X�A�i��uu��� ?'��;wb��;1���%E`�ZVI����=���"7ۏ�k��2~�mW������y{��e�/x�hб�Ԅ��7ėl���e�o؃���<�R�9cҩ4"iF�����jD�ly�%$M����>޼{wmCI!+�7 ��e��}���ۯ�c��/>�J�Q�HH��L^q�(�1��������;��,Y��[���8�cjm>,U�r��$�3�"�e�]H��p�2⹴��qYLa!�����j���}(_!�m��|�ST���k�?K���~���/@��T�3zu�"���a�L!(�&
L)�+�kdؘ����"�KAB씤�[*����<���P�{[��>v�P��*�0��;�����b,`*�)�i�9Z#�'n�_6ǁ�X�^z�ܟ)�헶����QԮ}F`��^��e�	!Sɧe2PR��E��>���OD꼼���2��>8��mR���ɖl��l���ǌ8�n���k��3�¸��U�C����ػsc�̫�̼k���Q�g/x����N���JY��>$�T �m��6���>��=�h���\5=��������%����{�y� �]�����ڌ��l6t(�����?ߓI�7L�A�㏿���}odY;q���FW2�YI�*�#���h 8Yy?F>�Z*QC��5�����K�QZm��x\��������Bl�6��V�+)Φ���,��kP��G�,�9P�Sz<�V��q�+j�9!p"���yu�T.���Ť��u�g�����nJ네$-<�;�Vų��G-�H,at?V䍖�Y@V�M[��������Z�zL������5�x|%a��Ze��I�Дe�=q^pSѿ�+�q��	����{2'T�D�:��$0��&ҽ� �~�	`�,�
���ةX�t0���d;t�$.�������Q�xj�?�q�5�8;@D�H���s/�r�N=�(<�ҫ��3/���`�=8)�߹��+.�y���P~���3{����@a/Gh7����[U�.>��'�wY���<�ڻ��CϠs�~����s�(B��8���(��b�o?��f?�Nva�w��w)-E�>���;oJ?�VJ�Үس�����|4ނ�"�f���#hU��J�*��ch�N�{��u"�=J湈Xj�<�B'+('��q�.'��LxF)���In�
��� �b;ϡ��f�����9�E+FU�*l�d�ql�k�����j���Zc1��c�$bM�q�7~^�3��%9�o�D��T��YvlK���k���L�7�@�M�S[���/<�����E˕U��k������i��v�"4��Lei
���{�D����ǌ03;��7���p<����*�h�I�ȟ��%���J&%���3{�K�p��vy<b)��9���L�M�r�~i�z�������q������wy���Q�������fξ�ʃ��\~��E��>�.�&D��~$v����_a��Qx����@@M��f�ª-��CsS=��N$"-�9u�1ؼavm݌XK��>�B�nʊS��]��RY]8Z������o�� ���vWF��N$�E�r{�7��> �m�X�`�!���ė�R\��0qw�9�p�f��5�� �}G�]�;f�U})1h_8������sg��x\@LwYݕ�M�q���{�"�$�?&*�n�as�@C�˜Ǹ��>ߣ�ΉK@�u��XhB��;)H�{<&��Y%P\u\8�X�[1���`�d~i%�� ��Wnz,u�xM �	����n�&�9Ntqhy�S��M�lS��WL���V�&S�]#I�}�k`R���&��v�u�ȡ)j�@0�EII�d��Y�z�ir�-[�aҤI���Bͦ�5�P���C����AMu.��bL�nV�]���諮CM: on�d�o۰z��7O�z۸KN���̓���مY���X���xQ5��
l��Kx�gp�'!N��U�q��נK�! [64�!�s����?���o�D�!Ŵ�b��,��*(*���Ps�Hޟ|�ivء2}�x�)�Zd��b�&�X�s`��    IDATqQ�!�o\$T=��χmv��6�
,�6	�^R"���F&�,��jC��E"���( گS !n�
���h�)�nq۬h?�W��up��� �ONP��;A����KW�ca\ jM��=�b�/��JK��82����)`Ą��@����i�ئ@e���18Z��zL}���C/�n�t鱵����#�+I���
n���.7!�<h�9�i���g_�e��;���(H$�g�/�,]{�<�����B�������܈Eٹ OB����#�!s�H ��4�	��|n�5u�6�����8n�17�2����p4�-z�_x��ں~��y�fN�vٹ_�1hk���������li>��G��k����j[��9��T+��v�W�����sx��Ͼ�;��=Ii2A$T�3�����ƚ=X�r9��f�"�1ͨ.�EL߼��s����w�B4�Ė-[�d�ɮ��%�`��;��q0�c����q��bYpw��9uᙒ�Y�Qۚ� vRP��������c������괚X��J+ag�?2��\�Upͨ��%���>;j�pk1!��u�Q	u�(�&���Z�;��δ@��[<_aa� �X���1y�AP8�
(${�u�����MΎ=xc�B��bv���l�KXA�%_&Z��x�����U>M���
vH�W�Ud�a^�!�^cAn^FפѻP$,���PXY��/�R@��ȺNZ|�~Z(fId�^s�Q6A.�]�vػw�4�cE9�C��^-� k�0O(�B�%���l�{��>}�ŏK1n�L>�!p���۸�/�&]?���(?T�v��<�+,acG2���(6|�������N�\����Sg���A�n}���f��v6��[�-��{�6��%��uh���%h���&������{�������b��� (��Msn�d�����CV��~�FJ���{Q�,]xf�Of
 i�G���[?�p�F�<'�,��̾s��W@�_
��4:�n	��0
�8M���7	rX��P$�ONH.��߅(��6?� �I�z�;���SvQ�G�XpNyN�����Q�*'�Y��2!I)�����ªĦ�΁ȁ�#�qҟMx�U������!U���π��6�^9/�uXV��1���l׮D�����������cp����}���;<¡�FoIq�(��VԳic�ȳ�6�g�!c��LJ�(K>�4T3c@$�Z�e�r�U�W׌�'�S/��er�7lz���'\x�W�B�qcݐ)O��۠���n8�	t
F������Y7�Og#��o܀	��g0��gWW�p=F�<M�{P�n���1��)�\lWIK!�h*+w�%q��w`��ؖU԰�?���(LmX�;���������k�G&x<�+��RHU���#Х�ږ��@����PK���k���ZjR����I�?��,���9�6��� �>�$!��)���)�fV*	a�&ZI��L$����VҮ�|�V	�ω����@� D��98y��!�34���O�!Nl��� נ�����j�LB�ҴK��Xb
(�`0�B&��*a@#��,�u���&������ch5k;@�c}^��H�9[�>�J}��p����{@YY%���9�M%���`DAqcv#�0*�:�� �	Ds�Ar��ؙ���U�uz���;�]��V��>�=oػ����J֦�8)~s.�͔ϩ�r��1!9A��d¢ �[��W+�]RdeA[4k�'����B�~.�hǤd��|�i�*�`�<���Z03��g4E>ۃ��f��)�M]�zu��Çˆ��d�����7�'��.�b�X�|�����=��:��v���ɗJn�c���$I���[e��/�'O?$���(x�zl��|b�t�;@v�,�d���
i��)'7H�}����j���֤:*��S�I꒥������3�E������o*�0��|*�5j����ı�Xh*�3���_kt#5�E�бc��@H����<�̻j�d�&��W��Vq*�Yl����k�x4�t�W�!�0	1A��8�@z+�fM[�w1�|7f<��g�Cz�5Tk�y��VC�/�hp-�Mȿ���{�}>�,fS¸���̈́�L���CSƹ�Uc�q2O����<��� ��f~U2��I���ftUd��S"�9"��J�C6CM��5o�儥S�E��푴�4��q?���\�`�Vg�Ա���_>����?�9��U�*��>F��|�v�!:$ۑW�Ry��8k�4h�D�U��)	������=�	��#��s��!��|Œ��=��N�m� ʬ�v�����Ʀ��{Զ�I,)��{6��/_���+u���\y�|3s��6m�e�K
�J���I��?�ٹy��i�ok`��LO�^�d�l���6lzf���Αy�)w�I�2;�+݇����;�B�w�.�g2�G� �ļ>,��mc�8v^����s{������d��� ĘZ�Ծ�4�§�P���%�Qa�J)�aq���v�W,C�Z�j�Zӵs[�*�,�L)�S��c���yj4��iAʀ��{bIu,t�p����1���E�I�19��q��w��G-�L�@SH��Ar��>�U`�j�W�~E�!�qoT���R����) URJc��$u3֜�֛o�\�1>�c��cOjQ�	��Kn}4��1��8Պ�ʥ�k�,2I��s�=[��u@��>�D?���B{�����u�vڢW�ʵ�[E�9���e🎓z�4���l�.����է|т9+��+�v�1��	�L_���^�����6n���%[�J�Vi2�֋$-�L6��[�v�ղ����R/+W�J�$��D�?f�l�m�̟=C�	�,/�4:�%$Y{��]u��U��8_�)�:�U#_{��9�'1��������������������c-<��E��@�k��)��B32Դ7u���񅀠�Y��_1-!���[���G�{4)����h�@9���A�p�%�@p��立��_~��V��PQ���	�8a��cA�zĮ��:F������DŐ��B�&T��w����M�C5�*s��k(���cڠ�*Q9���Rp
S�&m�5����G� �!D�����e���O,�	��M7ܨ�0�=<V���`���/���C��=��(�d��Y��DMD�|O?������o&�?��zr���0ٶc�n�RY�U��J���]���v�LH�&-��y�.�];�ʶoۺ��GF_���ԍ�2m��^WNx㑆��q{�$ʮ_Ɉ+N����G�"�}�M���ǤY��RTf,ziq�4�I����gY�|�|���� 3K23ҴT#�ڶ=�w�@�Z�\�<�ty��Ǧ�[dҤ)���"-)�Bꀢ$\�ycBa���d㩧jQh4v|/.�;���Z�N�y�X�kcG��PPC���DHL78���[=�b�W1�bR� *-58�tx.*����q�b	`��BZ;��ؾ���T���%�k�ro �[�������MA�xg �q�����ش,�Px֐#r@q�2�N�����}'�}�+��A>�!��i`.���!8�w�Ί�&j\a����	97y|s�y�u+�
��^�Rk��}��r��7�W_|�Z�H��?�Da��^���L�u��d(]92#g34��k�.
���.��(i�L���ny�w�U�RVR�%C�R�3��ï���t9�������W_y����|�c�~��c�C�f��W=������W�,�D�|��<7���6W�'ˍ����~#��v�=�"E��RR�'G<H�K6�[.���I'>"5Y
�
u���q?�.֬Y�Ezh!�{���3f�g�}�*xA�\(.��09��P����E�L">|4T~~~8	�U�8/��V�G�ƅ����j�`�y9AߵX��|�r���*�)��z��A%}��`�,AS���Ps)W�gxa W��BNN����nMc��7����u+T�O���֬^�;";! �

�А?s(�ŉ��Z���
�;��}8	�?�k(x'j��� -^�0��!%�_񀒐��q1,��T{�B@��X�m�� ���qo�ir��#1�2��9�1}�j�l�3�ݳ��ozZ��� >��Ʉ����y�����:1x�ٞ�D�3�LV2��ɧ��'�ۺ�LK�:��GJZ�>h�{�Iҧ�A��;�5�\Kӱ��ƌ~�Iu���j���W=��C��ܳ'MRK
�������#%;�JҒ����I��k��J
��x��y�IRV�[͝)k�/�f�4RB՘"�Y�?��T�2X^|�y�	ş2�f�Pf�L�vov��BȂ�leA���?u$<�ōV��0cƌ�O��LHH�d��/ �<6�I�x�5$���@)L&�{�t��,J����8u�̆2ɪgIi4�9觋f�Q��e��@�7��5xN틈`��Ģkuԉ�]�겘{�Tz�O�>; �I�� ���&ܳ�����9<bֹ"e�bF�i �f���yǪ͓��/kj*Ե��n���?��[����JW�f�x���իW5��(��,��=��Y��.���Onצ�شa�S�u�`egg��ԋ��i��Q�m�{<�h��ɑ���N�1;3Cb�))���d�f���GI�Vmeڿf�'�,�6]���;���ꦍ�+7t�c/�nҹ���D���B9�}�<r��R^X.���r�yW��U�IV�*�$�y�2�2�2�t�x�ٯ߁�y�V]���e��=�s5xm��9�+{`B�U�#��'4f?k��xL@ ���.�����]�.X��^��L�����⋺�Y��?�����"��
��ñ�\����m�B9rA�FF��JPm@A�W�, �EjZ��'.��=G��mٺɢw�v(4���������c�Zl	`ł�DB����B�c��1��$��(��v��5k� �M�ͮp��*�dl �=ځ�5����VQ ��� 
s�VM-]�oٲeKu�bC0H�CSAfL��h�B��2d�@�T/��ȑ��X�d[3_��
��{l޼��>���_g���?^e}�}[)�|���VF5%��D��4�xÍ�ȀC���;����6����]�����M=�ik7���ڧc���ʪd�7�ʄۮ���(���}�N9��a���D�2*��l�rۍ�h��o��T֭X&���}Fr�u�g�/X��/	��a�\�q�>��i�f���LI���(\��Ni$`�6m�@��=�"a�j���&�E�w���46l�
!�;y�����܎����}�ZtM���܀^%�oӬ�?�i���2C����U��q\�k�*N��Y8����ء��m�7���Sm�f�h�5�n������_`��~so���*`ƛ;fJU{r8�9��D�]<�'~���5�3@	�����]I�r�l��?�ijqMȻ���\Q��F�@#��6���A[���(�k����q/�
�#�=��ҹc\�X�S��/]�Lyh��m�N�ŵ����d��֬Y=/T��p+�+�R`�����!��h�D�R���ǝx��킋e�V��{�?�܊������i<�ǆpo�oޟ�i�AW<0��z-;��l�ןʧS�H�F�B��ĉ/˽��I���`�2��`�zy�-���U2����v�2I�,���s�pR�D>��!�^y���4w��1cU�)j�`���rU9P��i��r�퉟���^R/�B��ς�L8l��W_�����I�;Ѹ��#_<��E�܋��G�Z�& 
@�_~U`�����j�
^�'��5�ִ��Ν��>$Q�M�AUNS	�����������Z0�߳gw�O
]Z�O�i�&�r?AO�~4g���ߎ���`bT�M"wy�mD]$%Vϱ.|�]�W��V @		٘9�"���cZ�H�P<�*f�T�V��0���	�\����VG����F54Gu7G&,�e�ٯKg���9pU咓SOǻISsS-��O���U�Z8���>3=M�@=G"���C�Nr׽�J��d����-���?�t�!u(��m?���^}4�M���Kg~%�L#�dIU���d��/J��IyU��^�L:�l(C�$+~^"���������J��-x@����n��R��b<�G����qk׮��^�gDRV�u!Gd�	�8�U�0���If�'Bm70h��,�P�A�r�! `��	��j#
C��Ue܊p#�a@`qY��ay�LB���	�� �D �PBP�W�&���chsi�W)�N�2���}�4�B踇Ν�S՛�X��3X1���tUM/�����;$bCbVnT[&t)��Q�-��q&v�W�/���՞���/�3r���;`TkF���A���8;����抯��4��fH`�]� @����Sm���&��ຐ1D^q7�f�d�XE��唵m�f����f9Z)�¦H�u(���ŋ���Z
��)���!��p�z�L���1������Gv�'u��|�~ǡ׏{�����۶�ټr�����UQ*M�i �f�|��7ҩ{oiۮ�L����wʟd�&�����¹s4�8'�&U�[�i��s"��Ͼ���JAa���ꫲqӖ(ʱ�!�ͨ	P,&���Qz9�#(�h��$-͈+���fE���:/��j9�=���ǝ8��V�NBH;����E�b��"��y����Y�N�yZ<D2��.2G�Y8�E��4^��c���<'`�f�� P�qL$. ��{->�n�p.�����i��6v�ׁ#�p��]%E�,o�rk��y��#�Y\��[H�j�Jr5h�}���
��qF�^e����E8�̿si�������v�>�4^����`�z��y睯r�F����w_x$�-1E*�t#|�J7Y~7h��mKqc��d�F�u�LN>�T�P�wd����j�~נ���W7�#%W_;\^y�%����W�����>Ⰿ�P�[�e�����x�.={�Y1_%ˤ�7H�TJbB�\u�?d�O�$w�ƺ�׮�Yn��2)/�)�g̔5+Wh�6��˰��4m��|����J�fHQA�<��Z�7��|��Ie �� �����E��ͱLc���"������E�N�Dz;J-=E`:88x��r6{������/+@.�g���[	�O�ɋaÀ ��ic|�t�e���`�k��d���*�-,��������]�H;v̈́��8��3���(at�9�?�%A�k�fLM�� ş۽?�M`���&��Lč���cNT*s��A�a<�q-��V��1����
9����_�k7����{�뮻E���4@'t��Њh�Y-^���T�IQ�T2�&ZD��(���uY?�<ʿ��5���M�9`�{Ե���X��F����zK��a��7���5C��N �e����ˏ��֧�ϋg������v���W�ܹk���ɖ�y�ڱm��'W�U��)?|��̘��&P5"���,E�RP\ g�{��e���kuٞr��:x��� �}T�9)�̀ś:N�i!�TZP��la�9�٧����F"���.��"H�������i��h����zFNz��?f��Z����<�M��P�|o�����W� �M�N�q���34�@�����{�׬T���c�hن ���s^x��|+uP�����B��dp��Hu2������6�Qr��.H���!���q�����`�l�|�^�{*++�����\���<�񘉆lP����M�h�H�8<bQh܅�
��&,2	9�9�,��i�5��PФ�?�H���]*f�$�	s�F�Y�fx���dԨQ�H�f���<�A~(���S㕯9��sW���Ç�#@�r��!7�{��6]{vY<�{��?j�D    IDAT�������$�@>�h��t�Hٷm;iҬ�Hvf�;�y�7ԋѬqm~����"��;o��n�YV�Z�ZC�EL��K�o�)��1�WA���f�3��'Y�͖-�u@w�ئȞ���v�g����E{���D�gQ�.F�4�9�p��΅5^�p�G��6~��E�*O�:���.�T�w���SPkQ�ynTZ	"`8��
�7 @��p����L!�Ĳ`��R�.=c�Ri���Ď�����b��	�mO�t tr@Qs&p�98U��;��� !�w0�l�i�q�kp3��޿����*Ǉ`�q�P�s�h�� kV�`9���t��8oVZR$;�Ӷ��r(,��m�O�-jƜ��_�i�| �X��s�hi����D2^����Ȳͳ�΄�T��3�1�eM�#F(���>�Xe��"�,%��ɓ�Q����[9j��\7n�oWlr��o<�o������Z^z�~i�U&i�"�&�#c��"�z�T�b��r�=eС�佷_�?�W���d� �F�ɑ������@*�:�ϦaQ���ֻ�j�jTL"��������2��B=�e��x��t' �o�ĉz*!Z
n<xj���}��H������2b^/��ʓ�i�NN�Y}�9LL����;�e(w(�C�
 1h;z�F��7�����H���S�ǘ"��7o��M�	��$��s,�qv
��<�\���DJ<�8(���f�����\Kp/��ǘ��~�2���¹X5���ȼ��sD����s���D
��l4�%E��V-�U����R���[5�o��:�-�?�H6mܡ��6N1ΨA�/!y5[	]d@��G��M�����j�J�n��Bv�ء���-��$;�\9i�Е�^{��G}��ub�|���!�?��f:w�y�72����aY��d�M7���>�VZ�m#e��e��2��KI��拏e���U�,#ЩD��3�W��2{�O2w�O2��1r����������I���혨�U��#b#�KI�r���B�A�u�͙3��r�e�&&���
���]�E���E����sFNW�C�'!P?܉���@H�G�<Ɍg2�ĈB/1�;����Jg�ỀQ�x� ���п���;4U�˩��P�j�l��x@����>�0�c�xx�=��;��I�����Yh6D��5�q�8��?QX|<4�P�sq��M,����C�?*�X8�n�p.=oru$n8���N�IV�*�����R5M|�KNLQ��k�.�>���0�ݷ(�գGw����䠃�c�=U�"5-QǼ~�z��%'H�6�TN��a�`NY[�r�D�LyN�;�<-�N�&,�STP�&������a�V�~��W�|�ɟ�	�|�h��; E@���O}jߎ�;,���|��� �vI�\}�}2�ǅR�QCi�0[*J�d�ygh���_!;�m�̌���I���9�-W^u�
䜹��~N}M�^��
y��$'��z�L@��%P���4L*d��E�xw�֯����=�]�� љlHvj�����\[�'k���M"߁���Įf3&�r�
��}�u-��|��o�����Vk��B+�ݻwO�3~���<���y�i � J��mxs�g�b�x�H�Ǿ��HBs�e�<=ߴO"c�k�=ڼ�f#n�Ҫ��Y�f[�t#�6��5 ����ex�_#4�|N���s�v��umXM�Ěe����
��2�w�)-)��6[�a��J�Ι5[s�p3�rs�'��˗/S�⪫.�;G<��t�@!f	pC���?�(�H��<mK5��:T5�GM}d�{$ȍ�r*BSk����,;�Æ�u�Yu(_����~~B�N];�Z8C>x�A���=���e+�K+v��*ٯMz�1���7e�҅�AΓ� �paK�Y���ﾷ��U"�}�����K�/��,�i�s,��������b$�^t���nm�e�:!^oo���B��y+R��Z3�&%u�E������A�5-�D��M�����|���� 6��\����\�� �9#)))������<�	���{�#��a�
&Q�]��N ��G��y� ���'�a
UƸ�P�	�����f6��M�Q����0T5����R��j�E�.���K�V˯n��񴚇C!�N��>�)����o(��< 6;wm�9@�G{?����٧_E%OͥO�����z�4m�Drss���X疵Dz�s��hSJ&���ФXL[Oje3`�y���'��{���]x�uá`����k�h�q����Ɣ��a�HIA���׋��߶H��d��2��!ҿwwy���d���j��FS�A�б��˗�,�s��?^������m�nU��R}(.8�@&�?��u��L��}W� "�˼Dַ�Uj��L��V��:I�� %��ǂR��z���r����b���&���%��d��<�Q�����x���[c���x"��u�t
��E³���jls��*�mk�&�HL{����"[�1���M�?�B���q���Q\��m�"rص)L==&r�XFi�<�b	-@�8�����ΰr��~���f ¢F� ���+��Fh���\�Z�������z$XC/��x�F֪��w ndL*4N���=MA��.P���cQؾ!@\{�|.l߾�g�}v�$~�����z��'��۲����)�I��"~�!�^x�����ɯ�W˕�M�e$�ӿ�E�H�f�e��1	:P�@���K-�Kt���o�4�΁
A�p!����.ԁb���ɭ	���X2�v�c|�q��v��̜x^�v@���x@qu5�̤(�3�y~_ �������{C/�ϣs�	��'Q����������<���k� 05�1����:~�G̈�D+���4OEu�NM7�p��6�؆�����<y�~�|�I��1|���\��U�8���\��I�.�w��Xu>ƃ�>o-J��t��<�,�p_��<���S^&?����� 6�)�V��ʂ� �zY�Ҫվ���)\��9ϑ���\|�媝���"������a��q.j�dff�JII���3��~oh�Q�o���p�w+���G�nٺC����ț/����"��m�A:Y���]m��G*m��#IU���;oʊ�K�l2�;Qwž�zk�5�믿.���<+W��YL#(p(n���v
mr����C����H��,
��Kp��w�|����͓���'|����ݐ.�b��Fj5��q��B`q��@py�����k���$-�C�2I���J�GZ��/��R_byS��9��xc��AZ��p,S���Fa!�'j�fi����o·�J�ZM�)�E�fj5�(>��:��U���v-w�W��S����E���;%7��,�y�Fn���-Ӧ� _}��t谟F�nߵ[=c��N�iv�<��7��Y�6�/��wH�>pc��:R�������7i�ر2h�Q���>��ʢ���gfJJ����Ou(?��z���"=+�G���呻.�,y����QKNNc��Ζ�O:AZ7m"��̐�?�DC�	����ruka=�����Ā���f��)�a� ޿%$�BaqN�LM
�PKdg�0�,&���uQ=GPa�8��&����޴��z��X;�Uf܏ᳰ�9P����^(^;q��;�@���{��M��Ǹ�ű�9��@�~���} śīi��A��́�Z�ϗ���&M�J�y$'��'&��b�T��ռ�:(z�t��$[�X�I�cy�|>�8��]�A�c�so2�l�6�������96��5�z���@�g��5��2P�v�I�vm$/�Mo)�4U�y�H���!����t���$('��KM!�o֏s,�?"f�yg��el Z�,[\�}�������^ӻw�yu(h(�����m����\9mHoI�w����������n�Y�u.�h�ti�V����,\8O�s̬�1>����&r�7(�$�;oOՈB7y ^{[P�6+6�OwdL�
��~�ě0ph$,"�3�KN��\��c�&eA}�A��J��j�5����Z,���I�p��3s�nұps^4 O�ki�x6��N���,�Ԍ��8r[{X����/+S��F� p�F�!5`��Uz��t�+���&Ÿ�k��dA�|V�=��v|HAm�J<��� %�C�RЉ�L��s56��	(����BR pFj��9�p���U����z��\�k���t�(���b��%�R/;K7�􅕌T���DiѼ�̞=Osz�8�I�:j�\r�%R���<� L�n]�_}�U��n�zq� ʏ+�|�=�a��~)}�4�z�"�]w�L��X7o)�6m���J���/?�i?|�j�t%�z�G=Hf̘�����AP  x���T�&����6p����5�V��	��ͤ8QŠ��8Pw���mi �4q#���C�C!ն���!�������-���D����sz!'+Eh�d��1c�sm����gg�ۅ�k=�W�k ��X����O�V,��MJ��ʘ�V��^���m
b	ޡh����g�}��In�0������xĕ�E��`<]<`ч)���"���[�Y�
�.D���YgJΣ�V��zV9��R)�0�����J
�B�4i�X�?�)A�'�x��k�N�m�|���� Xn��&�T�+4O;�5�9z����7o��N e��E�/��		}u����PS_u��2o�:�T�p��3J6�[/�̕y檭� ��D���o���L������K哏?S��6�L �u��.f�f�L�ﱈ�%�@cMIf�D+­�V�`����m֬ylR}��mPÅ�ׁ��C�9�P�c��~�3�9u�Z��"��s>�����x6����9�6�@��c�¢Fb�ݸ;���Nv������	a�, ����0�^�?7�:Ν�P?�5����h�~q=w���(�"��u̒,�{t-��9(�&I��p�����<��#ϟ�8��[K�x@Q-)Ppi�_���w�e|s˸oOy�Ns�S%�	����3�dHP�KI�m!-[��HZ��
9��c5���4�
`]Qɍ͆x��w��m۶͙2e҅]�tYX'�2k��o�w�ĝ�y}'��Gz�k(�e"�\}�|>m��ﴟ�X�H&<���Y�T>��=�/�S�)�n�.���@<1�y���т�7��]�N���.�z�	��f	���E��뗘�K\�;j��k����;a�`���P����p��� �����}����4
��ع�޼7�oƇFfDN����}�"�r�@�х��0n��w�"�6�Tj�B+DÃ|����]�������C�O6j� ��{����ݫ���K߮Kma7k,�����qx�k��Cn%~��P�s�n�,����ܚ�gק��fݔ�;�R�1��N�<��L�L�"VKM��`ߜ|uSΚ�S�B�[��HC�V�	���"�U�[���tӘ�>B���+UUI{B� f��Gd̘1:7l�|c�����}��.�3e��]\{��I�����~�>�o}ɬ9������+�q�fR��UƎ�_6�\-�O�$;v���T�]��H9�$
Q\�D(�p���oԖ�a�h6]�D�<���iN6�n�m����,��}�NDR���1�"�8�xB.^K�<(�C-#d(���S����ga�F�v@�$�'�ݥ�;/�s��&�H0��EmE#i��p?��]��˫��>BK�� ��ݷm��K��\8'.U#~�j|Z���P���
�ιt�dC�ǳ6Џ7Y� b�O��m[���E�Z1�m;B+��xbE���#���S#|������k��:��v�Ix�Լ�Z�:�@�"�Y�j����z��Q�m��*����'������Q�^��M-�ڊ��9�?���ݺu�_'����_����T&������ҶQ�$���k��˥m�RY�'=p�����h���i�&IN5����ZTT��q���ɘ1cuWc'z���e���1��ɀCa�8��}��;�a�|�u��PE����T7������e��ʹ�l\�u��U�xU94]B�;^-W�R\`C0A���^�](9O�� 4�������!|��3��g��;��"؉1d�kP�!9x �<�5���"��,0�@��6�R��j�p^ێ�Lh� ��h�\I]4�I+�k=����UVTS�+-Ƌ�����k0amX7u����ĤFM�	�߽{�8:�D�ӯ��ph�tSL�̊�8{.w�3����fu �勑u�<�kL��b�W�s�
�RZ�G2235ğ0~bQ����㌆gIgAb� �-g�R>"��Ocǎ��O�>u(?��=��;������J��$I)����2g�:I�L�^=:ʅ�%Ϗ�$�f�R�-�m�ENv��Q�B̟?WC�iz������JaAqdC��4�恝#p-�X�� 7�0�\�cR8᧨/hH�����zA��P B0	�Wk� 0������'(m��|�9k�)�syH<�1,B�M��<����n�g~�Ɗ$&�\���1���r�֓����a7P b��Z�?\���zj� ��	�P~dڒs��q�  ��B&r���cE����r@	�6^�Mt���P��|��dtJ<���EM�
u�R"S��D=����+�۔TIMISy�{q3'P���Y(17v(T�����FI��+$=3]�4�G2h�WT���d�}�(�\z�Z�t�
t�����&##c��?ti�i(3Wn?��N������	��~�HBq�v��^�FR���!�Ȱ�N�[��^V/_!-۴�]�����Ϊ��]�Z#d/��bݽh7J��̌z�'%���Jȗ�Α�+�Ȅ�y�vr�\�WW��G��(���^�]\h(����;��pP�P\@c&P(���(��I;�Mm�4T�_@�FV�I1����r>��o@ ��X>w�og���Mf���{�JBƙ���yQ�ц b-(�Pa��@��]RZj���u^qGgefK�܆�{i��t�w��z墠;/����_ۼ���@�b<�W*%�����rي����,^�T��ܥ��x��2�Ε9?b��/�nP̛㿝��"��1m f-.�B�R��y��
(�bYhh���|���p�����sr��ǂ�{+ܔ<����G�uC��X�{�M#FL�W?����HN�Hy^�=�L)O˖5����n���د�<��32o�OҴEs�娪��R�� f�3�<�U�(�r�=Z6��`����AR�7��?Y���Q�V�'�p�����$P�ޱ0BI_vN�xk:�����ƫ�!ױ7��j�P�'m�6^������z��~;�-�T��V-�C��@��Xp��M�������(�{F �T�nJ��������9?�y��O>Q� Ӗ�!��AP7�(��~�"�y��ݺi�ưpn�q��-��x
 nf���/7��Ԍ�$P|N\�HKJ���T����fvy�;�t?�ԓe��Ezo���5��栬�j ����> J�� xB�]��f�aE�
�
���c!��奚�¦ �C8><!^d�v���v�t��]e pw��f\�O��~���{��4c��?���dۀ��wr����ώ@rS��x{��{��R��#�mR@I�S$S_yS֮\%���� ��'�`3\Ʉ�\ƫ��Rx�i԰�N ^%�aj���,<�� ���&�]z���i�zj�9g��u=Q�i0�Ix>�d��BF��M�ڄdo<J$�� P-��;T��PM���9�ǁ��qҝ,�`M�r6���.Rp�^D�z�[�� ������ZN�;x@�Ρ�.r\�xr�����vPm���V�(
�7^�͜z99�B�-��k�C���y�f2g�<=�1���b�M:��f:�f��S<X��8~!%VZ�/rTsג�    IDATP��a�EEyR��D���z��RЪU5��
,�C�<h���l�=7�����0`I���]Gb���v|ĩD�%nf���$dV=՞��CѼ��Tm���h׮�?a�l���wܡ���ez��J6�9W\q�g�qƢ:�Mn�o��z)ݟ}�i��"y�w�%�]%�˫$��@}�>�7�����ʮ�xx�ݐ�Z1�V���e���ϥQ#��ˎE�4���L�s$��p���=N��N���&T�f��g�F�d�"],"��3a5{�tc|@����v��?��?q��6B����9j��Nd��������NTs��G�`
o��	��E����y�	l��RP��(��Ƹ��1��(����� ��ВEK5��Y�}c� $4W�@++Ug��r	���K��z���e��s�0�Ռ���s���sj�ʕU�&��Q�5�������"`Ѽ�l��.�D���/>�����۷����K�J�&��k�< �oKt�2���.?�)��"jW���}��\�NnP?G�3�$�.��)���6�U9�֭��+���^(�Y̘C�������;w�~�9�bȐ!u(3�=��O>������q#��ݵ%_.��Y��/Ңվ2��G�wޒO?�H�w��T@ٵk��x�JܡQ���}���ݞ�.�O?�\����D#V�w%
�������B�-Fq�H|��y*�9@Ë�M��݅-^���PK�7y��~���Dh2i�������UJ�.�t�j�eut-.gO,�ù��1}��]�G��8�&Bɱ޷����F� l��ܼ�2���;hx�5T�3�2�� /E�TL��(�V�SӒ���X��R+ˠ�D�m�@ܣgD��%d�R��
���s��!�p>9��F 0�n]sGn��<	;��	�������/�J��դ�ޣ�|��wrԑGI��}���GH�\k5�@NI�Lj%�gh�̿ɀ�1 ��[��B���/j¦DyFh0	ԥ�ҶNl�BT[�u|����u��7�����="�f�ҹ׍��\z�����O?��:�y��r��ǞJ�H���#�I�zIR��L.��"Y�~�4h�P^z�9y��7��>�ݻvH��zQ(��FuP��O�4)�*�����] ��.�'P�[���^��~HB!u=K��B�K� �/���
�g��k!�� 
k<����fKy���� ��C��D���w�#��*��r$h���9�<<�؁�Sݷnݮ���W�y�_�B�� �9�|�{����jǔ���$kv���j�R!ބ�o\�8#ܓ�'�4T��nY�|����NxS��5-f�q3-����zRXl�9��(� ���Ƣ�B��33M��r1���׍���v�DIϰ��ŅERYe��*��"�n�&�a�m߶SC�_~�U��aY����
�q�B��;���$KU3E�������h�)�i�p�ŀ��Ds����_z�� �=��e�}<���]Rg&�����1ҳ2{<��=�";YJ��%�v�zi�o���������w�1�;2d�ϱ�Aƻ�KF���MG_�M�H'�]��U��j�:�� x\
Bxh~E��;��Hh��:9v??=���6�%�$�w�HB�9x�?�P��%���Bb؟���ڹs{Tg�\� k�1�ex%68$Z*{3}�����~U�M��9`L�7O�F��m�F5	@��W\��g�px�Hi����>�ک�g���f�:͜����B�ѭ�X��6�c�	p:��bNy~�
V&��u��6�� 9T��=�x�Uu�G�˕�u��ю	�6FÐ�n���%3-]�oߪe8�T���[]�w3΍�����9�8�{����6���w�.N򎍕1RmqO�U��2w?�F3��x����6�G�=��
E��w4j�p�e�]z�i��V7^�ū6zᝣ�g�f�zn�=Ҭ^�T���w��a�f�{�m��c�=&���d��z�"��ؘX~�N}�ᇵ���є�/���@�zQ|�/,'�,�vj��ʊs���ædgî'�uu=�Թ%�� ��C@��%]x8�5zl�P��f��`ɱ$����p�k���T]����ذpxv�, �Fÿi�f��+V+��
�����:�QQ�D����Mk��S�%'�K�d@�2s�̗�;i��"�	��T��4 �.�_��$�]��i~���z$�sI>���iA�́��x����V��	f�\�Hzlq.^�F���hsK�$ƞyhۮ�lټMI���{�Xl�n�0)��߄�S].��ɝhW����"w=�Ht~�#� ��a̚�-
M�1�8��Ju�U�i=5�i��A�Լ,��f͚μ꪿_^g^�y�~?��{��On�ɣ�fY"	�"'�|����-�<\.��"u�Z������TPTs�+v/�>�Ո�E�����[تђ�w(�'���o@�sYx�he-<��ǅ�����6@�W?CaIX��(]8Q�}2!H�w��;NI�h��/$�lj�cq��x���x_f^ے�XT� �g 
���o�n�V��d�@nڴ���r�ڵ�kJ���-�5w� E�Z���3��^Ԓ�h9�D9[���Q���`V�0�<�{׌pN�ک̳ 2�	u��v�!�P��k���@'Dƈg�G��X��h2��aj����>UR��1�T |ٜ,p��rF3f�V�V�!r%*	5�Ql��PT��@���Onn}�\j�������ɸ?����0[)��t�2����{�`SP�GU�4o�l�e�]z��'�X7n�ً?��>2>5;���QwI��IR�/r���HQe�~��r�)��-7ޠ;�.�vU��X�vR�!���������O>���%%{,�/��u�v�ģ=	˅�`i��*�Z��jQ��ٚ����������Pj�݉���/ jk R����=3B��:����D	��w��M5�Eܷo?�(�0��s ���)@eI}���#k׮Q��Gs��� ���L%aq3�,T�Z��I����-���i\ø!sq������"3F�����:����^���pP!3���,lz52�s���G@Qm�7��!N-���$�߽S�P��]�ub�g͙���qH�m"
�Ae'�tB@Pb �[r����'Z����6 +V���Th�1;�c�_��Ay�AG����'++k�W\v�Yg�U7�2}�/�{��'�TV����]��l)�C��ټu��r�_��?+�_}�*1�%k	zd;"�S�}W��6M;�]H�'����` `�5�>ݒØ,��Tn&����v7�11^@�����ɼ��k���l�q-159���G�(�猩�A�}x��o�w��}1!<k��B��	�����+��{�7TcA���8P>�:�}��*3����L�������E��"-5C]�$��J�����JKu�y�sB;�e{�<h33�TyU�gKN��5�Z�{�|s�{��/�2��ha=�y&��Ul�c�N�vN�(n��L�~v�j�hPl^ 2 ύ64{�<�8N�����VC��4�x��/�-���f���0��4��� �-���	r���ǟ�.��r��˯H�B��gLԌ�к7�n�醺��=���ޖ������H��M$�J��s.���5Mn��F9���ɽ��G�-��a�֜:I�CXg&�@*@�q(x ���"���ئ�AD�19^�/)��v�TOC�>�e��uZR�
�d˶�[T%ewd!�N�8�(!/4Q�C͢6��w�6s$�{=_-e	Bp��<����߶mk�>����'�M)̋/�HOGK<0x����s�n���K3���c����T�ՙqD�Fh�����?I��m�[�=n��\���;5�GB�2�lh!�j�ju2������\��\�y����AC�=��MB�<t~�63H_��릤�+H�ג8�P�Gk�P�*#-�w!h2]5����V��r�xol�j�:5s�7�=�_;$f�IY�h\�(�YP�,�  �uF[R%������0�N:�/
|�B~ܸǴ���yUS�c�a�ٯ��#F�vE��<��?��'�<����ǭ��M��%UE"�Pޙ���}�9��S����~�6ti=^Re��ߕ��6������U@��&��[�.&Zw��!B�p(Ԑ`X$p"����{��Ń ���Ύ�+���"���!��X��Y7ǹ��&KmJ��b�Ԧ� @���XY�����0�T�e
A���K���� ഺ$ ��'��5����y ��]$�s�L�6S���}��4x ���7�t����G�K/�)�~��·�Em1���e� �<��5��f8ߠ�b^�6ncg@ �aÆ)��%L܃�ש�ٻV,�^�]xE�%:n^���6�Q�V�����<��I�Ê���L�q�z4�BC!Ί{oۡ�V���= ���뺗2,&nX1�%�8�K)�$�k¼a�7j�O}��ДȪ�m�y�Qy뭷�+�;��Ú�>5j4��k����H����r���W������e��S�dG��}�~���S2f�(9�O�ʇ| OM��Ev������ jي����GW&�g���j�C'e�����'���IG#�8�
���Ph"Ah&�2~�ɼZ������J;7�N����A���B�do����|��bgX���B����0�Ė���"T=F,|�ǭK�����[�o~���-����Ç�BE;�{�H4�ݛ*w�e��:�����a\����	�
wx4ؠv��Z�|՟a<y&�={�v`mMi���}� X(���p�<V��Cܩ� T���7l�� �YO1�GnZJuv;�������i5]S�iΕ���&ٽ��x���N������ߠ��5�ԊE�Z�j4��d)&�YkU�u���ML�dfeH�F�Y���8��]����_ωi�Tm��:�߾]G�S��Q�MI�����׭��|��G]7n�o�z���{,37�S��by�%'Q��ߖ'�'/>��Hy�j�'<��3�� 5�h+��"g�y��4c�M�'��`$V�"���P��C� D@{��e� ` >��{gG&z��}&�]n��1�M�)�W�7aj�<���\����;��j~�Лo��W�_��ĵ�`�{4�E���x"t�U�2-�k��u�L����v�AGV�1�u�~�ŊpA�Sa��E�h�M�ѣGɊ�HS'YC��&B����.w-�wbnv]<$qr���4ն J4/�9�H^��q��{���<�4h�W�ݹ[{त�Y �(gWV�p��M,r�N K������?�`����\u�׷ޜ��v�Ͻ�
ؕ�b���.c�&�rf߳�?�Q����i��}kS�"�9YҼپ2t�ɱx���_F�-�F��޽�j�Y@G��䄪�ʪ��z��u��͒������7n�r����'GJz��}%�)�����8}���~�7��+Z�u�sI � U���P�o��:�V�7� ?G�D�m`���Dn�CX0�ش,LL��������#��N�@Q�\	�SBs'�P�p���������TM#(�(���v�=B!���^n�㼾GƋ��ko@�#��}�v��AF��t��#2�uSӢu�z���?�x��b�bf��Y��rD����?.�~T�
��l#)b�˜�0�-��ͳ1G
�Y�Y 3�s���)4N4�|���`�}Vk`��(2vOI���M�Z1+�	� ­Z4��ƀcy��hR�Վٶm�,��3�6j�cE����\��{���֖Zݲ�7�x���@�Ա�[+Rrv�Qe5��Vc ��9g�Km���m�ݡ)0$�b�2~ߓ�P��_0��;@�r��!7<:i|��m��ܲV^w��W���~�\y���֛���]y�p�"y���,_N�tU]!eɧar��[	��4�������l����$J�X4���>���[oՁ�����L�Q9uŋ��ޚX��p��f��/��v��n JhZ�f��/.�-v?��{y�$����-B�όkS��&������i.^T�/��:2/��2*?&ma^�L��f���V�)�rn��Nk�<P�C ���M�.��ʜ 
��N�� �` �m۶׹��-���5�G- ����'����XB��8l�?���
�5����Wr+�tAd�!7��&��=���j))��N:A�y��ҿ�A��g_��%�T�p�Ii/J�R�2��\S(q�H�z]�dG����p��D��|�y�g��~O�8Q|p�6KMI����9��S����g�{�?�:thݘ<�/�t�u�>3�y붝��6�scn�l�q�<����s�N���M	@v�geJ��dɁ$+�x�5�u�?ơL|�qj�G����<���s/�	^K�N�
��� ?��w\���cC�63$~bk���P�H�PB�������?F~w�� xn5_V�Tυyi�Z����+���NH7l�X� /����8wm�D����Ӿ�:�B�d�N,߃������Y�����	�$��������^���L�"ee���5W|����̵=g�|~��������V�x�wm H����q4��V��Jij�� - �\׶�q?�f}��ҍkw�n9�A�p��#�=U�5cd�ۅ�2ϩ�����w��2%-��(񬑵VȌ���wA,�����#��H�#���R����$V���9��+�Pl:�	S&4kժS��u��wJZ��w�+w�v����˲f�*�2�YY��7�k��zD��B`( �֣Gw� e�P|�#��� o۱MmD��t��EUu4/O�ˀ"X\C�}T�~D-HL<7\89gh��;�[����%ܡ�ܐ���F�s��4�/�wA@���]cK0�>4:��\wI�-����**��uvb#@�����<���A�^���Y�z�E�F�8�;r���jh��V\�4/��7�h|ΆA~���kU����`�<c�1��G�¨����s�m(Jι�2�鵷n٢r�E�������i�~��aŲqV�	jmZ*����T���K@@��,�*Z`b
�=ҴH��w���x��eYͿ(���Wn�֏<h�!QR5I+(Z;%"�5~���*�_crʩg����k��V��SN>M5V���%U����ǌy��uF�~�t��7=��M۴휿~��=�n�/"��'W\q�Lzz������OM�e�W�b땖�Q��%�BT%��}��Q@a҉�$��G����.��%��.�Ir�a@=������{�&�w<"� B�5�JB ��8 �$��c�&!�����5K�d��?xLG�/��MT�1+(�p��-�,�D/nd^���t+Ɗ1"���L_�,K�3wlR���Mc3�#� ��P��s ������kD,�]�wH�n=�;W�> %+���W0��Ґ���)x�H䆱�|�4�m;�| � <+U�1	W�Y��I{%��"V ��c��Q�A��i' /r�w 8���Y�t�x� }�vHtG������F]t�ͬ�*���]̝������H^~�j�|_9���P�?�]��>�2�٣�zJ83��LJJ�6z����8∺���岍��x��t��ҟTC�%�d�����eĈ��QN��1B~^�Br�Jrb�>�x��}U�?��}�0~�SZG #���PR�G#%��0i��*���E����@J�`�ۼ 届c�(�Q���=���8�hv� *A���&�l���"�/�,^#r �!�gu��u���l׾�>+���b�D�ۯ��ޘ�A��cS�ɣ⼌��Ŗ�`損�k%ܓ
g���;xP��8 v=�.ü�m�Xc�sz�r�̛ǱxP�/����\$�gKsM���m3����D��|��$��n�V�ły�L�ҥ���/�Y÷܆5�Qc��KE6�I*���w�T"�|���p��0��J{q*���͛I��:�k�hdl����k�e]�    IDAT�^]�+ܬ|��+�Y�BzF�r'&�	Z��=;���%�'�p�ig�J��9R�L�7N�5m��8�k��6�v��'��իWݴ"�z��#.����}�z�4���eh����2q�kr�yäi�\�����p�i�O#�S���a߇�A�:�5y�1��*�O�0�)�0�����N����N�"��	����`��)�1���#��ۧ�&��{3y<�,�P b��z#�F�ƛP, � F��v�Z쬻v���&��1�ژ5΍���� ��B\e`���Afjhط}n`W]$�� �x�B��ɕC9L5�L̽�x�8��:��	�����ubXI�h�7��S6
'f=rR���|��U�<�R�(�H]�j��c��=5��@J5�*"'@�X�����Y$���f��X'dL���T�x&��QC��6M9�&d�1�rWb�5}É�����J�2�(�-�LJ#y�5�@��p��cE��L<�m��r�UW�\E�RQ�~?>nx�޽���k�q����{ؐ^��.Î;\�?�pY�d�L�q�t谟��ʔ�'N����qh�H�7z䠁z��?��ƪ�����N�4�̝*�q���rs��"Ho� �"e�&s��<�K\��͖F޵k'Y���b�bB�?����g1�,jr�?�޲��M���
5W�0nH��.�V�y�=��F>`{�e��z� �wm�<2<'
����9�5
���) D�r/8�n{�b�v��FvS@D�����D5mx��X����Ut�7�0�!q2<C��-)Q~ �׷�~��z�>چ�Ɛ��wZ�֘&��>�����Fv,�*�0�,X{>kKڢ�5�߰a�z�֯�E��Is8�d�(�Д�K(����.��=U7-t�"�(���5 ������6&ϣ�>�w ��k��.,ʯlҤ����=<�[�nK�7�������_��0��1/��}ؐ���!'�]��xY�x�,Y�V�=6m�P�x�5�9s�$�%K�"�MJ�mUsx�W4A&�wT*]qLJr����eQ�h��Xr+���A�@}�l ���hC����e��%�+�6 ��˃�r>~|�t28�����h�T�v�EZ�B�I�+4�����r��c��0"a�x�f ���{���b5{�z{0\5�m��>΃蘔�����Q|�0��Y� �0q/c�zw���,,��v�r΅{qm��9����� �[���������'��M�sŽ�|�a��t�8S�e�6
X;u����������yFK6+�G�xR�B8oa^����c���-�{�z=ʛD����PBYa,����b����K��m~�Ol>97�Ͻ��p�I�9� 1q�3����BנkM�y�Z��r�؇��ԩ��u(���e���9�ˁ��]9�Gܫ�< @@��p�	�a�*Y�|���4����3�L����V�s�%I���tpv���E (�ƾ��{��<�Q�V���j_0(�d��U��B�DP]�O`�"��kԯ��i�T��|j1�qk�e�'�c"����k%T#%4[j�$g����[��5"��z��K�b�/����t������"ݶ���$׵]�v~^\�5��rO#���b.3�@������=c�]��z���\ffژ�F�o���,v��8�0cQ2����{��>'���v\b��y�],|��b�<����`� (������ܽ�J�&G��e�q  �J�����kaQ��v�ȩ�#I)�RZR��~sr���VX�72���rʑ� F��[P���;�y�kd�g���S���`�"�s^{��� J�N�}>r��w��$����F���q���G��v��_W-��g�S��#%�wʜYs4��s���K/�G�~�$aVY����v��j��vJ���� A�e�ˍr�x-*)�Ip���L8���ʱq~~�u̎����UOS�o��UU=���*�]�7y��j��4�P��cC�(9h
�����^�&�#��&җcvpj���˸y|���eq� ���p{��_��2�3�A�*�֚���ͮ<�d�|��jZ .~^ƙ��A7�<��4.K��Eƃ�oMz��6 P��ӵuS8i�niٲ����.<x9���h�����-����Z=z��ҠHӖm[��ɮg�[�% �{�� ��īv�������{��dNzsS-�1V36��	5ט,UZU�����E�' ��y~��裏�
^\�,q�^lD��r�ΛG�����#ﹱC�ԣ��P>\���<;uT������:)޸Z�{�N�WV"Ӿ�J~��W��1C�ߞ��"sJ�n�r]�uQeܸ��$ڄ�رu�$��4�܌�OGC����BZ�[l���䯐$G�{�oڴ����Gq��qOD&ZNL��Um�K8�^ѫ*΋@fV�+�3�x��A���@t���Am�X�iW^:�ݦhv>�D]�BT ��&���w쀃J�>}��	�6�*ͽ�3�+B�%�z*M�!R�����?���{�<�������D�/��h�ܗ�J<�9眧��Rx _ ͣ���uF�+����4n��f�}�\�<*E�13oMQ�U����ƀ�,���ժ��������6��^b!&ow��N�-;��.f,P'HY���U�?�T%)�0�L�·ǎ�gu@)*.(�ׯ߇w�y��:t�㵼�O5���?tĤ�h�����6m���~"�):6�M���?/������Ͻ������#!a�y��ӧ�%�\��p_<ӦMWU�a�ƺC���܇r�&���fPi���<^˩(�hQ�i��&��<��tOs*�@�5�@�2�bƕ�����l�ޢ�:��ǈ޸bK�1�NxZ���
��lW׺%Q�s��ģ�P5.��c͜�����b���z������h!��\�H\���~�G��|p1���j�f�#����4ϛ��e�X�f�&:w���=V�0	2|�u����0�\�߮���̼��Q/K5Z���~�J��@v�����fvF�~n|�H��l���`��<�Ix����	h3.����ܗ/`�_C�̛�j��C�z(��iQ�KIO�#fτ�㤬����X%��0�!��lt�|o�1 W�[qAy���1⶛[�n��N e�u��5���������ir��]��Δ��B���r���j�A�ѿ8;�ݡ|D����R�;C�QHTȽ���F�;x���q��g�c��Ixc7ڱc�j(L6��Q��-�@: 67EeB7��k����
~�G����k T���1ہ�~��$�~7^�u����{R'ъ ;��Ad�+�ќJF|� <��L+M�{J�6<����w�}#����b1�A����O!���FN��qm������X�Mƛ�aA@vbN �-��1U��6^y�%��'���-C�W~8���)&�gq׭�'�z�tRj�.d���;�@����\�d +�Tn��P3���KFr��A�HM�+5@��6G�A6yȻy���;����}q��Q��,*��E�b���cdm Θ��;�����	4dȟ�8����hn�O��~-;���?���;oiժժ:���=h���lڥ��E�����r@�$yz䕲u�FY�p�t��]���޻���0�
ڨ"5IA ����e�i��Y�by��y���c�|�@uCa�<�ҥK�s�o�G��Tk֬�����+�����^�f�k,����_+�D�BM\9���9���<\��c]�3/����[`��5v�tm����<;q|��M���a�W�Y�x�_�Vͼg��Y��_E�����.��tӊ���r3��t��NM'�s�E�����8�\ 	32�͂�9Q+��¹�w��y���ȅ�B�c�.��!p[�i#�}7M��`����i����+�*�������k�(�\��I��$M�����.l��Qb:E���oT�
��͢*�6�\��b����x;(��#]׍��R+K �D���1C�q"x��`�=��m3��,��I$�,	$�r	�;����Wu���Fx���]KKݷ�=a���]�W�_�<MM���<,�_��W����{D��eG����?w���z�С���<o�aWM|��ƽƟؖ.J��OdH~�L���%��Y6�Y%�xR���?w�<��2l��RߜT�S'2��LZ,7�H����J��>?�ў����m�d��"��ct�߶[{z��!Cuw�H��]�q�<C��g����D{���޲%k%���dֆ2il�`�����\@!l����q%�hc�5@'9�)�G`2f�N�K�`��㺎+���32��'���Ģ�v��K�E�5A�nd!�����3�3�>��Ź��۽�h��k�ļBޓ��\mlT �b3cs��m�V�,s΃eL_dw��'�8��s�">�nC�S�}�`(=�ھ�������q@���b|Il��� �3a�kk�+�&�[_��fz$r,���KA��ˮ,Yi|/�Meƌ��e�]r����{\�'����N��n��4g"�h���Y2�Ke��ղ�w%S�b�AM��H�A{ҕ�N�Q�6LS���ᯠ=WcQ�f���8
�t���ћa Y��8H�Щ�	�@`Ĺ�~�8�ދ��gz[(�w��Y�M�C�(�]��	��Z
\�:
>���Ba�x+����9&�W��]B��/1Q�2���tƂ����b!�HY��p�M�9>�1�&h���.�~�ՁŁu��q�����kU���9��z`�;{�Z<\?ϔ<��������/E���ɋ�����Eǫ���$aaa�@�-k���n�YO��Jl�ͣ� $�!.~na�G��5r�'���F�T�� � =Y�9A������Hy GE��" HM�����\ (z�WeUy�#�8�����˛��V�������������>��xኚ=����TL��i���+��S�(~�dY��<�#���_.��/���V'1y��Mǿ��ߩ�:"H���8�ioC��̈�X�������c*zȑI�w<,��s\�	A����w�
O���.���[H�ޖI�+�il�������v��s�Iv�Ri8��R��y������ٕ}��`5� (��:��v���ԍ L��?��e��E�����z �	/���V
���6]�׃��+ׁ�ı���|a�q�Z#ԙV���N������P�)�{<QN�F�D�rł��dY��˶���J	���<�y���	�t1�ͦ���$a0PnC-	�E|��ϔ���[7Ou�DeF�(�y ���{���}��4
 pg�����T-ajy��9�ȣKa{̈́�����~⢋.����a�n���Y9��_��fā_��)���D>^ e�WɌ�-[eݦ-V���"��u�tuX����5�_������E�B�ō���������ٞ�Ʉ����bc���L�Z�vT����p2����Cq3��[�R� ����2!�F���]�ǉ��C�չJ�-�9������PX�N���L`Ϭ�d8ϺK��S-�R��m�b⛼�b|�=��1��M05x�FYx����=�����1��Y��]�s#��s:�ܳ�
h߁�ɵ8���H"�ߩy���82&מ(/S>�S�79_OG�����ͽ��y�Us����Ȼ��k$$�����9`�
�ƹ0���f=N��.Q\F� ��֐�3�=�(�R��{B���k��Ns�~��Ƚtbࠦ��Ç>��_��\���_=��{���z�q�o�H���>m�d���d�+��c�&�=�}�6�_+�1Y�h��\LZ*%M��Le�Iҁm�t�̛;?𽃔���g��c���9�H� (v*&-��0׉𰻲�1y��s�_�>�>e���K�l�B!�A'a�wˣ7���ῇ-��։���nβK=d�d2�`�.n�a&��,��<��x�&�����TV�䁖F$-W��c]"D�u L\��vl�Ws|�pt~lX��J�U�s1O�`���K5
C�;�R��H0l|v+W��_ƥ�Έ^�m���ˀ��X���	�,�m.|?�2�1(�E����g����WĈq�Tpa0b��ZE T�9����S��3=n��v�P��įm&�:��W���al�<��0t����9�L����|TGGG����ŗ�5j�Dy&����+�|U���_���D!'};7�Go='3'O���`��ȥ�ɢ��u�k*%/ e���l�$�*1?����7^K����Lт�3|�;-N8���5' �Q�7����L��]'8��$���lZ&��HaK`W�Hآ0��� P�n?3A��xɾ����Xa0qp�x߯�v`��T:�;-*�Xd�_w?�_���x&���)Dؚ��ޤ�ON8
 �qb2�������>�i��g���1�D�x���,n3�M&�E�D�?Ǣ_;=�D�Y�D�|��dR
6_:�H]$lBg�u�n��� �qems/�0��V0σ�ɠ���¢�ld��Xt�a�t:�H��^�V�v���Q�w�f*�y˷���>� �D�R��6���s�},�O����8�y�)O���!O�N��D:n)�ýb5���W�\��5�\s�n�)s����G^�:6h��2	�f��?�C�}�>��u���q����kB��D��ѪU�����ʤN$�W[K��c
:K�2�Jأ2��:�=ڲm�T�+ԪXo[Օϛ�h�;'����]2x��[��Գ��u4͟LK@ߛ�έ;P����~�*��l|o����3�'�{T��h��{r�vថv��k�Z�@��t�`"8b�7>����q9rϒv(�ɘ���xj;�<��a����n�.��M+��4�s\υ]�_�>jQZ���l� ���O�i�J�U�$F&�%xA�g�9"o����>�#�p\,K��g�|!�7��m��Htk��ӲO{X�A�>os���k$ ��	k�_O�[�j���uM�Q�)wR0��l�)1���,�8����k��
R��Hf�^jČ�����PSW��@il�s�G&�y?��|��S��`�`X����Zg̘1c	d������-��G_�&2d��ק�R��dD,+�=.#�:e��G�I�G�W�1Ǟ �lV~{��\�$�6R���ă���^������O�D4Oʂ�v5��g0���o(I�C��套��d��&��>c4]����z<�  ��D"�����R80�u�@q��am�]�X-��7���v����H��t�$�Ju������:c��r��M���&	n����)�2Fp[����HPhV����`|8 ���:�Ewv2~����ba"���Y� 7$�~pc��� ��.S"�`�p��c��瀸�h���A���\��$��w6 	�r��P���H`y؂6n��Ay�@��[pY4�,�V1sN]��UckG�B�b�5���}��឵uv)Hڱ�#�T�@����T�;p��N�`�F�V�#��|6��Z<i�PFO7�_����r�u׫�R���wu�ʥ����!=a��/�u�]��@��^�F��9}}gB$���|��}�E�i[+�<��dRm�;t��-���	�Nu��]>_�IIt�3��OT$��-IUk#��+伞����֞{�E�.���ij���Ld� �ʪu0�!!�� �$�eқ?)�	$����Z���Yت�����@�֌?xw_<\��C�\�F��v�a��I�x/cK;/j�����{MM%�>�	`�ν�;ɸ��A�y�5�#��k c��y�?�����J�����I�������sm�������UW]��͜�5�u�?"5_t7��[�l�>?��F���n�#P��7@!�=l���\;��4=p� |����!��$z�\Tg����ˣ����{�cEy�В��ٯ��    IDAT�l<��"�WIᠭ������w�x�% ��Y�1���ƌ����Qu;�L����w��6}�&��\�L��9�}�X�}�م�n����&�^@��c/]������Og�o�N��h��������rи}�K/��.�Xz�Ay�3D�ŲD�s`B0Ah���\�Ǉ|D}4���e,��x(8�B,,&��zҘ~���R�AZ��MK���29�V��΄I3�2�ͽ�f�{��t@���<J���|b��h$ �ȴ<�.�7�e��f]�M����߰�<��x����s� ��G� aTv~jv�9s��eZa�]��
,G��"����0�}8� �񉪰�s_L` �� �j��I���<c���x��k�n|ˇT{&8� 9bOm��3vk@��8�'ۑH��eIj�W�U�,��(�*�-\3_���.�x4�ű�HQ�ŨQ{��i��U��X(�])��ȵ3&��8����{䄵�D�'�.?�:�J���TŞ�Z}��7ĳ斷nk�������/�J$����:���+X�*��/}�K�����&=�����P������a���1��|:#�[�KŎOd���Ϗ�'�&�\r�|��U+��M�+QƯa� Y�d�]-+yx�^xI���:�e�����j���@a��������x� ޓ�XD 
�ޑ���c ҳ�J�p���Aތ� 6����gSzk&*c߃�aVMNwg��l(�\	$#�G������49��&-�d�)��B���� 
n\ �g��b�x�S������9r�V,A��΄�ZHY�
��Z�9�[�s�M\�0'҄X��e0'21l�Ԋ�lg[(��zq(%@��o�Ό��n�7��FN�'2w�ܡ��_:R�����S�Ћ�å[��Cu3����[�Bf� p�o0��y �����ՕR^an�E��%�8X��\VKc ��7ޒ�O?C����&d�f��릺�Fv6�J*�Qr�����6�I^4zw>���}o~��k{���T��Ri�n�*]��Kn�R�_��W^�*������Z"
j"G��S9 `�111���Ф�ݒ�+tgj�cQ��W��Uƾ�k�AP��՛��(�ܥ�M���x�'�O��˃������Hs���'~P¿�XA>�Hea1Ytp�r~&��`<���Z�)Q'k�n�>Z� A�5�ј�XL>B��<x��'%�*�Z���8,���;�e�Mh�	��̎�/\�8��X1�t��'*�󝳾�@I��}56ʫ��(U�r�@	�9H����B��=��P��ӏED&���A�`�=�T�����0��V�2�$2 �ƺZ��@3�sʀ�����ua�g�0���c{z�YDA#� �\[]%U��^�\� @alu���)7�|��|�e��]FeE�К��j��ri��c�?��k����&>0��1#vS��#�����_�:1|߯oL'$ۙ��Ν����d@�E�]��g����ܷߐ}��-S�yN�/Z(]��'����ț:�)�Q�9�X�1��D�\�<�K`A8�idZ$ B�FP�r�@�l�脳�n���M�O��E}.Wj��V����-e�=�1���{�����	�V�0��M������%����u00��������n*����p*��baa��� M/`K��M:��cLn^�N�C��}T���;�m�P]m��,����ju�8/��bd��ڔ�ZKhL������z���>�^�x��A���n0��;B�Y�q���K��^�v�Č��\�_7J�9�&ꚿ�[C���0��c0p ���
�&f�@'X�~��ՄB��#�PU)5�X�6��Pv�yN�o���r?��2u�3������$��H�)5o�9��/�^ѱb��'?��E#v'����+WŇ�{�Ʈ�d:�R�c�t�Y,M�vY�p�}�x����ӏ>$��/S�>-/��lݴٴ`���.����������IĠS[�=�`�8�����8�@��7��wW�3ե� �b�P]9�K���͛����!<��f��9�"�^��Gp|���k8�I9�Ϯ����L:��v횠4��c{��]�)���t��_Au1nVQ/΅+ ;���p���e�Z��
kp��C�;���������cI�<y�����s��<X�b�r���F��e��=\7�ۭR����0��7�� n��-��&�@o/j��=�]
v(χ�b�<Xk� z�a�Q#U��g�+��7�f<;��%e+�g��9�hժU���`�㋅���1Y�_ 
4��Y�/�8f��a�^����c��}�뭊 ���<���>�e��1��yg�ڏV�0u�S�h��=�<�Z�ϟ�z���бgnɔI�3-5�;d����Kj#)Ar�ܷe��ɑ_8D�/\(�_w�J
�
� ��Ȅ�:�(͂Čcs�� ��䩔���_p���L�K�� ��b�/R<5�ʉO��_�0%�-�~>0�}RyKLg����cs|"$ޞ��Ë�a���)��ͭ&��D�8&� �.6푙�YY�<avO�kik֐3 K���-*�W�h/O#Jdјd	��J�w�o�w���ŗ&δU���[w�u�^F�5J�G{�Q%K}�\��r9,o�W� ��{Il���^y'|V7��#�~���m���9�8R�6���_��W:V�<p�H*(�SaY�N�b}(��}���&��&"r����j�|��ߕ�&=���܀�j�T��C�P�RWS��Hk{�~����<�����N��c�?��r�9���W��i8^�ղ��U�399��h�Вe��[[v<�ȣ_2v�n�����1����cC�~mk& J�l_6_���K7��u+������eق�e���A������֞��Ƃ s�L�l��r	� �=�.�CV���X
1?c�����4["���9���
�-����+�&}E��;�I�B�[�r��`Ab���Y�D��<�*���*k���7��p-p�f��-���54LP��,<<�a5*�C�&/Ee�$��5z��>\逸�*7�p�	�䙣 ��X���.��H}�k�*��p2XS �y��T�y�9yz�T]n5��Nb�[h�o�'(
\�	y"=��gW ߈�"�]˲�����Ƣ&$�eŵ-�^�D�Os�U���˂����.[�mӐ2ϛq�?�S�UE�p��%�Y=^�9�:F���D��Yy�6���>������y%���-�L���֖�K�ڿ9��m-��B.Y�<k��h����I��;�q�g��?U�+��i���P2�iiHwȇ�-�%�ɂ�]�P�>����䵗_�	��3S��Y��="�<hbR���A�Vɸqh�E�r$�:�5�3���zq��/L <Qv$vP�K���5�t'L:�we������;��Y���� ��9�C�zH��XcX1L&&!Q�������IN��n,|�>�ϳ����u�hGb�S�j��3SF�1��hK�w󦭪��8�;�}�vb�c9��5kN���9�aG(� $ #�@t�
;%K�ۣN�F���q׉1u ���@�nnx���Ӟ�`5-����t>�����|��p�;A�d�sf-��2��3X�dy �aU��c^Wd}��*ʙ�vE��+K�O��?�cu\��!u�~�ƠI�	�Ŭ�	
�}4��X-삥J�q̜?�+��l޴]�Og*���6�7��1�J�eg{�4$�;R,Y�5�%��'������ڰ� e���bC����tR��]R�钭�Jf�F�S!�wɆU�dΫ�Ku<"�7[w�eK�C�t8�٩D�x�q��M7�Tj`t�}uL&̔�бsN��y� ���v��e���~�m�i����E[�i�8�&�v&m�f�c�W){*:�?�-��q��וʔ�ȼ��D1,B@�}�f�Â>b�ZxL
;9),T@�kf�^���Y*P��c��)|��	�,�s@������OLQ���%���=p\���Yq���>vn�q-�/�"O��LV���$Ԫz>@Wk������˰5�M�w���>&j�|��n���b�Hwհ��.?Н���2^�G�q���5ǵc̞z�)U�٭7��1�a�gR]fy�]tڊ0��-Z�u����U.���ܭZE#Ԧ�I�>�A�����p��n��������s��?����k�z-�;5"�L�K!��ά}�IҞ-Ȃ��y��xd҃w���#�Wo�-�r��co{z���!{��=�t{F�3]�n�����HFj*��r�,���?ȗ��9�������Ws��/�1{��
G���˥o�F}`k�|�Y�,R&��O?��Cm":�q��'��;5���g�2�x�M]�]|{��s��x�����aU�L
&�YQV��.�,ް���ä��|� ���&��}RX��E,L��$�s-�c:�5��c��@�"������r�LH"*XGK�.B�E��'f2co�Z�X�b���n��;l���%%I!%�5���~\57L�3�<MV�X-�]v�4�
�"v�Z*ʽh�/�E����xEs/�gB������u������%7�)�Am@�#��ś~���D�p;�m)n4s7����3�p���6䋚/"��tuvj����5&����}�E���l���$�,6�8u�����Kc�P��F�>/-rMeu�<t|�\r��r��IuU��ؾ��F�&�҅����#�|�l�Hɪ5�0�;
�Ԥ��r��Pr�����u�!{��#����4沲��YR�K2��LW�d�7�ɇ��{�z�l��,S���L��o�.u5ՒI��OC�邖�uw��:<
n��h�M���w�Fd|�7�zdǳY���e�]q��l�r�<aW�{뭷���p�}������ʮ���LE_�`���, ���V>��ezL@Le�xpct?7�g. �$q]�.�o}�
��9�>��;2	9VG�5��*�����-���� �	�&g���z�L��輒^��0����G'�[o�ֆP$�a	��@$�`��R��F��g�$������l���)l}8Hmr˄�a�w���t�(����p��� EZ��ݼ�ߓQ���?ys82��%�ϑ[B<7�ҁ&�7qv6��*ˤ��^f1������y8k滺���g�t����J	������@�-f"a�ם��z��?��4|���W3��J$N'��r�'�[s�K�Z��G���~`��F����-Jo@I���6��}$���"����J�m�wn�9��$[�l�i/<+k>�Hf�~G���ASj�Q&�̙okālK����ؙ�RVf�	�����?Hkn$- ���Q�&�r��d'e!��c��{/X���8O��~��� � @�X�,n��Ik}����v�I���Jq��\'�8�Z�����w���;\��{h���=ܲesPӲ��������1%4�L�?:��O���E�[y�-�(��u޿�Tf�`A�rm�k^���<HN9�T5���� ���',R��0^�-m�\]ٌ(�Z�!�Xl�wk�5�Q�`��/�d:O��^ =]��J=�W>��n�Xx�9Z��9����D���p~N��s0~My�\F�]�!�m�u����dg�v�^I��0a�Z̞�E���B�*+ʥ���ܩ,�:m޶�������Բ?묳�y(-�;�{�m���I����F�����$���DDb�=������@�u������ꎬ�[c6+��+�LJj�b��2�����˙�/屼�Z�X�:���3S%��\38�vS�ea!���裏���Cu 'O�"�̜-���m�SM�LF'(Nk���%��⃐t�?oA(Kh�Ki��8��;��܌u�9� *,@��r^Zt���,u[�5p����8z����3a��ph�2Q��>g��er�	Ǫu�5X�ϋ��ֵ"jyQ��dw׭(Vd߁���yXLpj� G��d*�IT�| ���a� �mY���zuI6�½���<e�,~2��C�&�D{XVQw�`a�,�W�����ʡ|�t�2Ɵ��Eݓ(ai�մ7+���n@aw��s�)���4ӕ��Q�z���˜L�L���{�%�����h$0���vT��dܮ�d����}ak�TҊ+��9FY�b�>R]]�2
.���3�!C�S���k���n�Y�46�~}��ةE_�h�x��1RHT��-�R�TB$�^[��t�]�ttM�<�]���Q���X�ϭ�θ^����bR�_s9�h�,��e�"���|�K�)/f��g�g��"ߟ#�Z*?�Pjk*J
S�l��ص!�&�w��x�q������{F��-$�Ddgg��,����e���M`7>�h#�H-�4�Q]�0��	Ϥfg�lO{)+�����v����L �4��;Vw�JX�K��5��	(����>H]H"��E���3v?�� �[D�*����r�LT*�\VQC���N�ۣ"��.����Y�p�up�?���̞��~߬2�N��⮴���ҋn�$]]��!x;C6�8�P�uĄh	VA2��F�.�h�*_�=h����,IGꎯmH��5c�n���� ��v!�H��	��Y�F7HY�$�_ݪ���,�X�6��/�Lޙ5[�� ��ްa���ܯ��h�I����5��bN-�|`����=�:���<pq���H$�*�ͥ74�i�>/��!h}�������?'������.P������s�������{_Y��&�ҙ��Z)OD�j�G��K��Gv�&@Y��mϼ}�4�:mG�|��LJ�-�'L�lF
��VdRұm��}��Ҷ}�����R�(ʜYoJ2V��r*}sZ���ѥ=j��Gv����7)����!�����W��e=�� c��<Q�?�����`�3���i���3q���>���/Be���A>k՜��,:��	�,X)�Å���4�����a�߽��I�y���z�na-,]�\'L?���1Y<�u�6���b��%����zR�D�`Ƕ�ҷo�`</� �C,��y-zea�X��8^���e	�js0�B��X�����3�����E�Fs|
�Q���S��BN�����*o�r�*�l �-:�/sjt&)G^Q��K$B�I�9:��|A�<ü���IMR�\'��	����"����Z ٿ��AL���E�r�̦ϔ��<n��B��:.j���
D*4�  ��ŭ	w���F�<Y�.�%�Q˖�Jm�d�������;�"�ߒs�>K��������$+%���I����B�������du�$c�֚�<�����1i�-�r��+��������<m{�Z`֧:e��P���D��(K(��l�(}��rԡ㥮�L�����,�۶H��Ѥ!ăs���x���o�7^]*i�����O�EKk&�-�_��ń`a��I��'km&;�]][-t�G����	�f���.���<|\�Z���bl޼Qù�Z!� ����Z�D� �k9�GL0_P��,�\�N���b� *0�w�~�Z|�3{��S2w4 �4R� �2R�U��#FUSS�; �t\��D4�D��4�D]�P[�t��k�r8ncd��'�Q�J�@�]8��N�Ǯ����N�k��X/���o�y�6���ׁ1 ��o�����sfk�P��*�A�,��4"��}3������7�����zz�^4���g�q�ZU�Z��Ǖ��N-J�^�ɘ�<ZH�/�{�/��Md6�<���s�=G-�[n���[ĐR��^�ʳ6�kkk���*��R�;�{�F�x]q��r�m����_ ����ت�|�x��#<ۈ��x����YHU�P�W�H<�m�M'=��m��X��.^�T���W���io_��?�k[�Qɦ�R��5�+չ�$Dh�bA��h�Kb�.9�cd��eȀi۾Q���SW�- �,cA7(�ϝ'�y�m��SO�����u �    IDAT��t29A�iY �Lrw+����p׮[+�^{�,[�\M}�������LL� �K�� ��D�� �}�Y9묳tw�L��e���t�L%i΋������Y� ԃ<\r%<����#��=@�R��9��|!��i�@�)�}�s���{��]�P1�s����Ef��Z./�ڔ��iؓ4u����fɲ�D���W���ֶ#(�m��;��~�c����	���F��~�#ټu���G?�h�����G�3aӥ{�;���s98�J���P�4	Ц��������b\����\w�K�P���\"Ӝly�<��o�]�͛�?��ʫ�TY�j6�8 `���1�6Q���%��1��?�;��{���o��#ٮvi��O�sIe�+:���e�d��V)�;D���̎�d������g�L��|̄��^��3����a��]�᜙ʡTƢ�E'4�%屢�GE:Zw������X���4T�e�K�K.ݦ%�X;�A��?�HCt�}��'�	��ƛ`��Qm�t��< �%x�6),7`��%}��A,&����?�P0���$#����ƙ�:0�!Qo��f%���D"Y���Bb�|_0f)� /�k(����巿�Rw,S@ R�5o$��	�8�����̎�n�n�$���;��*\>; �L��gw+L&䧺/Abׯ@[�bF�؁��@z'f�Hʩd��3��FI�w�%����Fw������u6c
�fa�����2a½%}W�^�ې�=���8���wPr�q�y���4b�X���[6�$U���O>^�9E�\r�n^N��y�C	�h#,�ޡT_�e���y~$��$)����9x��T��!C,u�����h�x�7�ԩS���^���QRW]%5�B�O�'e��A�w�`yk�\�&%Q�� ���V�(<���w��_$b=Y��-��]��3��)��B�Ȧ%Qd�`��%V�I!�%ET�j���o�g�|T��cr�=�K!�!5Ւ�L!^�]���6��ɲ߾��-M����10␱泆�������4�{(9)�Ո�t���ʭ����� ���^��(���݀�1�Y"�^n���4�.��F�� +��;���ʡ��"j�EX5��٩��
��{�}���28)�c�<gY �s�����n~�|��,�u ��*����W ����Z*s�����6��tG��l�#U��"���]�l���7���w�����rՕW�9Q7��&�Rٶm�V���{T��Rn�S2�	�Q�ԣgNO���[D��p�4���)����`���;���1
��ނC�T�����KDM����SN=I9�c���9s��Bp<'���X6OħF�?�����V�{�<��U����7ߒk��Z[��S�f�RY� �v��Y�QV��,;�y��;Xe/f��'�O<�؝���X���T��7�,TV�ߟ+ J����$ A@��-H���LW�T$�Jn�B�S��$�t�l߰F�~�%��L�>J���Y!�0d�`U9?�S4I��1���F�aAb���~=���:�.��L�,[�T�}���}��~�Z�a��Č}��"�Wwuu��C~�<	_�v�6���PEPhE��)dLN�e�f����?�I��Ձ%����wxy��kXX^��$�1f�*���!�@�Tx��	;���h�'��s��V4��wn']�1q7�C��G�����5�������~/sޝ�|��8�r��a�z�.�
�A�k��-u�s1��&�Y���WK�`����=��\GMuu��f\��ؘ��G"<����X_�����?=�)�R��=�9 ��eab� ���#�̹.��!_5'&ș�2�EZD8���������t&׻|�
-��c����)���e����˒�Iy�TA*����r��[k�������G6�&e������RCP U�)�p�l�dqJQ��:+I!捹X�Xz"���ʄ�� g~�Dy��i2��d�����$c�Ȫ2���4���۵Jx�����)w�}oЄʒ�<����V�B�v'\�yk�Ă��Du.,5�+����J���hW��_����8�ā���gBt���W1˄4x&r&G�M���??_����hX��J�5X�J���Fa�0�h���7Ll���T�Ԁ���{�]���[JA���P4yٌEc����[*�?���N��C�!�<��X �}�i��(� ��K/�Tޟ��F� ^�!YmC��b����qy*�+$�50[J�.&��&��8���Ãp��b�7��P��Ҥ�J� Z.���Ks,�M��[�h�n,x����~W�^0l�����E�8q��KC}�e�'�K��bM-*q1݄T"��J�7c�}����ʫT�1%�o�fZv�uHyC�ER[� ��IVHg>"�ƾ��c����x�����=wS�@�{���s�m}�!|m�C>^0W*Ȑ���.u1�Z�a,.�.���ѼM��o�s��5y��g��wߒ�CH'�X��j��2�r��7���==m|�˞8�iJ%k��UZXÜ���BM�=�b��VG�E�_E�#�;�0�,02U�N���:��ux��'=���LWV�jV�5~g!������P �p7����߯��Iu�2&`�ag_�� ��^��2�Dn9hD(k"L��z�����T�JdOw����Ԙxt��w��_P��$��wޑ��͑�A�$(�����O~,Gq�̜9K3��9J	�'�4�'��JUM�t�;�����xd���CkS������5��n�-�+��"�ٗ����7j�4/'�&9_WQQ���^8�F}ǧ�*�"�5iA8��,���o���C�\sP���(N�HZ6�n/5Ul�D4(86�D�P]��c�<#��tfr�����a{Hg*'[�[%K��d�HY�Fђ��Ґ�?��#w\�?�����.ς1wO�4����˓�x$�PtG�n)�1�6i�J�ч,�[7�췦K2�%.u��)uj����zY�n�TVWɳS���M��+%�_�F%���(�j�Lt�Q|��E�y�����Mvy�3�n
($�1�U�)��n�>X�Z��yo���ILv��܄U�"nը��ZY�u-?���9��KY��Wp�<��s�����j<��ws�	�+ly�-2�zΚ��T�b����OGD&�4Q
��y]�@��G�U��^ڻڥ_#8	q]��ѪcFj?��
`E�r��������޼q����iD,���x,��8���z�9	ߍ���˜��1,��]p��<����̱�peIgP��ú&h�<m^�֭���HX���3�o���j�^f.b9�	y�J,����8�P|��� 1�;Yπ6V�?����6�[��yꩧT���RVQ&�w�I��ҧi��ߴU�q'��%��jM�TUUJ�إ���#w\��tg{��j�R��io]Wl����]�_Q��.�,�@*sX%���;~>Ј�c)�$VȨ�s�^#eɼY�a�Ji�.�b�5�¹�2|�<��3��C�	����+�L�*d��-[��['�`�`ZZ�&CQw�~xiw�|����4!)k��>�u,T�1�xu���7�R��5�Rn"c�0�TD��UAiLX�i�y�s HpA����p@�oDjV���k�+��]�b�ƨ�=��I u��c����{a��gY4���`��_�B݇�O?M~�Q������R z8|�]�Μd�����ʥP�L8-[��ˋ~��뢋.28��=�� ��8q��Zx�ꭄ,��c����,ܲ%_��v#,f\��{s�06�S�R9�; �|qݚtʂ�#L���ZE����:GE�BY9}v�+�9F�>�tn�� �!I^���x���U��IM�&�;l�l��!���I�kħ XN!b���py���;/߭�r�so\2� %����6�d��RI�@r�3_-f����+�2RN�b�S*9��C%۾M��qi�.��j���4��t&'{�=Z#�r�&:1��D��m:)�>i|�YV�Y(���$s�&�E���d*�VsԽӛ;u��Br���S�v vm����T�w��:1���y�_�b���{]�ѕ׽f�}w&?��8���9:l���H�dw~G��uGMJ.C4�f+ts�ϢYEƃ]�������8S���k�R3�޼F�q�1������:�5�]墨I"}��o��.�I��s�/1��=�[X~�a@�k���KѪ zG�Y-��bv��EA�%)X(� p��,}�2��dy�rsyy&�K*�Cx��Q�Җ@d�f�S�K�l��� J6OG�*�C u)� ]2�q����r�
X��X�ǔfc���o���e�Eґʪu�/Ƅ�PVS���,vlm��~b�]��D:{&ݠ�Y��y�Ķ�<����cOې�I.����VY�d�T��+�BҰ�W!j9$�$c�dR��fe��#d�~2����e��:X��Y���d%��ˊ�5'��:��s(
���R�yυ`&y�t���,�����;{���h�������&��,E�t�äQ�� �L\[��d��tvj8�c�?N�k&
��k�g���:A[[Q3�\�R��wf�X��מ�b	�<�LQ#� >&=�5���]h`�;�Br#�%*�������al�B&���ܥ:���L���x�}��o�)pP�׏��r��ulqX�|����I-�����C��B������]���7 ,���_B�3�
�˅ �����Qe;��Zǜ�E�R@�
��P�b���}��t��ڟ��-�B�_&.�f)-C�ҵ�{�5��	я�L�gH�9�8��y����6���:�<L��IY�q�H���tITTK+E�5uRUY&eҹ�1�}��G�v�n�Pzc�>7>1���=����t^���Y6,] 5�>� %y�G��I|L�K\���Ԗe�QC��1#d�̷�7^�~}A��Z�p%���ޝ)�v�Lz�q)+�^�������5��J�^�`(����0�`�v��7��_�� 
���I�A
�:vW�\��U�j�Io��ϢBe�Jk��)�������A�qlj��C��h��Ձ�+Äd��ՠi�A�v�0N�!t�aK%���x�X@%.�N��̄��<$'r�X���Ͼ�d����Ӳ�^c5����[g����3�0�K/���	�q衇kX@A�lgx�2�O���I.�O �K�^͝�7����q�����½ڪZD: �y�Z���r���KZT��g^j��@��gd�h�+�e.��ڋ��2��c�TT%5��5��}�+_S�h�-��E�Sd��n�&�qGW��UTI��!��%#�ZR����4��x�d�b�����r)��Mu��Ó����F�N|k�7>��5�ǝ�R޺S6.[(�Q@)h�f^�P�IV(��řMj���e`}���-��ꥋ��OF��ۿ� %e�Zw��ŋ�k���5x���,�S��vG1��o1j �Y�����v{ܕ��ۄ��DvY/D<��0�II�֤���(z���ft�Y-쪮V�c��|���@��@Ru@��S�M���Pܗ�� zX(R��+a ��Ϛ�ND�B:��V*��f�<��װ�믽��Р�2~<`óc�>���@lR^>@5z��+V��p�Yg�����7^�!W�	0ѢG��3��(��?{}�ў�������
6�WW3���1�I��G��@te��}徉(�>v�>���l�&����y�^^��-��nR6'y�� U�>���L�HN*�+�0e�~���9�;�B:t�����Ef ssæ�r���RH�˚���ҕ�de��I:_�de��TY.��M���C���w���A+�n��{��[��Ҋ�u�lY�D�0�Hls�^ZUZ��[�3��U��E*bY)v5��?�W�k�@���?�*LG�#v܌�E46�iz;������S6m�&��-j��rנ�Wq�P�qûq�Ba������Ga�����b�-��
,'vlv�������k���'��RN<�$9���e���
��k,[�B����3Lo�`e���������Ba�ǯ�qW�G�s"`��V �(LK�	�Y�h���\c��K3��������T%�	�Ѿ�jkR��r�h�Q���69`܁�o���W�̞��,Y�H����|��J}������?g������OdM��̥"zMTX�kV�U������g͔�&?�L@��Uf��Fu����vV�2]sQcR�,�V�k��0�	
!� ���G3~�8��p��x��r�����">Fm��,�;��@9��Cd����^�)�lm���F��/u�dE�F���UJmu��S�ʳ<��W�6@�������7&G�=ikgN"v�Vٲb�T����:����b�'J���k��S8�.{m��s���?o�UKJ��}Ux�&�$�����a�2�����[��AǕ�U�c>k�5p�������!n��Y߫���.2�$��6Eb&>�5��ب)��a2��G���+V�҆�o����; �A$x��aZ��n�[#�}��v��8h��7��S�k�������]��	E]�X0�ys�X�������O?]^xn�Zj^�\�� �.i��,'�T�����_w�lٸI�,_&5�U�Ɇ�����p,���ό�V�E�X��yFf5��o�'jnG����:,�DԒ(9���B����Ң�#/����Ӥ��]U�p����[M�-W�F��5[YZ0�޺U�t�K^bфU`G����� �i���߽M�R�>��|~���Z��Xߠ��hUw'_�z�!C��~�3y�����M�H��J9=MՏƤ�8TTK}M�HW˦!e�?��(^^��������1'm�Ȋ��ݼ]�_;��H�2˘MH<P̊
�c)N�P���x�K�#r�qG�ʅ�d�{�H�&�A��"5T�驛�,S������-��i���%�\�K:Q�s��`o���)������Q [8�[�vԴ�w����� vMQ����݂�x�[��)��Bwɏ��ca�;a�0)ۛ�	�_O��z��
Pt�?l��ｄ?���vfI~�<:�y[xLhܑ�;P�J^y�UM�#��BnM����~�;~�i\EB�N*3^���%�ai'W��wa��F{� ����.^�xbi��DU\�Ϩ�]�"fXĚX���w�{����G���#F���$�X��G�炅��9;hQ�Ľr���S�5��a��}:1���d������tܾ���e��c�v�袋u�;F�g���)��rh��R�j�1��o˖��$��T����Ŝ)ƒ"�
����6�/����zh$bu�x�S�P�e�������{���=���l��%^��[>\VJ�������#_?�x���[e��eҧ�^�0�3�>e�Zu���7�p��y��d֬���
&�){)��:1��9zGo��^�j9���R� ����.�PLh��Ƌ�yј[6�@�<'Z�o��拾��`����gJ�Du��;��v�#^t��<�.I���p\��o��-��|����]i�k�xB>���X,T�T�&�>�tK��9w�
���		[v���Y	���mm��J�x��:�--;���<�rkz�iJ}���`������X�;��k�g�nˊU+eʔ)���9�|�J]���Ch��ڲX4���L��kV	��>��@��YS_���k�+5i���MF�Lɲry��G��7��PY��j�h9���l^��99�����M�dފ5RQ�O�#��jy�����	}�s&r���W�'Nx�/W��D,F��(���
(����P��\�.Ϯ,�h�u4��3�9�IY1#���2jX���W�=#ӞyJ*���D$b1�x�Ll&%�5X�{� 7l�!2��b����35��,��y�l�RG�C�<(Yc�����q�#�h.N��B�I�
�W���D�\��5F_d���-��=�H���
C�3��z�j�]p`��'��"�+������Z�t
�|�8IY1�#��z�5v|6	�/hCƅ��Ʊk�ˬ*���$9    IDAT=�3���t��5\z�%��~���D0�ѷ���1���aHog������ĈÔ�i�٬�8g�\��&��=`�@�8��0�uO>����u�����5?��BY��ؽT��9K�Q�r�y�aҿi�΍s�=W���_��W�1�ٺu��J:��q�%��֕�چF9��˜���5�XU����x_���F�	��z_Q.e�Ԧ���	���(�N_t�mϽy�[(�\A�;�}
P��C���dg���h^�$�K2��X�S��E�w��r����g'?!+�.�p$my��i=�A�%����7��*�L�-�N���[/#��^��8��ֿ:��7����N
`��AŮ�ew7��w^^5��Ԓ)X��G-�ޭ�0h(=pA�H���?��¨���(�D76��[n��K.�9e�TY����\>�֛�k%2�G-�����	/�R�s��t ��Bd,=5�1��ֿhtd�;o��-5� �8��I�
()�xιg�F�'�m-�
,�t<��ܮ��ˋ.����fz%Tb���-*aA�O�	�-k�T9��X&�*R�	:&�������e:p�x�܁J�E˥S�Hp'��D,!yT�$*��;X2��,]�Z���B�.���4NDL=PŤ
E)�i�*�l��C������� (y���C�:qs[Fbhf���)@��ǪKPlA�4-�EM=ɩ*~��E�W�WO��lX�R�����S,�b�Ţ�	�5��L��V���;���B�hH�ZG�c�on�'�нc���.O)5�M��H��}��¢J^����c�M�I�]��M�����[?zm����z[+�]��n��e(�~}�@C�����̈́&��P����	����k��<&�,z�1;�E��1�Y"�������xu�Uع��#�	l� ߦ��j��}��Jj��7��u�S_'3^{U%xF�/ҟ�(�#j�}�P%�	�B�B�$k�|����0��v��t���)|�ɧ|E�(���+3^}M/^��+/�>�wy�IQ��H�F��2ÆQ �9,Q>rB�_y�e�k�=�[�Y����E�L>*u���#��y����-��|4)8;D�
HzRN	I*-u��M8ݺ�u��	��v��r��o���	[�M�7��;�%ē�WJ7�x�J$$�k����d�J�k� i�J���G�{Ａ\JN���wJu��h� ��霜q�ץ��Q�Ĩ�\�f�sY���G�OY,%�gBܮ���e�%��.�"�g[$�E�U�ޘL�SAj<��[6�|�E�U{�9��3����S>����
pTJ��B�ZL��@��`�g�]��ߪs���*������S0�n%�4�N����g�f�Ksڦ�EҮ2Иy��,�ҁHA��Htc� �=f�|��i��㏭�7��E���T�jQ ��<�G'=��&�8��A�j�a�KGW�	��5����o/�\��7n�_���������'�T$nWT�͢�h����u��J
R��uJ]�=G�*�H�fRS�{��T��Қ|A�3j�F㚬��2j��R׷Iޙ3_"�r��MT(�h��֌mx�V���U�k�j^?������ӟv#�,?�_�)2x����B�� ����p�@��t� (�� )�I�r��_�x1+Ӟ�*[7��rBy�����E��x�w6�@@+���.�r%��&e}Q��G������?k1�w<ltO52H$Zv��5x4���Ǡ׋�d�/�U�n�8��\�p�`H (��g�@aw,��J	h�Zϕ�鹛�)ן��LڈNS��R@aA��=�m�W70�Oo��<����ȒY_fY��q����E��k�%��Jg�z����T`ĹQH�<X!�x����DDm���w@FA��S�����
[�l���sU[�����1��O>٠
t��SC�.K�5��E�(e	�Z�g\Z���M�r"Ӧ��BـIMM�FI)yP�J��#j���$��?T>Z�E/�P�$�]9�����$q�����%^Q#5U";?޿������H$b*a�x�S�<�<w���͹#��ԑ�xA$�usw
�
9��Z�]��������:�E��j�������(M�Ur�﯐����̝���2)�DF�� =ٔĘ�;w�h� +��i���V8f��	����m�v��õ<�Dz����,��=�D3:�b�:?�� 4�R�,p�\��ym�17������h	Yn%�A%���Oܠ�=F�&`�������Hq=�������Y�^}��^�r�HwLͥ�ЍrV-R%1-��E���ax$8!H!DQ�#�AtCw�qa���C�?@��ѸRK��i/+�	�IK�M�7h���\u�[;��W�	l�l�5Rul*�j��l���[��i/ː!֯��(���@���Ϫ�S^��
g�&"��C���5QYV)˖��W_��:��G��$/j�k��pgs�ҙ�9�T������)oRQ]'��)F⒏'�-Bj�ަ]T��O��D�Z֎��ǩw��H$�32�����2a��q}i�M�Ï��I`7�TE�'' O� NY�$��%t[(�I��l� e1��2Z��ɪ%�o����O}�>ٶi��]����^����"�NRr	�����0�����k��^p�E�+�q@	��4�������H��*�9��%��]�wq�`�)�s���ĳG�:=x�P"�g�D�>�pw��1tQ��U��M] E��Ani	
��疸o�����+INI�TW���4m�>���1(a��"_��1���#����V�݄i�X���������R_۠%4:C��T��B�kAe,+-�ܧ�fI�Jwi�bmC����׿���r�u7��o͔�CG�Ν�{1�R��u$�A�"��2�y�y�8��)I4Z�d¨L�<U]4����2�ԓ��&r�h�B�������_�Z>޼C��Q�H)LD��E�s)J�$*U�}�%�j]3�����w]{o$�{�o�=//>��W߹)ߴǱn��ɔ%��]�,� P�7���˯Q���K��d;[%^HIy$/���W������\�JY���A�z���-�2��N�[G{k�Ew���c�M�o���[�6�p炜,��B��&i�77e�;v1g� �� Fţ������{��wپ����4�T�(�~z��?Ξ �(K#|��x��"#ŭ���s�gw�X��ڹ�A�����@�	����q�P�c���i���P��<x�.d,7ׅZ���k���&.��-��Ѷy�iҷ/ٹt���U"1W��k�^���Xf����9뜳�8�\r�6R�i��J��8< ���v��TQ/�	p�xQM�6-��B�#�f�����}�.�Tb񫲛i��X��W�G/;�S2�����WH�Pq�8(�m�B-M��7�	oU$a�ZW����Sn���H$�1w���S-��^�?����ܜoq���l�.�.�jm0m.
��~�����F��h��tIU\$���-d�a����N���_�E�J!�k ���cb�ϰ�M�a�&���?����=����:�&/�z�����T� Y��.�	��[)�4�a� ���!a#�S��k:�L4`h�����5ހ;h�AD^��8z��p0";٭�Y��+��@�[Ī�j�=ܛ�щ��}i���	�K��Ģ���q`/[�D���į�X^�j����~��օ��g=��~�Gd��aj�`�h�<-=��cɯ�,��	�(��2����j:;�c���EC�t���G���oI����O=�uG�_���2l�sK���w��԰Y�.\x�GMU����!���D;�yI�B��x�+ӥ,��>�e������9z���� y�%�܅u�v
�d�j	Q_�`1�BB�jr[4fJe�D��W�5�ﵓ�z���(w���swL�us�i�/��|��N�ߋZ!ސ:(�)Yј����JU�2R[����������}�(���Wɦ;U��X�0��)�d�
�-;Zt��W��r�m��	����P
����l8�D7��q�>�N����	j\�@ӛ��0s&��!R���O<�e�e�~�."�b���I��(��D�9=35���&}ֵ��a~gW �֟���"�=�|O%�D�����W�BD-58�f>�xu?8.�k>�H��+�) �h��ח��We5x'����6X� �I/�rn��|�罁��J.�����c�ƍ�D��K6m�"3T��H��.tq������(/׍���E*�˥���Y-8����lڲY��m2�e��m2�O?�Q3F��X�d0gry�'+e��_��TN�/�Hʪ�HG&�Q^��1�ѐ�9�"�Em}b='�꥚T�����w��[�y0������r�K?�H�G�CE�.����z!���d��R��Q�=��ڪrmSڿ�V�l\+����������Ӟ�l�ˀ$(��	��9��GA����W��j��d��N�+�M�v籨�R�)�����L����1܏p��z+D0둖����NU��)S����V%�����:cR�X)|��
�®�IdJ��M/$b�*aҶ7�+��E
��@������ll�ܘ�\�v��T� ���7tc�|�m%h�f�xU#+DD֯_'����/�!�s�9W]��+�Ue/O�J� (�c���oa���ձ_�|�f��f��
x@��$S�~VZ����G��<���o3d�p=ׯYҹL�I���2\p&k>������G%�>!�Q)lm�:K��3g�J��>ү�V-xD�I������2��KÀA2��Ғ.H1^)�D��eFJ��H���1b�y�W���IUE���v�<p��������tϟ���׿(wΘ}sa�ȣ)԰��m�i����0pyB��K�@���H-��荡�[�ˠ�}�e�f��X'�[��~#��_>B�����^��tg�f�A��e`ĵ�o.�	J��9}���4@�����^%M������\ %����P�Iz,����c��P���9Z�>0 ��r�q���'�$��}Rj���Q����pҭ�GD-�d�v�@�ݞ�5�Bѡ��摺�>=[�;��A����g\��@�,6l�F]��+�a��tݟ��`q���G
��rX%�RY  ����˵.F"aQ"���$F �X����ly2�ѝT�KŲ�mۢ��t�cQ���3f�}�{'����7��@W�@�F-p@����i����X[� 2l�`�� �9~GgJ�*��gΞ-�d�
������:�bA�u��$**�Ï��;Z��+Dʫ�� %)ED��&�Q�CAצ�T7�W�-t4�_���Ҳ:�^��Ӧ7����*E���1���/6PA1�� S�$~�bK1$�BQjD�"�f�~Μ~���{�k�k��Ό�������̜�˳�繯{�k]�Z�w�����3��p� �K����ko{��UO������
F3�])���ڿ���ތ��bza��ղd�hT%�Jں�Ƕ�+N?I=h�\����Q��`(���M��	���2��RYN}��r�1/�=ʟ�����#�hJ��j�5�`E��]�$�� Pz�a���B�G�*!�r��K���δj�rٸ�@�A��91P�7�٤ �M��1��.'��>#��{t��!z�8��B_(���� @ҫK����XĚ
��EknT��v�=�m�;��t1s�8�s�2	W�"�Y��_�V}f�?���?�[N���9��j�� 2 D  �O���駿\y��~�;r����^�r޳[~|�-r�QG*P����O>��МN�&|'"l��MTcZ#Q�;?��2�N&d����^���LM�J5�.-�OL�9��5_�d@�#�}m�p�Z8.[�FW��r�-�DFR�A���J��8Ӝ�%, eq��=ۉ���J��S�|�������+nY4@�������?{�����S���W��S�g.�Ȯ��>��w�.$���D���l��F5���f$-uy�Eo��ݛ垻n�=;7�I��3R�6��)_Ћ΃ݠR��7��Z�y�˶&vcx�[��m�� �1GK�N$��)OtǷ��f�ӕ��El�r�ڿ��iH+�����UÐ�����3�#�C�ݧ��@"��*nr������A�Һ��:���L���X�l��L9OC�֜�,�awS���T��T�	\��E
_����l����h`�
]�4B��Am�R��G?O��~���2��9K���3���)�DLd6np|.��\�W�M���G|r޴o%��|��&㐣�֮����eK��ɧ����I����[� &z~84F��+�����Ք:g=eD ���Z#�Wp�)�-�exlB2ټ6;����d��[dh�_V._�M��ЛuC��I�Z�C�|����j3��6�XSX;ve��I�aM�M������_�詯_��R����i�?�}_��n[T@��ݏ_SYb�k�$9>.cO>)�VL��ɤ�"��0RM���/t�0
>�d��wj�b %��gɣ�L���$�N2�FLKI'A�\�5�ۣ�ڹ�ו����/�,����۹�D�h3�;G����8�S�$�"�V�F��c#�UЭ
Prc� �b�3���j'H��Lz��cO�B��y>�э�]���Jd'�u�"+�ƤX,)�%,�REwz�s�V��� �&��c[6�T�w&�֝uŲ�&�L�׊1�<oh�2[�53��`�h҃�`1"��9>�'�n\p��ݡn%��뮻��:�����t5���|�����3�RZ��:��Y��{��vS�����l��7�r�<�Rq�)s�֭Ye�>�������P�HJ��o��m��Z�TEo}Y�7�I)�#-��<&Rk4��f��Jap��摧��f>Q���-���O�e`��N��>&)����Jur��'�����n_T@��ݏ��t�)]@����R@�7����
vy� ������&��<�����֧S�Y��T�1�/����ȅ�4�������ü}�s�o\J4�r$�%�1��;�x�4�b�wJ�ײ0BwN iJJRm�k2���Q��H�\_�76��Y@��3\V���z���}������7E���B���v�.&|R�zxo~�����f�m3}�Th���3t��N���.��S�!r����6�m�%,�X|�߇�¿��t���( �ٽK�>�(�y4��~�#���'�f8����h��~o���=���<��k�)�ʅ����']⸭��T���^��Y>�^k���}D,����p�S3219-�f[�ݱ[K�ZQ�f��kevrҬ>�?�JG=`��%9�#e�����d�ؐF;%mu�Kk�J�!-��$s9�I}zצ��;���P�x�'|���]��7�g���Q@ɷ�ꇒ��Y/nk!B�F&{�t��Hw+)T��ޮI:^�veF�9�e���!�����O<*���ǌ�L�,;a�#��>҄SO=Uo~�<��̀����Om�(�2��䣾����NY��,_�L�b@n��r�57��6w�oh�Y3��gXb�~۝
 �������I��A6�#ci��ͯ'S�͛����D<���8����M>�5ʥ�SaB��vQ�rn~�կ��ܸ�ƛ���
F�� �֮�_]��������_���y��� Ł^�ϗK�1�J����E�y��r�oQ75 �7^C��q��.l޲�5�߮R���c������)�G���x��G+�.���֨
�~���0�xGrT��-�3:,�:"�����nR���^���dr|T�l~JHO���!�����.�y��aI�l��V�~ KM5�&6F���J"�U@iΌ<|�q������E�P��2��(�ĆG�(�?�8Ky�(��'�Ճ�	s��7kEI!n��SN�VyZ����7a�9���z�#( TN��|��/�.7��T�#>?J��qDA$�o�v���|@!U`��FU�5 �    IDAT6]��Dw}눦d�h˴�K6HD�D(?���H ��*,�׽��w.�o|�[���º���<���-O�ւ��?�OC�����Up��9��:�v����}N�'��o���ZIJ���z����z�;)��Mo��y3"���Q-��w��:w��Ԥ00�@��
�s/T��L����shTW�k���$ AI�� ���g�,&��)��[AZ�z�T�����}��hVӖRIϣjE��0�.�56ⵜC���$��<5W�S�>"�Z��zRf�&��_�k�r�wh�����ƍ�뿧�g��F��N�y�	/�X� w�s�.Y-�8�cR�T)�xuG��[�]�(�<���O=��|�C���ʗo��_��k*K֝�0�k>� ����wd����P�q>�Ҭ���֮e��er���Ge���R��J���fZ�4�F�٢.bBGnln2�n��>�J���Ӛ�"��� D� �>�1?wW�sڼcm�(�< �S�E0B��W�z����?8�C�ǞօND��b�����|����*�56�G}Gi�+�+
6�|����m�v��"��%�a�������QG��hn����o}G�.�sQJZt��ӪzԽ/<�hm�c~�����G}T�ȼ�moӴ�ݗ\����s���ͦd�3T��erl\m�C�F�0��w&��H�Α����T%Rڴ�Ѯ����R�����S;�o��8�qL��s|���,�����XL��V�#t(�������Qהp�JJ�Y0�i��22�K7�F�J����]{�FY�~�<��V���dvP��;���6�����rT�H�(��,X=`6՟�xu�Wg���w������E�/���K��Ӈ�)/]w�tSP�tf>�t7�P��hSR��(Q��_��	qPJ��h�ʥc���%�j '+���̦_�����d�z��9$3Gbi�D�7�dv
L��
���`6Lz��D&�9���P���K��T�qDF��
h��  �3 ޓv����T��\R��K���=���𣺠XX�܈��{��=19�����Ew��Gh�r�����d��R��.�XG�#ԧ�87�t������p�K��sΗ���m�j��� �����|����O|��Kgtǆd�[X�5۟����]Z�¼����/XD������zL�H��o�V�hDM�v����06
"��w����_ܫQͮ�=����ܠR��y��r>į3��X4B�#�|��pI �@�Yy�O����{�/���)�w�Pҽ��9F=��rJ�����P���L��)uV�\&G��E�ctB6=�E�w�M%���IPv���N���R�{H�T>/�|R����<�������}�(_�得~�.�P^6հ�32�с���&V��?�5>z�Q]��<�6е��B-��FU
��J�r�����9���?��[��,�KkY-U@�^�<����pSr�l4!S`��C�yl��-(�/B�L���SZZIA�Ů��K�4 J@��4���5��5O����7��%����8yh΢�.Y>��c_�`ō�a�Ar�UWɶ��T�R���4 6���R���g��+��Eğ#?Z�;�ղb���W���o|MS$F�)m���U7b�LG*�f����d:���⃳������ ��z���d�����/��q�F)|�M7ݤ���Oc�R��|�-V<~�	嗼j�����׋���Y:jל?J�2���D�����p�*]�2�_�B߀�Vj2<2*��V���Gݤ�2��9�~8Q�v��g�u�����&�l�<��6)��RA,��K�
g��@��F̿P��ds	I5��;����K���E���x�˾��Ǯi�X��a�]͚Jq�v�ԭ̛� P�|u_Mz��6�CO<.o��M�wr��K�4.{v<+۶<)�vSg�R��2�K�:������9ph�;�� j�c",�Vz����*<� -����皖��ߗ׿�톽����m�xV�Z�88ޮmd��� ��ǂ����ŋo��g���Iyzz�(�\r���0[4i�/x0����ϧe��m���FDp}��3ΒK�t�k?�9�T���5�@IK�!�'
��8�+��h;v�R���7����Wwh�s�35=!�s�|��Sw|�"`@N��0ђu&�ߗ4�ꫯօ���i�Mw�|��+��y��`o~�^����V��0���Ьח��P������M�����#{��b3����b�rr^���d��i�Ѹ�+�SoJ�m;!l<D��A6=��l�=!�WK����zz(뽊+��P�UlF�j#"�̜W6&B1@����ӎ{���s��(_�道�՗����RM����}���69077(�ʂ<����"0'�D_mĞl�$�d�OB���s��)w�v�|���E��������L9b�HX̢f��Щ���8���X�פ����/���*��]�ͨ���c�Ѧ7F/���(���P�eO65m������X��0N���n|��kV�4@0��x�q�a�5<��c�O}Z#3*0�ʥ�y�r��}�1C"洜}��r�aG��G>_S����rd�I'�T��]8�"d�ܢ�`�: ��c���#u�C���ܹ[�\5�e��B��`����V��>�+?��g�*�� j�h	��}^�p5/'��?�s��6.��Z����j�_�kEĭ	�h&�Ro���'l��23��ONͨD=׎j��=������-����p��@"�t6'�zK����#�>F���-��Kap�4c))7��^}gq��mK�;�µ@ʃ��q&�Tk��s�8�=W���ŋP���ޓ���ǯ��8�D �*��̶m
(qNr I����)�p���xhʍ�M�X+6�R����[%g�r�ԋ�r�ߑ�̘d3�9�$�*W�6�q�j�D��"�4��3�����<��J�oN4�F\��j7'Di�dY� 
�����0�$<'�x����5G&R�����p��m��X��쐣c{��|��giiuժ5��O~J�.Y��Y�8���ĄVy�A}��GĆ�ʳ�n���{Q�AY�5�灌�d̉�B��=˱`#�	�����wg7%}y����xy�8R�LJ6o}V��'�@�
��N8h��*�c���"���y��'I��TJ2�T�*�VK�r��m��g��6՛B���z���6�yl�ᆾ/�WBO����ާ�	ה�����I�R��)ך�ʻ`O��ȣ�`�ɧ�H'��|�R�)�$��)�K�Xjaa�o �vT[搲�����E�1u�g���޵�)��~t�)�|�#��Wn8aO��J�aG۶I����b�0: �z���
��Z	
B�;x��H���:ެJ�4%׭��V-�鱝21�[vn߬u�t�]��?�,���4�� ���-�F,�*~�έ�Oz��u��7��H宻�Д�4���Q]��1�0�����{k��oq�����^�B�	ݱ�>�tM�����W�zH����^>��+,�_�Wz����K;�/��RM1�xO�ح���NU��
~�ͺr�)v������g�5(�/��C����x����9�ߓ�N;]�O�r�@=*�^"R���(��5�y|?"΁��y��>>���k,pצ8��U��E/�>v�$���ư���q��s "��As���_�����~&��Y��l��p�R�X*��GW���
Kdӓ���1[��!�JJ�͇j!��DmB°�xP�� ��܊�=�}OIFǝ�$Q����ӎϢr(�~��S���'�i�<�� 
Jk�N)��!YH"��1@�>�H�ξ��s���Mk:�N��ѫ@CayVRL�����n��O:N�3crݿCvo�*��KBw��%]��Ee�r�	��;��ʩ 2^:dqD��'nh��wq@�e����f�x/zǟ�Bd�d�r�-"nL��eޚBv�ѵ��4=��|����`�n\9���+u��?�c-ۢ����'�@c�������p�x�u�qK�
��_.��z��\��^{����!�h���vBu0�2:2���3���|�_����6�MMN1����Fj\��|�����Q�������%�຺���	P��J#�Px9_yLt�)����s��,c0�݂W� %�����uS��\g�'���]aA��?z��5h5.�z����P�|A*՚
�Z1�il�%k��M�l��JK��>�-մ�S��"��6
g�QJ�m�q �.4��d^/ I�4�(��k�8���wQ��7������k+�?Zih�RۺU%ߎk7q�� (�V���d_�B�,�F�r��ZU.**�'�=�i�5f��#��v�o}B��=z��hC�|z���sp1/�~��E�r-˩�s(��F�%����)}�S(o�k���+_)o~�U���S�k����� 
�\J�~�u������Z���`����GUG���-���vꎉN��|���P���taI��F+i`FS'ߏ���.�իVis75|������M�f�X&���������D.=C����WV��P9k�f� ���qM!p9���_������NA*�q����|�����/��Y:R �P ��kj��Y��?D'޻�)������h���lv6p���lrtD��\��������VG�mO*��R]�6t�,Y�J�ܶS�gj��(���h��3~��,�J�@F�c7@Aj�$��Y���[��N�� ��w?vu4Bq@!Bq@a��:X���@�Q� �)LT� �T�T�I%���{�c��ɫ�|��q��������٢a�G̃a7q��?7 ���DoPnnZ �ŉҹz������
��\��ݕ��vl�

|�֭������
�]���%��X ����Ж�����Q�V�
�eF�2��J��rQ�Q����^n~�#"�C�(##��L�|�
y�ٯ�����* k�s���8[	���������y�MIj��1�+aݷ���:���Ԉ�>���kDH���?�I�܅F&�v�@��M�j�R��+4�����H�H��r8/�8�� :J�|�e+L���e�}J��Εd��	���0�zz�u%�!2D�H�^ �oX���LOM�ʥCz�\��̢�m�|�%�[hW1�9S���!�$���J���I��4I��yi�������6γMt��:`�CQ��(7t(��J��#��{�?���My<Bi�:��=��MKyf��r���-i7l�������bv�� �`��ĩ�p�g�R.��4�Kj��d�@F�8�x�̌�0����.��7�!��� �M+�f��c����Ut6/�e>��Kznn��cᐃ��+f���:��/|�.ʮ?�hW%j�(��)y���\SJ��w��EJ�
$�֩k÷����槜�f����j�>K��F��Ri�Ǭ�N�)�V��t����}L��ܽ�k$�o/-�f�0�� *<:�-���~��_�ȁj�}�ޯ|����Xh��ߘ(���_%g�y���{d��嚚�~�� �Z��;DwVV�����f&q�yp� d�RoYP�Sۦ�M͘�hhYHr ���q�?�|F�o�&�����fh`P�S_*m,�-�v���&H�/Y.�<��m��H'��F<���x3kld.��oF E�b��� E��DO�gH�T��?!9�$X��^�k�l|��]{ǯ�n��p�L�#�f]�۷Kq����p��A��8���,��]���M\v}�>�>�����|̪�ui|X:���s�r��k�G�G~���X=�ۥ�usW�{������)9���U+B_i������S%���T*�G4�i�id/ �����W��$-FAp*욌��I>�����؝�&'t�������9c!;��;k�&^��r��5�:�E/��n��\z��4Bpu)����E00���t����7ّ��r�M��>��
��V�%+Tk���ԦB�/��w�� ������T�F�k:���O��~k��q'�X�wđ�{�����۶��M��^�(^�u���?8/�tIZ�9k�psq���ʺ�'�&&�ebbRg�T*Uټu��ھ����@zO�G	�m F�O�@����0՛uI啄mX��`;dQ��q4v�BTҭkh7g�7�?�z�$��K'��$��BF�ő_��	��w�r_�����o��響����+8�X�H��P@��e�Б�2؝&�s�x�V��;�8�̛<H��ika���JyZ����k%i��rܱ/�#�(�;��خ�4��xL[�)g���ꣀ��+��4�U��rJ��B9��b<7*�÷$ʣh�i�$d�R�-:Ә��V=jV�]�*X L��3��>9���˺u�ˍ7�P��Ƨ&M^6�\zkX.�b�Y����W�"?����=|��_��B����� K�����4�>'ޛ�f���k���2�(����\��w>�Re���d�9MŖ/1�������g�����7T d?_J"M
U�sU+� u���/8�sL<�G:�Toa7X�~��	�P6������8�:�;��$U�� �$���D|�n�֝	ŽE�H.߯�+�1^_A+lc�����R�x��ҊɃ�>%�l���)��3'k����JP0%3'g�N
���Hq��Zl@�������_�\�����tef�N�0�D]�j]@�[H������p�":6���A�=�ꬖ�+�3��B&#���r��e�SO�o~�KɧbҗOK�XTn@��P�g_e��Y���6lԅ����7��b,H�+B�2\�`�k,�𔂛��A.�]�Z?�������U��O���IU���f�I�;��K�&�c��4��׿�����VHvoA��J�C*q�E���k��Z��uh,@�X	����W����K��\�=:,yͩ����sϽ�P��ɇN�G�~hoL�Q�6��U��}�`1����A_��%�X������x��*�A�kK ��e��0��h@x�TT q_x)���1����+�A&����X�#�2|L[mK�]���!��e�Զݲ}ϸ�X)��o��!{�Zr�k�3]�� jl�z�&SZ����
�|�G�8�+w?vUmɺ)�t�!By.�(W�;D(~B~[���u����U+E�ϥ�^.J�<��˗�==9%����#�u�-��~&�zQ�����b���@��s����gT`�=�pU-)���~�G�Y/U�����/BnnPn2U`v:2[���K�/ӛ���qlT��,��!� ,���oʕW~L�y�gT��AZ������V�����)w�u�J׵�����	`�!P�R����Q�,�?H�8O�g&'4� �p�#�"��淿��B;��^%Z=�L�ꑡ3U^�y4���$OO�{���G�+;�J�E��)���s]٬՟��%{EK49m��j\=3�i�G<v��3�,pmy.�9�?h�t��,]!k�;@2}C����st\���O��iv�����p��ݜ烊]k{�G((4-B�$s}2ؗ�Nq���8Ὃ�����������T�־%�jHc���5P�Hy4B�ϡ����f>�(K��$���A{�C?�|F��R���l:.K���o�>ٺ�Yyݹg�������O~Xv>�����0�Eo<"+��k���9�bDt9�<�(���.�U����o�щ~��lGp"�sq������	-�5�1�\�,�)	�;����Iu�#�X�l�\w�w����Ko~<QX�ʀ�7>��s�.0̨�s�O�c)�&�|?_<,$R��~��]������=U+���+�>[�.�����s�g���R���#�A�PP�T�_�,t��Q�ڍ�#u#�X���a��up���
i����.}_�*�Ĭ�05�1@��M���"J$:���1��
����q\��+��O���:�z�Q�|�:yb�Vٶ{Tb�d�dr�,�l��qƣ��w�P4zv���&�B�C�F�C4KN�c/    IDAT�BR:���;��K���E�P�憻�����>SXs4��hԤI�g�NF�)&�C��PxWo�6�]�k��D$D+ũqɤ:�'o��g�-M*S#r���%���˓���'e|d����p�NL����7\�>���`����ݞ�����Ds�Jш�i�d�c��l,��(�{M|�:������g����a�h�V�K&�>�i��u9��s���F;�K$��ýV)@�P���D3.p��g�%}-�ƕ�|�!5:�ԓ5��pe��?��}��&���t���@�Et��뾫��)�sz����pi���*�æ��D �	eCj�s���S8���R�cn�@��_���K����LMN��6�3�����F	`4S����Hgrz_��M��Ɇ���k��cO<#[w�H�0 ��A���.e���
\�>Qe0�K$Bᜆ��LH,��T�`�2=��W�v�%�
(�����iק���?�B�-��7G��7
�����>qP�;��L���:S���ai��n���C2�t���VM�؎�ڕ��?%�mX+�,�G~�+�
P�����n(6�z�.��X\(�d���Й�I����=��o���]����y��r�����E8T��l�"vF>�+)z3�F<H݉:�dzjJ�g��#��z�`�t�7�� 
  p衇k�-�=�R�F�](�vk_S�ry���Y,����!5b�җ��i��8�t�ح�?�蜫��K�mߵJl<���|+��*h�}Q򅈏�ёU���r�q�t��~�OT��F�r
~�����0��3�g\�pZ�'!*�z��)�<��;��m�<� �h>�T��t�,�W���O8IrCK䱧��S���$��)�K�#2[�J�����q*R�J�F&�M=BA��@ɧ�3�������~b1#�����57<2������(�zuN�⤬.t��a7�S2'�?�O�.���S�;	���:s�n��J85� %�Y�b����4![�U���nɧ:ҟ9�äZ���۶�t9no���G��qv�.x��	9��Iy�lU�܊jY��`1z��y"������%eW:q�������@y�)�YEݹ1/ڵ{���-o�����8o!���a!�����*�  ݭ���s�T��NL����I�d�ũY� ,>f���`�s�Cd����j#ODHy|�h���aQ����ND���^tz�VY��
�ϙ�����q5�V��i�s�i0�сu�ۣK#�-=�h-�<�G�7"q�4��.�d��H<��Z��Ǆ��k�+����}=����csA�mΌ ��$3��듁 (���K>}�����~;������u���M�?^\{�
���83�\\�d$;F�y���"7`r`�(p$�.���X��U�٤%�zU�>+V,��U�hq���i�%%M��J��XK��N�N�G�LWk7q�V�=�L�7���	�����Í���*eeP%�� 'zSZڳa�8�w0݃- 8�hCw����������(HL/��
R���
D �0Tph�gA�jq�(J�Q�VM<Jbx�N����o����[9�IG^�r�еbŀ.�l������� ���:hW��w�D�E��	9���f�� 	���r�;ۓ����q����6U.s�\�=c��t��K"A�����k���ݧ��,��r'�Q/8F���#�=�E�ز]�V�U�;l��9�	�]W@�^�9�s(�Q�x� %��Ɋ%}R���O/8��KP�����@Xs�B��U��,�N��Q������v!@хHͽ�����hw�\������
u���F+���jV%o�@��5����)i5*������*P���ȯi#�a. Aʡf:a�qS�۫�j���jC�I��.���-UI��-7O�����S��f�H������!��#b�E���-/�ص'D3V��R�&ܹ��.y��f@/�~n0����Y�A8@Xdj��õ�i>�8�]j8�&"0��TC��*��ϐ��o�����l{��4ܒ�9*@�@�����g���X�H� P�	)���>Ou��f��������1���䨣���bY6o�%c3ei%2�=�pMm��d�G��O�E��>���}&����M�6# ���H"����9i�o���SN��o>����]u��o��G�?ZZ{�t�R"��]��`�Jq��6#�ڪ��"Ch��&�] R�l�(�j�(<�˜��l�1�20hz�>L�#"A�(OK�Y�L�)if����靛!�3��n��>£vhg���Z�q̴+��5�51&bP6��=��J� Ðq���*N�.���V^݌JT�#�/d'y.���	���\W�v#��T8��B�x�ԍd��!���;y�]�)�>=�l�>	���}]��z%l�cX�k�����d���۔�P-H�j9��"B*P|<���{�q�\��͍��>\��!O�<���e)��7�%2��cDhY�N:'�LA�D#|g�l(��}�w�sS����E�O�����~��`��\��|RR��~��߷������7l���� �];ev�I(�1P�7�����r�v���4j(˗�Ώ_i�&�!�/��h��Mj*Ԙ��NuV2����^�.�/Lʅ,Ho���hE+@��G�rl�Ȕ�k��47;��k��G(�9+:�ϸ����P�`)����^��������T���X�i�m�M����:��iY��F h=%�S�L�x|A�&](|�WN<r�o�N�s܅�p4�ca��&l�z���ߖb2ͱ�%�=���)���^%nՈ�ݞ��M$5��\�]�d���`Kkq��R~��2:{�OK�͐��@6�N�w����T'D�4]z�B����BA-Ke)��H�S������g���oxd�G�Ckה���P������$�%D*~ºш/�y��͍ol��a�{����P�J����H_�`�N�����\J�ͪTfƤU*J�S���=����H�(<|V�e�4Z3!��&>�<���x~�7y*�ъ��^�����5����M�)&;zx��g�H]ߙ���T�S!~�^0.kiG���pεd�FEaƜԇ�-����h�{N�B�v]�U=�L�F((�i�$(�)���Դ��a�m
��~��|�Q�q͌V�H�ꗔ����HXl!ܘ)�xɈmQ
§��cDI�I�\��WH�RYi�1���az�pMY9!��w��B�Z�\���Ţ��F��P��6@ɦ�R���z���}��w/){��n���P���R�'���2�S�='�+�D����Xy��uZj}W��H�ZQ�Z���u�Ե�W ��j�>6^�EU�V$�iI6%��H�^�ziZӠ�ԕ�u p����1�����/(�V��n z��#6��K��U /G:ɫ�dB�+�� �#݈#tb���.�i^�����;u��EH����l>����� ��/����K:It��i�}o�G<��c�=�eJ.�2�}?�g��	@�;@J��Հ[�� �ws�[mʥ��6er���}:�	���T�jX�zJ��h�B�A'/�p%!�XV�	�^m�$��o�֤����c�I�QnP����\�IwtS\@Ԧk'T�0��h�M�A*#\�Sm�5g�|�K���O��O�˥���6~�;���?Ք��}J4Bћ*����":�0�f�6�h��hň���sz�,!��
� �`T��zKCW����` (�X՛�5jҮW%��I?�3���I�ʄ$ڶ�F�
׮�snP�-��@�q���P���k���.��]��[#��?��j�����la�����:w����;���H��Q0EJ�� �������+��KE��w8^h/{{T�י��n�D�ܮ��5j���K���£Fԩ�'`��m�n]�QI��z��-e��T1@��<m60�O�MG�0�#eҌ%��	����ĉH�U�S�7�]�^����h��4ۢ���/����(J9���O� �'3��夐IH�2v�k�:��{��~���r�#�?Z[�ߡӵ��kui�ڮ��<��T`P�<<��#����:mZ��B�y�9�c�i	O���*��UK�/�KΊ}"�ۜ��������OCMJ�,�������4fG$�4�;@E%�Ϥ`�x�fӤ�z��\�(g�I6Z�|�u�M�H�A�����`mݴ��IoJ����S�n"�:�Ee��tG�r_�KE��d� c*G��a�S{�~�Z`�>� Baav�����0]R��Xt�49ΜO]��t���L���l�w���=*�.�z�������Z��!��SB�o���f�D�A�0cI�^Ɨ FSy��{-*��0@II3��������������ij8%���cDb\����m�����;A
�`������=���݃��
H��du {_.)2��'ox�����oxx� ���x����?R�_s�L�-IB�훥4�[O#��j������<��&�z��QwɧH˿#�[;(����py,
�2��͖�)(��\�T걎��9J��Z����<t��r*$"<%|M�ҨU%��k��C���.i��S���nOuڒ�7-��([[�C�QǪ0>윶w-�v�����
�*\{~��E8AQ�0+˼ ��(�R���t��(Qʢ$�X�.\�2f$ޞs�ݻ���<�������P�w�<l�x��*W~��| e�"��b1Z�un�R7U�Z�&-l"<2�����,��=d���^�R�"t���.u�G36�Q�A�:�ՆD\uUD}q�ē
��#I�ubLݖN"��)$��U4V(׫on��]n0��x�����5)�Zd�������^���l,<O�& �FMa��B�й���Md�Hk�3�M������_���\��E��G>Z\s�t��iAc׳Rڽ�(j����z�c��[�2bh@�#�9��+����m7$Ŕ�RIZ���X��R�("�DZj�PIIe3!�F*���b)��d8DV�V]�[�Jj3ckVU�o�$�(J�^iV%�i�3��.<. �<δB�֚��M�|��<g���Xd��#?ݔ hh�g�n�~�[�W��Ԫ*�P����M4�.N��X����^���Wx>���l�j)��@���K��[&:=��t�[ʸp#z�k����}J�u�T�K��k�x`[�p�KP����4b�� J®�0�/��;8�;k��rI�t|�t��p�=�{J���N`K��<�K
���A��(�.ġ����+���X���
u�l�_��q�O���g�򁏽�M���\}�]o�~�������������)������H�XG6��[Xv�ٯ�����j�?L��m������xG�,��Ĥ�ԝefF[���DP ��P�9���bm�4�:N�!�8��QZ�3{��{͈��Jt$������z��L����Ԭ�xء<U�4��7����f�G�C�i�;����W�<�,U�ҽg�%�s�.
(~���6�
D���̏�uJ� TRz��k�������m��g�0f���ֺ>��������y������9�)Ǉm�FlY�b�Ip�P4XHH[��c�4��t'��J���J;��4��9�#B�ʳ�A�� e�����ni)kT���s�'���["+�&n`�m� J'�\a@
i�ħFn{��'/2�\��o���J�ڍS����t��⮝
�� (���_��y�歷R~���s\Uk���4k5�R����G(��K3N��V�fu�(�JY��R��J�B���u ��"��Z5Et��#ٸ{N�U�*P�Y���4�ng:�ӡ�������uG��k�PC�no��p@"�\`�ɭ;aX�������^��ש� U"n��$p��|����/��9�@q���?/-X��=�oX��A��|�����hEqL�꧞~�+���_�$#�)-0Cް�@=߹^DQzO�I�َ!a���nє�o�C<Y}x��o$�\oH��ѪI<�ը�'"KH�Փ�ր��`T�o�U�1x����o-���.��/����F(��C�����-13��7�{��|�7��\�wWy����?�ަ���8]e�fX��ٽ]IY���{���q	("]Na����P�Ŧ�E�M��ToJ�8�)O'ޒ��+��I��V�tezV��J��S��Cb�-B@���?�F�f-#��P"a"JIt�Z�IƚR/O������u��Ue"�yK�1�A�R�vLՑ ��E?�*I]�!�2��FZ���`;��d)�ld ���ë:J�&��,��e�����=����c����y3~�Q��luAB��Ǐ0��1BBs��7�=?][p�F �C�H�̳�"Kݹ-Uմ�ʝ���T�o�ZR����H������5�6�*Xc�y�,�Z���������?�4�3u��s��r]�9/�r>���XW��R�Ɖ�J!�Jc�\��3>�޷���E�����w�����k6���FMdx����\o.����9��)֋9"�N4��2�^�����"}5
8Z�kH�ْ��rQ�	R��J`�Ӓ\2+�k2��$Y���������0�������j�����M0���1��.�zIZՒ�*�����h��%�V�ᵂ�����B��BP����:����2��9���?R���pO9����zV�>�B�P�&��E��@��?��iJ��8��e�hy���W���xd��;�� �L
�n�E8�T��� s����^$���	 1'8�4��*�l!���p_(�ɵc@W2�Q@�z�0�>-Z$M�]A�-='I�����ӁD�o?�y��s�Y�Ȱ�������c�)���C%J?>D�<[7� x˧:�lu��?yùx��_�������?�����͹��A#�o(��^PZ:�r�^_�Vw�������}}�h���`�!���hImfZ����C�VH+�0@aמ��rqV�=P4Bi�|��Tkhl2�"a ��R�6�e"����-ɤ:�iT�C�3 ۨH@�¶]��g��6%<�Q8G��b�b�A����V� 6WR��7+')��:c.�z���)��+��+E�,<�A�A&�Ob���u�(�F!���*���}|�)��<�Ng��g��9�[)�%��v�u7��ߎ.Zw >vEW9��3�RϽ���H�t�-��N2��q���MH�X�J�&q %��N*)u�� stI�m���`��t��< >S��tA����g��hE5�Z������,�#O��X+[��o~�����ӟX<@�������F�(���o�RW@i����.A�p�Zx}�,-�\��2v��>z��P��F ��U�ZIA�!B���z�������NƥVe�gP�0 ���$��I�I	�d-!������lL$Դ�o:��Itg�%�_M'ERx�2�2�U!��
q|Vl�5|���X��<B�� F���f�)5�<��Rb���S�6��$`�z&r�܅���B;�x�9ʩxD��J4J��Q�3���G>�ӄGE�e.��(��͙��|��Io��]
����%i��\J��ab�vǣx%E�\g����詬���7A'�8�D'���_��Sz_�RIi�@�FM�,�\ʺt 녪է����o� g�{����iJe@���"@�<�l^r�v3W����o>��E�k�������Q�[�nO�,�f[�{vHut��è>��4QR��!}�#h
����h��#?��J��B���@%tP���LI�X҅K�B�Y.�tj

��d�ri'RS��j�o����C(������z�$�m�/��zPfnT%^+I��aJ:^���3�ER���Z��h�]w���C���~t�)'�B��-HK�A��=A:�&X�$ՙ���    IDAT�����$џy���G"������G���:v��Pn�ffV�Hg0��X9�#Z�`�y���L���P4#u�AP��\�+���l�#6�z|����(D�����6�ҡ��OFS�/u⺉�bq)�0q�"���9i�Ρei\��t��@�PD⺑���(�Cq]
ϛ�;1}JW�bm`lK��O{S�-SJꍁ���oݫ.����-^�s��?}���_Q�[�@I����@^i_M��wS}#�Hy�%Z~���jĮUK���o�X[�D-L��o����q�ޒl*+թY�g�-_�`��J��`�tX\(�7��O��w��D0�	ߟ��!�q.	&+��4��P��$��I�0�h�A�9��h�He�q�%E7j݆�+�@�)��h�X�zRfC�����p���(�D_��>��(��8�^/�K��7�E�_�N��?3�^�sT<P�X=��r?Q����]k�h4����G�SYvx��[�hv�J�8��X:/�L^b��	��B�1�hK�XҮv�@�ުk�:}#шe-&��H8��t3T4�܀���ޢ������ 9�{��/��t���ߘ��oXd@���?}���طz�x��G�wIulXwo�& U����޼�go��?
S�JR�Z�k�n�L�-�k��r���k�I�oR���j���a`���MH8m�K�Ρ�C=��Xs ��;�Y삚��;�L�/��5��Q�V��"�VE2�h'��0Q�*.\dҒٜ�k� ����*6v�z=;�����%2�.t^��ht{�#�]4"%L}�p����EmQE�;���G���CO���B`��/)s���x4���9�
}Itsn���mВ����V�Iz	�<"U���Jf$�T@��h	=5Ze�
e�`4��e%��N�'�ԅ��Q�ߦ�>���� '
&{�y��a�$�N������iI��\m�?{���-j�����|�OM_1�_�f�ސ�谔G���ꀢ;"�pFo$o
{�s[D���_�m�=D��@�оݒ,�,�8��.r��D(T;С����^�'�%˖I�D/|��u��J���ӧ��z$�4=��ҋfR}&c [I���a�v�(�FEҝ��Z2i����Y���6�m� ������!��m��^/�Ev���gg45������ �׽�#}<<�u4��1\�p=���F?�>��d~�]޴�{�/���ͼ���t�&�Z�b�>��$=W6���/�܉Vw���[��e�Ev`P���J��|�ԄG���F'�?��4��Si�(�\�6�GϚ� Q@�꯺��5���B�����p��K"����$�P�ty��w]���/>oS�O~�Ko�R�\�j]�26"���(a)
(za	�C��|`�݄s:�<�5�Z�t�SS erZ�D)��,�o�tRt�vTc���6sp���
(�)��t��Pt���s�3L������|p[ic�5���V�q��YUܪ�%ё��9��(�]@5(
�?�0t��s#_��5�Z8�o�9��}�o��\��_� .@ѿ صsr��鋝=O��ל��q9��O���W�}<���f���9���ר�%_�,::x|�R�Bߐ������T�T�J�єF����/Jf`P�M"��h�GJ)�IC�o�Lḟg�k�,�<�+�Y�~�.����Bk ���h?Z����}J�zo�&��.B���\V2�z#>���_��?���'-N�����>�;�s󳥿��-[;]�H�t� %X7�pm��ڛ��L��P���C��4R���n�9�@�6E*�R��V X��j%�~a�S���ٙ)�)��X)�ɨ��,��R��|��n���:������C}D�����:������g
�հV]-�RJ3�R+NI<��1�����T��:�]��Tس�){PhJt9?�՜��J�Ѵ�ӈ(��L����n�}=� ��9 �)<�W��| ��7Q�5
b��Z�*�v�ԅ�H���#����Y5���bz�$3e|t�nf�4�܈A9��v�:��U��@	��+`1���Sb�=[��?���su3s��}5!�Ϣ�p���������_�SM�-b�O�Ca�2�Ҟ�y�e����/z�"
����ny������u3�Ju|�M�W; �Y�����7�F,a������O�{��M�"���JO��J �t�#��Im����[�����ٜ
cIy�kVI�f=@��6Q��<�j�����5�T1�Q/]����w�{iT�.ɦB�x!�P[���3c2�s��ebhd ���A�L5.Zo6d�t%lt�bM�Q��|Q����o�]��� �bunZ��̲��+OU���(�#�\��;��s��<="r����g�%G��Er�n�J#.�׮Wk�]{�d�������r�T@aAIM
c!�������%�2�lP�v���?\��T��s��G�3b�i�WR�M��	��&�����PL�c��T@�&���֛?�޷^��E�o�z񏷗��J-���f�,��a���ހ�c��E�s��g@��)�WZBD�-/�+���� Ȱ�M�i4�6=#�bQ��кU��C���:5%Sc���ʵk�c!U�!��PȌG�d+��{�x���\���Ïپ_��u=i���il�x�9�U�&:�,���䈬�OJer���O˖'���9`�A����
OtR���0j��`i��-�hw7�7��a�L�ݰ�D+A���k��+>�߯�q<��ƴ�7v#�TB}{4��:�x4✇�䵛?tܪ
4�����HN�fC;���Tj5���y٩�I&-r��-?��]����ex|Z�-���I�D�j�HtҧC�qUӲ2s��UiI���VIǏ�����I�?��E6��%́����P���9�U��ȿ�I"�K�b̏�<e���֑��P���h��ό�WA��7,�K4��=����K.\\@�����������rߺ�S�����&F�69�l7b,��!��$a��AP�F��f;ض�7D7��H���|��I���<I�i��ukj-�ӐL�!��q)3�/����+G�p
@i�ebx�J��쿿��j�7H
��]�CX�-������0\�ܶX���eV���R���Z��=�袮k�a[rɸ�*�2�K�1)���K�'�����_ʲ�+etrZ�i�sxs�Y��;e�XS�-ƇX��Ld%�Ȩ�m�©7�Ro��H���7V]j�$�*���:��Z."���2�j�TEm;�w�B���P�Ng͵�|T�Z�y�1FCg���P6�6�3�ѯM�0�����P"��1�}')R�T%�K��O��m�U,	@-z�3,S��f�ToH>���̬\��?��}��ZD�&�W~F��Z��<�c�T;1������H.ߧ�P��*�T�u�R�f�R�#^9����~�
� �⛻��R�&ӝ�g>%a�8��{�ڜ�X��¼.}�؂ߋ����y�|��0�P��d�Z���|���������v�O����RvՁS�����a�NM��+�H
@�m ��u��U��u�0����v'9iu#�D�0�dj��ְ����@/X�,5Z�K�]1@���\v���¸řJQ�i�e|d�*b׮_�H:�׷�Y���u�:7��ߡ��Xz˺eq�s�T��*H�8%�����XFg�����^��I��Ϳ��^|�|��k$����V����VV﷿�Tk��ȳ[wH�і|:#+�i�3�B�dG���4k����x�Q֮�D��Qa��1m:;+����d�w&��Z�s���h��+`�&(�u.4ig����J�i?�zR��J��7���\��?��dDE�^V~�88D`L�3��g�34�Z�^����v"�����Ȉ
��9�y�I'�����ƞ�=����d�����l�.��\)���=�>$�t�T$)�LX�+H�0(��~+��;Rk�aۑd[��H�R��RI���	�uԦU5>�
��H�#���W(�F�!���������Z�E'suBڗ��S^6�I�S�j�3��r���<����?��ُs+6��ÎҘ�#Չ	�YѨ�Uص�;ӐS�t̠�ݹ������n�����)~��ry�c)�Ms\<�^{z���l�&�Q)OM���jI�s�.� m'Bi�S� (D(�6��a��.��y�'�rvK�x��{k~�@d���
�*}y�\*!�"�׸�\t�W�!KrY9`��<�˻�m�{��.Ծ˿�_�O��g�#���-k7��v3Ɍ̎����]җf�PI��T&�͏�	��d�I���%r����Ò��\!Ⱥ�mS�f/����g�&XQ��K:�Qє���޲��QwE 	a!s��i��l�;c(lkS*�������|�|�gf�Ht���;��q�a�q�F�~���C=B
�Y�TERI���N�͗�MY�b�������;�����KK���²��楙����D�"�\,-�FM��I�TKZv�>-IߒA�, Ku�'R�� &1�P��9{0қK���މ��U�}��.�?�.k��c�NeP&��r�P�wכ~���_�d��́�ό����t�(R�oV�vOO$�!���*EM�R�s4|5	�S�6���\k��@&/�B��{��RQ�t���/d^-U�vP�(�LMi���I;��b�,$�3%��cZ��z�z<���(�̏P�ɪK�*���J�`�U�S�I}vBZ�qi7+2X�[w�jU�]��d�)�>�I>�������V�����\�_�u�*����kerzVV-[.�xBvn~Jҝ�4E�f�b��T2����NCo"̥�(hCP�0�i�q	ͧ1
�_�K[R�F��)u$R��hR�j"+�'�)#*� T�i9�E��H=K�r��T[k�CTƭ�G��!��ش:�l��@!)c���?�#��%�4�<Z��I��I.��DtéW�˧d�&�g�����ֻe`�:�6�Z!�%t�'�B�C~,!y*:Ū�g��T/J��$�o`@�u�"eL���'90��<]n�uV������ou8q�r�m72���$ec���@:��a��[�V�o�������o;�'�������K�������[���D1��8ʚ Jib\%Mʂ193eNv�rQsY�4�����b�R�S�5��j��(g���D2����2}C}�.�Z�d����h14�,%��Q�H��xR�Nq, ��T�ƥ49�'
@a2Z�Q���
(ơ��?ig�
(5zfԹ�"�^���u#{ٶ��y@';����r�ZQv��y�K_(G�Ff&�H*��_=�k�t���	�f����@�=�\�h�W�|I�����К$�|��:�@����ﰢ��ѭ[�4>"+W���J�����bY�ek��V��2	i�+�i�dI_Nr���鎕V���q�rEE^�r�`�Ig���43�
�E��hV�1MG�U=�T"��nH�>dJ9Z0SX��P����g\O���zC9���!I$$�[)K���L�)��=-�;�,yۛ� �tB��Yɥs
̴X�ci��	�B��Hs�l۹M���o����)��d��H�����Ǭ',&���+W�51#�bQJx�fRjQ�����9"�S��s�#�J�J��k��9�`O�o��rx��F��{[����r��l�j,�1��j�Eʳ�������W�8:��߹���<=��r~ա 
JA �:=e��Ij24���;���ѿҮ�jũ������fes_&�c��~:�ˌ�[���N�c�G'�mz��cF�ˇ,[��ɪ�Xzy'��O���	�Ն=��I���v��d�5�OO(�h%g�AK��Ԭi�Ҙ����#�����2ii$
(p(X�iI��u�aH��Z�H�ǋ]lS��{�p "��6��r����W�K�[
�cڵ�bKʭ���TAp�מ����d3Y�5E���*������u�X2$+6��r�)�jMV�d�#�Iuz\�����m����zU�ҟ�LZ�rY��[29�]�w=+�vU�͆L����i��j��d%��k�4��
�Q�Q�F6�$QD�9p��q�yFy�<�l/5�1ҽ�xU��l��h"%u^��I���D�_����L>oBC:�9�t�JlK�$���2��i)��-2�V[��CJ���\�(�6'��7�����d`́/I-������Vke00�iK����I�]�	)3}�0�I�]���r(�P!XK�嬀4DQ����w�L�@���}G)!E� 
F�Z��֔M�S��'�����/��m�.b���o�v�mON~�6����JGj���'ƤQ�a!Q�a�x�|:;�YY�����ÅT���N?��W�~��>���w1�q���ۿ���7�x��mۇO�L���������x.S �f'k��҈3�$.M�P���4�>3)%��v[V�A♌T;Mա (㻆P eQ�6�)��]<P������0���p�j����:�Ͱ����̌��h����������ǟݑu��=�\�	�@��R��x��)R�"�[Z�Ni�"m���q"��������������&GI�/��^/^�������y�#����(�ք�����6�b=E��C��H.���"��_�eW�
��1pTW���Y�6�j|~t-]�B*���& Om2�ħ����(��*���Z$��E]؍��j�e����Z�O?��#	,X��u,n������u�]���P����2�n	)�i�fhP4����^o������=n�v!>2�K��_�ڶ�HkN��K�+�<}	vKd��D�\��D��*�uK?��K�T�%����f[{J.�%{plY�D&9�BOK
�鋢q�t X��Z��&�]|T���$C*�m�6��f�!6�����Y�$�]�0l����^�o8}�ms�u�7�2o���ږbc��;�����ŀ��RU+���e�|�6myP��U�-�8>�%πbPJd2�'�5SMt�/������#��q¢='N�n���OV=������U�Ⱦ�K��HJnI>X��ЭI���7 ��TV��%�������o ����tZ����&�U�|�O��4�Ο�yi4���j�>�>�gH�����Q[ӂ����ͧ#�q��;_YM���u�_X�n�;��SĸwDJ-r��e��AjxU�j�m7#�4����O������3K
5�|rg	-�����K1i�4���+�������k��LZ�S��~�T�U8ϵ�5u�$�>��ס��9Uź�&L��IӦ#K����G��UH���!�K�W����eT�L@�_�x��ʡzn^?���$�[���Bv���U8���0�)J'+d��KB:���6�PW�ȃ�� =��X����z?Z��iS�*JPx��(�QP���ȓ�p�`��"�a65���Ԝ9;����k߸�7��(����e#�ѕ����?�)�lP*�;o�nG��H�v�٧\~�3Vn��������_����{��W�ߠ��ǧPr��$�LV����-5��ڐ6�ݵ��Ⱦp<�?���ܓ9�K������M-�j�c�C�W[���A�w9��mi(R˓J�dX�im����Wv��R�`w//>���y�&t��V�Lq_�d�3�������d�=�[ϲQlŚсjф���.�3�O�6�����Hs�򆄆��+�B}u��H�2����"0�7ଭC����w �=�V�����G��*��~�>r�$�>8C�^���L�lCSu��C���k�*,\�5��h�������,>Uնl����k����J�U�W/��	�ⲋ��b��8N�s%DO����a�%�{�r�����4���W_{g^x5����M��e㶵0�������<�,��}�g,�t�8��X��cg��j��R:$xP0��4pȱg��֣(���,H��Q@�$�].��D-�$���ԡ���A�����;�Ȟ�؆I���)[���
�sTK�j��Z�������b-k�7�:�ڤ��m�y+����sf]q���? i���    IDAT�n�VUɯA/�nꦠ�u+-��O]p�1��:d�-��-}���n����g~8y��稆8E��]�W�F�`G	�Ph*�L�(9b;}Z�c��o����̚YV.�T���g&<r���:6�b�g)����;v�wȡB]�)�;��:�h�:��q�Mwa���� -�WtB����sN��[`�������#�Q�$d-	f���Vd(�ҴqI�[��d
�j4t�C���"w�<��s��*���3q���">������[o������^|m��D�q
N�ӊ
��^?��	�����>�, "��^�	>�۟���s��Cc�����4�a��%8��}q�YǢ>twg��S/����Љ��B�hgPK%'�pASKX��3�x�{���@.� �����,M��fa
:�:�hհ �>����\���G ڌ�Xu�h��=0��.�����kB�į�n�p���`#�cY���
������*��\06��
&�����B�J�ǞR%큮XɞW����yG�=iV(����ݠ��'�5�C�C��<�����̺t��WO;�;���5[����A��m|��E�w��t��uX��3o�(ts�Ĕ���@:��-�^>q*�2���7cCk3�fe=�옾��X9�*O�̟xeW�ה�nt2��$��9�����P0�?<�1�yh>-��Ó��&�Ǫ�����^���	/��p��s�Ra�j!D��khD�0XjP-K�_�
�Ld4<~�$�,�	mq�R+>�'^��]�w��*��w.i��|�&�:���Wx����1mO$.����O�P5g[2R�#Y
VB��=�;�<��/�q̬ட1X�ׅ����R�_{���1�1�����O��_��I8kZQ�(@��C%[�d�̺uY�zE���#x��cj�J*�r�KC�
0:$����p4�:����� |ѭ�gG����i��M�i�D&�P�j�8
j�ۅ@]|�:h��	q�m-]��?�4�Q��Q��<�o��yغQ�I8��j�M���Z�0��ώ��ȱ�k��ژ ���+���5��y��n{@��j��ѝ(��wb.���ӄ�*tV���}v����߬������G}�o(au���r�;,���Q��E'�5�d� ���[Z �|P�<.�Ml(oy�x��'�D����pYm\�P*B�>ic˾J	��?V�_'�4�8dkT�L/:�^����Y�S��Ǟ+P!R��@�+@O!۷���ch��![�w=���~��qpD��m��+�k�������&SUGP?�95�	������ޛ���~�M��$H��]
E��9tSvP2̾x��J �2�B�H�QZ�sZ/Wk%�V;H�`)P�V��3���_]�ܙ{�n��1L���H���]�!$cыʭ��z7���6���x���%m�Q��3��-�J�\
̒!�4h��i��D_,��!/v�}s�1��{�#���Q�����p�]�k$��&�u��L�����kQ��!�&Lɂ�*�`M=T���F�W�2�f�U�~6�-I�'7��ڞQ!���'�(�\+�ZIW�C�Χ�1/�٤�6�f�^��9R�/��S�:x�ɫ6wo~�3��9��E#W����C�u#Hv�$Q�Q��{�3���.��N;�������W�o���3]��S�@c�&xa�Y�,j.�B6�<�ps3;�S��Rim<8�ڭmm0=.ފp&-[��'��5^�[�m�����Xf�-Œ
���k`�>���Н�p���j�{���~�v���E���䃢fQ�61�j!����񗳙z������݂���a�kᮮy���J�V��ף::�NeB$��gﾁs�=7͝�`��q"���
�X���4�� N9��i	�X ݎ�����#N����A.�G)��9�f����T��]��'7�{��iәs.�?>Y�~
��`*�ќ5���|F�-y�z�E�k�7�_���\����H(9h�
����#Y��X�T�y$xJ�.-�E�� ���8�'���K�X��^��#O<����:T��ۚ�α�eX(7��%�a=� ;n��/Z�|���#$ä��(���W�&��oo ��%F�F�ֶ5߶n怯Q_��e@a�c�9�Y��o����n�s���P^x��,�J�L���;��V�b��t�oN��^��>t���-�lx�}�8�����+����[݈|9ٞ ��d�Wr�b�47��qC!3�z*��p����0\
���<��e�����D����|�WT�V��qP�?�FîL�R8���{?ֱ�.E�0 U��+��1��&h�rC(���za���s��uw�f�TX�Zx���(�����˘�n�"&�
2�.b`��䔣p��C�����?���a��n��q�D�w�Y�}�<#���ώ;q�G��@5���،�q(���yIi3�?�m2��<X��s.����9&��S��K�3��`�wcð��0��,|�U����֗�s�}p�NA�63�_1 �
\��"�a�ₕ|f�u+���3N�/�"��lY^Ay�y���+X�C}�v�m�@�@|�8ѽ��ͼYc&JD���Zթ�d�ز�M�{����8�����P�V�ᚬ�����o�l�����!�x�Ӯ�+����p�g]}��c�]�r����/KF�僭��h�䒈�!Pjp��e̻��Ӟک�a'\�����ДG����{�r�Yryxo��eQ�+(��6X��U6*.&R��(�*�tvB�E�D�'��& e4#�~��+"G�"bSꉼ:Nv}��?�_}g���xa?"m�1�ס��%��O�5⅙�E�g1�{�D�"~�E���P3v2�It��Hd�>V.[����+DǴ�W�ncՂ���k/�1텑�?<���c��9P�Y8�U���8��Cp˼�F�xG�~%V�!Tw��d����F�9���e��Γh?ރm�x��kx���_������aO��U4eTy�U�~G�p'�~�H�<�W����P5ywK�e{�"��VD<��	��8�[��8?�o4EpӼ)�Ǘ�����O>�k���r��n�\��������&�-�������F(ڈ�(��-��y�~�$�
���}�d+���Z�-W(\��򌞡|�-�ް��ų�����,[T���L� 
oy��'�Egz���/8s�K����#�򾦱�E���,�|5�l\X:��kN��� G�?�cO�m��ο;����U7K����e�����Ɩ=OH�E�RH���'���;�$�|�ā���)���uIe�_}U�O֟_2��V�D�c"��(n����/p�n�x��y�~�m��}��Sv�#TW��7�A8�FX,�ӷ��ۮ�'u(�p������D�m���N7�x�|�Bf���Ԅv�nȌ�A����nƴ��Z8���!�P�ȪjkkQ���u�0S}x���# y���`�p���E!O j%4P,�n�'Fr�p��69��xm�o�ُ�y7���AM�X�b��k�,����>p3<�6��;��=������Go^�.���IQ/Q�Bq�$#���/p���㜓~Ѵ�d*��O>�уI�m���D�`5ɇ�d���P[S�\!b^�-��(�U���L"��^ɮ��f���蘅Q�7[��P�7f�T�ok{��R��F�h`��le�/
U($�����
g@Q�t�ל�Շ�1u�����t�r������W��y_Sg��!�j�ix����-է�s������򛟏��{��8���rPv�|��<�غ �dX[�܎"�JJ̘4
9�ط���\&:m�Y�o��{��t��Z�Ґ��4�߮[�f)� l�;�LR�����{�CcU��q\t�-x���:�f���e0��~��n��K%�Á3/�O��>\U�TGijD^'nid|�x��1cҌ���*�W.�k�SǷ`ђ�8q�lԴN�ᰝ�I����)I��,^x�^�T"s�8����?1҆T�X�n*�(r�>M%Â����з�߸�K�������Yx���'�d��A�������nhm�C�0�pY7N�}9\�0�5P��Q�G�ֆ��1[�#�z�~���=�t �:���\�����
U�(ȁ���8b�:d����^�.�s9�;&�����<^���ͤ�ƮDmہr�v�o��kz��>����_�$�>�)�͕Ji�y�h�e�k+�ɜ�����1ex�{ T5��s�:��c��i���/�u����s���v�O�fr!�*5��w�U?�wɖ�����?�x�����޼sG(*	� �n�luh6�q���v&�Q�M*�B��F�dkkk��i�H4�2�pd*s!i�A��t�<nIi=���Ǩ�R����%�j��s�c�0��x��kq�����KȨ&n��>|���(���05L�:s/� �!/̒��rN>��� G#�up��(r��DP�`��0�����y(K��e�����n�� �Rp�7��/�Nf�t�y���(*Y�v�8���핏˅��݃���Ꭲ`P̂]��d�$��6C.���jт�胞\�'~Əm�y%.��<�㦜!v�w������\}�w��7?D�ipU7 S�9o�T�d4N{m��&S(���^�朆SߓU�R���V���,��\b;��Dn�:���H�zԴ�E���냪;;vM�ame�^cl����U�1�|��eS �ي`����_k��u\��<��P�d�{�V�4�ϝ�Q���i��z|�ʵ���̷V�/W�Mm���
� �]L TL���ݦͺ��]��u��7��e��ϼ�껺���`T�<a���Q��Ns,$	Ӣ-�0������L�v�-ͭ�������RE�a�AJY�P�*����}��-�<������%bh�����ZtT{��#��/��S��L/Y��	��¥ ژ����[��W��1k�F�i4�i��uC��e����ƺ�a��ׅh[�2%ՙX��=���o���ff�(�8�.j���/!J+�\�| Ogϻ��#�H�(Ù�R�����#_�ɀ�-��4�X��˘>���~D�An��!��XI�J�5��3�m�>��_}m�C�du+�P�����5�ނ~O�
EBq�M.�r��"%J_0/������-H�ndQ(d�L�!����gk����`���m@�R���d��R�8����ٶgk���g�v��msKۥ�6K���9J��<�
i��R�.���s�Q����]۬�����~���ey_sk�� Qˠʙ�?���cN�꨽m���������|�e7ޓt���J>����外'�,�T"���j]Ȫ�zܼR��a��h���r٭;e6�a�r;uNⵔ�⩯�y�[v0��*U8�K��lj�v��K1mm~.3i#��D�l�U��9<�ȳx���1u��1�Ӄ��0j;���FY�B;��Ś%K9����Ӧ�6�-;�v�gx��w`�	5�9	�4�$��o������4��AdKN��v,X5�A^wp�B���>�:��-.KG�* ս��[�Z>��;{��L�<U!?T�@6�#�����_����;S
���Dm9��1Yg�C�AÀD�1��$.=���YK�,d�4��B��:8E7�֭�h�v��PR1�x��G�`�=�����~t6�*��y�F�h{�VF�'��@e[�}=�M��v��3��)g?�X���zz�?h[�+3�g}�-T���O�v(�)�%�w֞y�i?��?� �ӟ��+�x�mܓ����٧T�AK(�d� ���Q9��#"��#62��_k{g�$)����(Ƕ�ɠ�1yv��Gr�+�~����J�@�S	~ʃ<���:�#����a��q衇b��1�5 A�ey�Y�{/��-���+��ȗt�\�t>O4��q<T�g�'�ՋC �M�5�H�\����p�
\u�I8���()&d�Ê�P����l1"����M����������C��#�ɱ{m���k���|��i�c��jq�k�ᑻ������{>��C��ֶ�U��,Ĳ*V��`܎;#X׈X��d!Ͼ5�Ц���F��,�U�?Y��Ew��lda��`Zg3N<�htt��/���K�e}.|o���G&��w,�`����:����Ūf�J~����gW]��Y9��Q�\^?S�O�ԍ�ٷb���������l��3��r�B�P喇 E�3J��x��O����m���<׽��Y������[Z˅B���@Vb�ɑ�u�K~q�QOMv8����|�q�����\���MIɹ�O��%"�u-͜�R����H&��H3ᬵ��ǃX2�!�$�6�jg�T�Z��������j�d(�D/J��@^QIF��e0�~$c�$>ً:��Z�N��f��4���3e7l���0ϳ��PR�x�4~ҹ"��ԓ6f�2Y��5c��rK0Jr���.D%A���f�H�R��ҕp��!�ij"5�M��^�`9����u,��L�94�ա����N��X&|d˘���k���Y*�+8���W��K/����a]�P5:�n����R�)E�o8�eR���HCX;���(�C�9bfG�\���y�;�`P���>'�v:r�4�:�8�ڑ(�HE�b���57��<�翣v�T� 2Dd�N[R��@��Ӧ�2���\��كn
P����m��3gEoV�P<�������z���X��Z����9OcK.h�z(#h�|�P���S����5���;5�����S��⫋�w�#`
S%�B6�D��'Z�yX�Lx�>$bC�f(F�@Cc|~?'�N�Xa/p����l�����t��o�3� �V�*b!
4&t�q��DcH�����p���#�sx������Y��`D�����ŋ��������;a��U�\�U6�p������}�_���ހ��N(%����nt��]t-��%�T�m��L��b=��^�v�-�h�k��|�tNGu�$��?ToIUg��,/i9�>��>�e�A1كݷ�������� 7��5�\_���;}�?��&
�����S!���*��)�I��b!GQE�"*x>$�z$H��7x�����:����>�g^|	%3��~y�;�6�Y2��d����e�
8��s FZ઩G����$���-JńѦ��(���ͭ��b�|�Ҭs�3m�ibD��d=�P�5%g����7�lo;@���wf�uu�򌷩��y���)�J
�<�ᵯ�p��W�9f�������1�'_�fE_�'�P]�ԩ�/d;|Y&2�82�$��M�-pJ�����s)�TU��D�1L5L���mgX�űcT��vܲ[�o��4 �q
o5H�A��N����O��K��3�����ȑc["��Ӷǭ7�EU��"�8��,[Տ��y�-\]���T�i����!2�xC4��Z'Q�e	M�&B��cSC�{&U�p��������0~b'>��m��i*�ɏ0}�dD�>|��Ex��x����vڞ��2RE��F�v���U���n9�r���5t-�?�g̜6{�#ƶ�W	 �����f�>��+�a���p�2�'����v �V�v��u}�fGQ��#�L��{]�*�
~y�8���X-M�w�q���1�d/.�s:f�Sd����?��t:��ӧb�S1R �;�lU�H�C\(�l����ƀ�}d4����)�7OL�_\��(��&Ќ�ŀ�L�>��-W�2��j۵<�>��]���vն��J�l�u!��[��5�{�i����}�o���>�ܟ��rY�y]��4_}3L��(������`�T<�׍��FJ��Q��C5��!�N��<B� �յe�4�m���mP!����)�&��\����"[��Z|    IDAT`J�����TH�[���7^�=\ ]0q깿��>�~Q�[����Z/ovȶ���eN�s����8��gA�6 ��୯BM[+RJ����<>�Z��-7i�nkeH�[ĒO�������೥)̚}6��;L�믹�U&�ӍD�6L�~�(��u���7�j�����0�����2�z�4%{5.	��:֮X�S��4����p�?�.;L@s[y�^���偾��7?��>���d�7���^QD.6���0�iӢ�1e;$W������#Y���e\}ۃ�0e:>���x��c�Z$Gp�!'b�Kp��sq���!e q.Ҏ ��n7��,��դD<\l�
:H��gRQ�64�'��ƨ�ʦ���k��̮+&N\���P�h�-�x�����fV(�ė�LJ��={�ܴ͗ǘ�u��o���5Ͻ}�]�+SrM[�L�sy8s1J^�	�b&{�yԏ���c�����[�yr�?���%k��ʔW��?��jU(�&�#��f����E�����0��슯��<�s��Gk8ԉ��e8D^;�cѡ�]�*�e���m4T��$�%�Q&�Q��1��K��x<p�/�:}��E8v֙���������} �u�~��X�r���
�7� ��κ�~���f8�2��u�,��~��xO/�Fc�n3�T�(�Yw-���o׆��v�e�@,>��]����IQ�{��B�t'�U{z
�'�)}AQ#��Ks%�R2y��4���ݳȆ��B7��,��'�(&S���q��8��?�76���k�����
������G�C�E���Ibp��W��%�ɟ���+}�ӏ�	���\%�v�%X�*ƪ�=�е�CVi��� �yN>�T�"�9d6���p��ݥ�!���Iy٢���e@���r�o�uS�÷��z�}���6��~��6�Nb喇0��~@qٔ[x��.�ƀ�̻���Q楤�v�̇���PQ*�����".�?�8s�����]?;����;�>�?�o�����t1�Ce��.($ �'ظ�*�@&�T�:S����3����0 D����;]^��
�1KTz�{8x۰���g�]���נ2���C���E
���_� s����D��\r�x�w9@{�)�x���8 ��'���0��_r����%�r�p�Uw�wO�����A�hK3t�N�s�%�[�1�b�Z�w�B�šƻ���w�1�[�~�/�A
�t<���h�!�5p��c��e�{�E�����	�|ѭ�pq�m1���E/3W)��B���"�p��llKz�A< {JAD�g5��}����6y,��g�p�Q�n�4�"K�_��E�TZ�NC"�Gb$�X� |7�� �a�l/��}��6����ƑG��H��Co.��|�?� ��*��N8CkW��KOÜ��CB�9��J�0X�A[+Π��,�k噉�����m�ւʦ�[Z#o	���٘8�mC�rmm�m4C!�1���K��� ��+n�cLն�P�}�S�ѓ��#�CC�x��)��' A�X*����=ϟz�A����} @鿂[��?�;t ��9����c�� ���_I�Ja_�)����o���3�q����E�}D��"8���9�I���R)��;��E;��F�
/���E��r8:1#��x�n���.�-�7�y$.8�`n�f�}=Vw�#Ʃ'�3O;�IfO��n��A��j�><�䣨�8q�5����^Am�8&�5������#���F!=�	�����0��|{�<�\{>����?1��9~���o�K�������5+p�uW���5~�l��r>Z��DL%�h?��Rh��)L��[Ģ�D�8!��,r��q!�:�V�D�{�F�8���c�]g R���I�!�e�Q�;�O��&B��X�3�tFaHMu.����0f�
V~����q�(��:}6��d;�C��nNJl�����@v��[�;权#�:%����,d�AT5wb-��|l���T��N�\����Aa��JKA?��౥k���lP��m4���PP<f>)���z��������v-���<��ʸn���|�\�AZ�
p�)�gQ������jϛGt�S3v�5������ʯ�?�<���&|���C{S��1����!���.:a��I&E�%��/�PR	�
m{ �?����ɲR�7Z,a"IT��5���F��(�����/���ɯ
��R�oX�i3�Y\�����=��3Q,Z�uʙX���$ᥧC{{29'�>{=+Y<�胨����+o��O���1SY�S�܂�\��2
��l��@/<���^	�d?.��T\x�ap9L���_q��`�ݝ��
��?��c�8��񁈄�8��cpŅg�!9�ew3<���4Ҹ�8���]8�Nt��"����!(�Adc}�d�4}:~�߾�c�44F#��b��)���;�e_��g^�WkQr��38�,��#P��qqkB�݀lBO�c��:��e��ko��C�;Mc&a괝���M&��������D���䁟w>
r���`�L��k�
�x(v>�Q �F����v���?`�n�-Pn��?�m�N��6 n<B��8Y�+V���P�k����W�߲}��w�ʼ'�~�{#�+�R�9�0U�D�Drϖdb�h��*d59�.��Ô�3fL�|�ɻ���8
�)�}����W5�X�z��ޑ=���!���C"V�7��B�l'�1r�NxD7��	#�C:1]#屉PU~��#��M7�Lt���eP1L"UW��I�^r�w:�
�W��5ry0[iyhg�b9�`q }�#�Dv`��s��"f�>�У��mwa�λ⥧�mO�)`�}̈́�F�p��G��ٳX�{���7�_CS��Y��r�����"E�ljH@�d�r��Ļq���+���ѧ_��g�F���/���ӧ3E��g?��>��Y����]�@�Ѳ~|0n�O�:|<�%N�Iw�V7�;RrplJ��ƪE�F�0�����mG�8c
�t��P4!�/�0v���?���/���ǞEwOU�Z�A�N-��j�~��ߏB���T���v	~w�u�u�8n�|�Y�t����Q[��k�ޞuhl��u���~�۞���_���g�n�t���&%�ۼ#{XA":�NH��-ʖ7=�Uu2<6u�ln*$����،_�o�L�)�(^��P�B�g�#w�p��o�6˲W>���>���%�p��8(�ep���0H� CM��(���Q�r)�$���|K�N�f[]Mo��κE���2��,�,�X,���%�Q��L��tFٮ$ޘ��C�[�nDZ�Q%䑑)�a�ND��\��n��D��&��
�T�����E����$a'�:y��2i��i�2Y���� �� �^9$9҆�s��f��OӮ`�c��)�����عލ?�w-<$dӳ��C���w���w���gˆq�ɧ@�Tap���:�ل��9��O�.�����"D���v8|A��*�+EDM��J��j1֍]gt��n�,�x���0k�i��>O<���1��p�)��`�ʅ�}�Ѹ������r~�e���JB��A�5k"����⡈�O����n��"�S3,��O�ߩ��t��Ě�><��S�|��������22��(�\�y�o���q#G�+���a�DCP��Gׇob֑?���_ �+"��a$���o��O?��Rľ�}?9x�"^������){����-J�^�۷��N[I���,�h����?�ܦZ�-�o6%�8�z��9�e�B!@��\ґX7���i��t�?uiBՑ�<{�%\�X�Pk�L�9Ȕy�Ӱ6�ZВ�O<r�+#[�g})gZ��`N�kNo��U�2jx$�f���2gMA��b���#��Yq�](��̒�n�(��.�`�(h��L����UG!P^�A�_j��L2�|:�"�H�
Ѫ($�qMg'/��\�wne�D�\x��?�a+9�r_}�9��sfegS�wAC�##�.�w+���� ���c�]���W�iк�)�q��H
>���yZ�W�
�MmB�JΒ
�0��Z:�d�jx�,����n�$����ӍI�&���t� N�p.�Z��ŧ��;�ǡ���Ŀ3/��~��13Q��6?�aA'��ɡY�2�/04�C��n3p���A*�ҙ|��#X����n>>�l1�s����!_("9Cb8ΛB]/����P�-=I7D�n��N7.j=K��H)eh5�~�|���A&�O�V2sgF�$�3�H�ח�8圹����X7���B:��)�~���L�nw,�m�@��7���1z8:�F�ڊeK�M��Ǯ\{���Əg+�)�v�c-�	��{\$CI"�5��_߲ME���?�|�[�(���p�B�#�hcB�MSh��9�����\	S�8 ��;D�	���tѨ:�y[�Z]@Q�@ɓ�����!{ P�7��7���$;�;�,�ײ�2��,V65�F�R�@�:�P4�>tC˔67J6%���W�.��X��t����R�h�A���Ȥưs{ypK�Cٽ�S��Qm��X/�^z.N8bo�(��m�,w��I<���;a<�{�����-v���7�=w?�?>�:v�)ECv$���dq\�'������
\����D�k%v�4�Z�qٜc�#�1b�isZn���x�orPۡ?��]w>c,��^��R�ؤ�PH�l���*���LN[���`���x���0���-�C�<��/�S!Tݎpu=\^�yPi ��#Mv�Ԯr0��pc#�Uad�<�X�.7ky\.	��"ַ%%��H�]+8&��FW_{�a�8�l8ӽ���p���͏>GU�8���A��SD&�D$ �,�_)��R��NGў]����gkAbt�R9��q�W��*<���F{�l*5p4?��-O����&�;��8���d]`'AR�F��w�u��z�77ݼ{Kt��<ҕO�uɇ}�Ei�:B"5��4C(�S�&�Y���%)�LC<�=��)�@+�'*o]�M�L�t8e8]p�^rN�T!P�)k+l�0Nv�(����r�J"?���S����zz0��*�pm�\����������ܢ�����Q⋞����IC`'_��e�OTu��,�Q���w!ֳ�� ��}T��𫁑8�\��o?�+�\*����|~��>�t!|5���Q�k����TE��F�}>x"!A/D��٬������ z-�y�N�����-����ʞ4���W��+����	}]]��spʱ�������;�L�e_�K>�v�͆���y1+��<D��I�Vc��(�#�<���Ԣ���8=0�����(R��Ɵ��i�������a�5}��m�T*�#�ͨ�t|��TW�0l7�����|����a����|�{�|���t�a��5\݅�:`y��K���r@|!�B��]3��d�)��ᡸ	�h�� �^�o���h@���k-IPF����Q��r�W~n�ǭly�J+��G
y�PQ-�p�i�
i�R)��-���=�ݼC�o�����fY�8o�[��߯���Ѫ
���(f�l�L�$�1�pW@w`�+�U).%r�!�%�@�~�P���d��)�|!�P�B�)Ě�� 7��@�bo`����A�@�_z%E��V8j�~'PE��a���y��nŌ%���+��3���dȣ��,�m��/�7�dھ(�g��RI�ih��N��\�uCK�@-�Z�0�N4� q��D<>�7m�(�"\߀�d��T�r����>y>T7���A2��*�.D�׍l|����P���{����}���M��ā�X�Ս	M-�0��,ayw7^��tL������f�fl@a��m����d�ֲ.�F1ޏ�KBmu5�Z���#�TmQKSd�ʎ�ٌ�͉�����	��`�mr�'�;�K�˴PȤ���y�E74�&M���s(�w`����L&���PP�=������b0���l���׍Tl>
��ϊ���k��'�i�©D�g@��
���Q`�akcؖ eõ^�>R19���T(���p��(>AK(�_=9���n١u�:��P�y�߼�>}N�U�K�y0b\���|����iGYN��x����{�N:�9��)A�Cv�J��|tcR�Md$���Y� ��н�ɻM�L��H"�wh�D�C�y�K"�1ml���-��e+N����B�0���p2B�*E/+QI=�Y����4ӡe�]A	�ȀJ�Y+O�R�7��֍��I�F� o�|U���K�$�.Z���SIB�`g:�=Čs
hhj�*���&&"Dqd�Z�T��`)� o8���A˩�\�Yn/�N�E'\>/�Z�9t��a��ˮ%|��T���-�bC��G� �JB�42|vR8}���"��jxB^��( ��{���\���zQ�*��_S��N���@%H�>��4���lb�����Ls��n�����]͗+eR��Z[dp�a,7��Noȶ}�q;��ߨ$6�;�Px�C�����[*eㅁ�O?q�7��^3��������o�'߳,K���7��g�va�]T4�k�b˿%�مt�%��h�W�T�<أ�O��<�*�Z�Bh��ah�ϕ�d��ʇ�)��qp�q����5k�5�Fjh:�d�_8 712}^��$�FV�u"g#Q�'�/���B���e���!I<����*ڀ�����Dv�0t���0��	�(����*�.�=G`Ma�+�TA���E�������N�p����I�D���T.�����D�E��a"�uA��2؋:?�L%!{\�iE�s*�h*����
��oD�r g8`X2S�uS��Y`�/OөM����!g�|��~�Ai#����Ap�a�4�����a��CQx"u��"��冮�p�4�i�^� >��X`�TA7P�Ў@�d2���m�F�k>������m}vb���b
<sRLY"z\�KJ�<|^{��OG�E\j�
������u�l�p�1�H���٘�:�j��
e�{���g���*::I�I��d�me+�╉z��#����������
P�+�|c޻=�O
��Z| z:]����g(vb3�h��f{�1Z��2����T4A��{⊔��Bo�T��6Z��T�ʬ�NuZm����VM��(P��T��Ɣ�'PbKֶ�.ֳ�%4�$6-o�<n^i��+�u�d�̪�
�@�'dA�,�]��̧��g,DCA�)����T�T2��׍4��>$sE�L��GuCo��&(�
_4��T��ҕX�K-EKk�A?2�
C�����jd��Q���:��YR��d���A��bK���퇯���B���4c07�tdn����tNAɁ�5+�������K�k�/�42p�h0,�!�)E��,c�t�y��ԚZEJ"%� m�i�7q��� ��HDJsyl���_dq��,��}��E��?E�0K�t{ ��I%�������5S��u@�kհl��o���������������3��P��nLn\%
J��I����o��_O9�Pc�;�*
1e	P��~蕡,	��$-����+����b|�_���!���h����:]��	Sj���NAU���O9�+32=��Pn:����E(�\C�샚� O3�( ȩ�4���*1j{��"�'� �j��SC=�R1��^4VQ̨���1H�R*$�GNU�.�b]�yC���."۹E(��a@r�\#XE��8���C�U[Uu��zeT�xMZ�B��	�m�������e��;GR)"��6aD_��:�~����-&�����T�X|C���0R�p�i��}D#���(�4	��zP2hep�&�7�� �.XY(�*RÃ��v;!����PM��^�A$r�\R�    IDAT�,Aل�P�Z�b:��H�I�@"�C ڈ�����|8�������ܞs�fǬ�U�� 7�n�cf�{@�}C�S�.*�m��_e��*��
2��M3CZ�:���2�<��k�jن�"\��W�ӫ�Q<u�р�����2���B3[�˓��u+v{\I�fe
:=l6�= �Y�;
p6&�T��/��W^�[|�PXY�J\%��A84���்d�g��3��i�L�W�~ �` N7����,4�4�o4�C��PHŐ��B�4����� �Y��Nbp8EQP(�&�{��q�p�����Wt�@��ֵ��F�F�z��YK��q�$��<{��bkG�Ǵc����G!1�T�$G��PS�m$:&LFcs'���WT��2�i�;e�q�n4ڼхNv����AS�^�S�*��h��E|��_WQˣ�����u��+��Sی�S�F2o��
��V�M��5ѺXr	���B��*���6
M���6���.)��a8�)��4�#�����P���ڷ�����V-#�<+�u��e[i����ѷ.��6([��|l����Q��P�B!��� ��+�j���Օ�O؂��V�ۖ�f(7��ޥ��~w�B��,;�S�SH&���'G�)���T��_��ѿ��,�ze�X�{��r�b�E\)Imc�ͭ�*/vt�`��Q�i�J�r�F�F�bfr(����Bg�+�C�.
�����Yx=��)�r5�u{�W���%���X{�b�q7,h(�D=���*6
�$��E�(��O��iS����n��/0�|��j���p�>��c�a8Q�O���l�,�op��C���0���E!1١c��N��5��T�����ވ�>{�B~7�싖��s��I��?KG�sP��x�,��TU���I�j�4�(�&���(t��k�;�������3���m�nvC(B1���H��@ A)�4��h@�XP)JU��?	%�PJ
I�m����u�{f���,I���?3���n�;s���y��Ћ��+�{Аp�A�a��S�nGKS=�<�t��N@CS#r�6�on�	����8���j�[�Ptudse�0З�x���Z���$�x�{��j�lBϺe�Z�G��>�x�Խ���W yŪu��������#3N��Hc�ְ�;ϬE1`�=�B�a�-�xjQGe�J)��>�N
y��ȿHo�˸��+�T��IlEgS/E�4�Ph�0(kH�8��6����n��7N[۹%4xG��?z��냯t�u��!s9=��v#���*XS�>tAxU!V
9�1�i)Ĵ�GT`2�p@��D�b����^=�J��8�34�i1�����h(�
(��&a�\��:d�`$M����i3������l��Z�2�bX"+�%��������l|h�ވk6�/Z�L�3/�M-c`�1	�Ҁ"�a�������s���OFIK`ޫo�5���>�Rup�$��
Gß�@=4&L��}n�A�N�S����4�7�����m׉w���F~Gɕ������8������X�t�]h�1����Э�Tt�=`�)���n\�gv�7�y�<i֮\
ߵq嬯J�xMR�Ar8>��~s�l\6�*��8	q,�t����7����J���	��Q��tS��SȢ<Ћ�vnE�s�.yq�~<N9�����?���DH��Y�W]u�������A�2�@��0�7;P���Q�I}���B�j�V�F#n+�DV��g�C�g�����P�Q�����q�%�:(n���������{
(W���o>�1���l�!a������閴1M[�c`s�l}(yv%^��J��Q	:E3ʫ3�S"1�y��8:A��TY(�zT�HM*� t���E��A!��sS�#�X*�a�x�����������H��nW�$�L��\BeLhJ��ysqM��+Q�P'����4edz;;���$i�s?u���#8��Ē�>��/���u�)"|�q��&�:ó�pnłg0&c`L&��{NDmBGgG;�u�u3�e�o�`h�YY^{Œ-��٧��������K�pej'��֝ї+J�3M7%ݝ����b`�
�hkJc�ֱ���}ݸ���ń������Z�{� �|��~�
�yd.f�yO<�_��۰}��&"�֠���P2�z	1�m��
[k"��c���¹����O�ni��y�V\�9R�KX��������_��85�'�疠q���4�.�[�"$r44�I� F�k�
(#��w�B��R9�#k2��,�q�P�}�B��dn��3o~/]}ֽ^�TG��l�9�g�����݈5Q|�7|���P�lKe 	2�b��";wۡ(0�ӊR��0@ٺ���K}�P�r��Gf-��y���\�\�l�Y5)4N�\{�zL@�8�����P%Rl�6�at�����ՋȤc����c�Im�|��(�I�	ȓV�b�8V�Z�~�#�b)��,X���J����P�`/"�e�+@<pD,z�k�ò�p����E�ٰ��tv��7<�G �D�Z����/��E���ǟ�L���_<0=����6e)����<[ e�����݀C����cْŸ�Ο�����m�\ϕ�5�bL�E��޾��i���tt�x���h�u_5Mp�Zh�Zdˌu��ˀb�:N�܆�'ྻn��M�眆1-�[R��ؘ�,�X�-�2��p��EØ�8�_����,�]�Z���V��P�?Q�6��$��n���:��o�[�h���A���Ж�
�%P���o��5_�c�z���ry�+~��Տ��/*Ռ�ͳ��Ķ- �ϪK�C�E1[�
P*����.�DL�u����:�� U��G��v�ꐯB�(HZ�:�xB
ʘeF�&$y5uh���%(�i������������܀��&�a��u#��T��ϲ2�I� ����s���}/N9�b|梯`􎻠f���`�Q(2U
4�Xp:�����=Zq���Y3���]�c���t�b5��C���lE�D)�����>�[r��ܗ�+��uY�<%M��NAp]���r+_|�N�o_q).��\��8�cǋK�`��(w�6���-�FT@S;�c���7���>���u��QԒh��'���p|�[˒ r)ߏ���qOG[c��3�J���N�]�G<�R�����DpEs�� ^{�wp��~�����m�+���J�-xf���"2�1mX&�Mm�E6�;3�}#�ֶeC|+�g�8�zo���W�xH@�%8�p���
�;5�W_wٗ~�g��Eݢw2��_s�?f=�2w�S7�q�j�l�ؽA�<P1�<��R(Q7`�#;�2_=���,��7��y���\���(`���f&�f9%�t]�twK[S��k�0��^�@./<NZfu���0�:fZ3����6�2e�]<?���a�h!�?_t��%V��]�e�2����\p�e��{����Cg	h��+bc`$2(�t�ȭ)���������g����<>u����&M�e6�FE��U�[�D#A����4pٗ���f]��>|֖4���>h�:I�JaMIAV�8_��L|��sq��g��oF�����n]Q:��1*N�RӰ`]\p�L�zǭ���g`��NL�w:�T=zX9��=fYҦ�t�ÔG�?܃:��?��L�m'!��I�N�L��`�o����m,Z���0�����G�c��jGK�tQ���롄fO=�jɊ�3o[ �_��>3���1��rCEQ/T᪲P��0�	��Ǹ��b=(��ۘ��~����e�����_r��>���������)z��(nZ�Bob$:���_ ic�zp)KQ_7	+s飪c�!;�K���-��#bEA_&TiB�lS�&�5�oY��
h&�~�ȲY��z�eK�m�QMh?�iѪ���ւ"=�e�������c�Ic�*��yÏ�|`�)��V	{�=J�Z.o�>wU����q��n�mw܈���>~��Gж�~��I8f
��!�4�s�N,}���g`����c?����Oޅ+Yz!N� ]L%��a(�>b�ݞ��}�kW��܀]��.=�L�d���r$�� X��P�>� .�ܙ8���ǎ�(��.L�o�pd8�d�&���Y�ڄ��S&��A��Ͽ�������3�h]7Z�~?��z�<] Ŷ=$�����,��o<2��H�y<��$�ϑ��(��y#3IBeD�����"N;�\\���W����֡_OH�)��	(|�2+��șB�K�/�
����P0���+�"#��?q%f�����S&�_�+�{D�$2���;f��nx����,\�ּ�^�,��v�}�����T����U�&���qM�v�T��0�<���[�p0����
���Q�&٩ùƐ�TI�@���`;�;{�{��g�·,Դ4IS�4nNd���%X��i��,�J�t҄z쾃����c�<WϺ��u�Ѝ�g1�$S����Zoƭ���7��c���R\<s.���x���󃇠�l�B�-D�ۻEԛ^}�Q�8t�}��8x��p�i�_�e5{���, �s�����q��wc�K�1���p����&�&�Պ��ir-�vF%�4��x�~����k_��r0���g��aL�dA{:�S�ĚhY��q�w��o߄Oa&�=��4z-{����t5pr�z�Q��ڔ@��g�ݾ���nL���
�VD������zl+����x�Os�ً.�׿s#~��x�ǁ9j�X z6��!�P�2L[	3?Ë�ގ�%K|k�(�C	w���5�Q��;,r���ˑ�G���DQ�/r�b�	���^mM��{��ک�����p߇��Nb�nG�����5�-��oQF��2ܟG���� (␂�AwgHu�j���^�������d_���Q���mdu��:�YZ�>
�?�ʹ �z{�
(�J�aK�a�S�U�9RSc�ti(���#�{q�)��<��<��ӟ��m�`�riZ�K�%j�-�g���<���x~�J�6�G��e��i�Aٮ���>V/z�i���1���? ׹��奲�[	C��aP6({Ф+9о�>�Xr�qH�7��_���m{��v\�^U��m�'�x�I�S~��c��W�����:�t�4y��2I�%d��e����aɆ��HeZ0z����/�O�ctۮ(���nJI��5Uu�z1����^�k�a����;oBCc
媀/��G�YR���"�r�GQ����;~���q/�hGP3
$?H��H�$��6�wG�DS�SU�Z_�����T��,��Fs��5�]��p:7CMZD�{*6g�SJ���t�$���Z�5	�9�X���������qì�nmi��շ���:w�����äO�������rɑ�W/���֤��gea�MB��sa6�*v� D�d��ڬ���Q�&<O�n�5j�����SI�ER�H�2��
\���Xt}#�yX�#}qنA�5��q��qX�8��&4m"�9��������]s��I�B��
U�!;������;O����_�yK�lBMc3jG�@2���	�S@o���&>����1Q�ۄ]&N�ׯ��%�%�[�%H���J���/AGO;��/z/.Y�1m;!=j�A��W�:�b94�M��}���Ҽ���ٿĂ��.[q�	'b���a���j
R��cd&b�y��x��q䌏cѲuxn�J�2�Q?�MJ�ˑ0�y ƍ%ۍ���1	����7����w->w����x�r�kG@ss���Ƿ�w�|����>�����d֢��,�d�p���(WA�)��ʝ^����^2Q��1�)��U;IE}�X��(�&�~_�*e)�\�ZQ�'��̓J6В��B����6T�%��g�� ,�ѡ¿�R<��uҦ��g�O�C�m�]���[�{��!��������ޏ/\zj}�ngv��ق#)�ZYhČK�y�V̐݃-��E_���FR}=b��ZS�1���[=�����W�%
P�Qms쥹H&�<Ebs	�RNAvZ!�������T&��bR�k-Z�c�_(��=�$�=�|��sPS�L�,��(�Xtp�7b�S��#���o��s��cc�C����v+5(�DfnM� �شz9vn�Ǿ��a���?�(>�p��.A&S+��t��}�l���3���spȑ3��7���@��#�،�1��.(&,���F\.jb����S����i3��k]7L���G�G��L=)��`ل�����q�mw��?�'�v6Vo�����aC��q03M(�P���H�ct:��_D�͡Խ���̙�k�8�أ0~�81��lU4�z;{p�M���?����c��++�>P�c�!�/ن�[8'T�R.�P��T����+�"tV e�L��h�Ʀ�qͨ���2G��)�V}�%�͠k(�!ͼ�#��Xv�ۘ8~�;�,�wu����?����2M�`�V�w�B�������s��]�2ᄞ�ߖ-yR�JIAJ"zvY�](ːl��a%R�_#��J�-rUF2�x��{��(��������>#�V��CTT(�Qab$v,���4Ud��!��И��������3O<�=v���h���a:r�V��
���~�}�8��"�ٕw�ʛ�$�XFK�M���i��D@*�k����w�#��hۄ�`j%<��H�>��O����ƍ��òe+p��?�W_É'��u{�]p�b�&���!��|���_᳢ʙW,���ѻ~��[�2��c�=�8<��|\}�U8�c0u����҄l����ǟ�<�6���X��,k6��Y�H5��k�P��5I�S��	+)i|�)	�f��4�-Sw���^Ɯ?݇���#��O:QL���N,\����7�pp���"]׌�o����׈d��{��d(���=!�8R��+O�9.L {��N4�%9LR���Nx�\�q%�JX�9�6K�ql4�p��,[��\��ڸg��C��}�g-ݦ{�ܷ��m~�}a��+�}����rZ���'��������V;�ZvVex�ߕ����2��-i\^�t[��w62%+�y3�#��ؐ>b&V�Q2#4b����]���Ї��X#VĔ]Z1�9���Cq��=�T����Jףu�=�X�����������:�L#X��P�HwpN�^5�IJ�X����N�Ԋ	��1�FGϦ�x�אL��uK�����C��	�m�"^S��\��.ib$3��5��V�B�xB�~i]&�I��eS��x+���c5F��qL#2�	l�؎��:�:��`�Ey�6m:Zw�%WC��>�U��S�n�"���kH����p�6jk��Ƙ�Z�n�ORK4�)�);�b�sOc����N$�J�*�B�]0��#�zC^_�������cɻ�4��,%�Š%���@URaK�b�8�H����A7���^6! L�C��Z�a:��)Ҧ���XalI��������kž?\{ť������n���X(�-����=z�3���'�xfb����R��"7�<b~ICр�`3�Z��4>B��E�S��#��0��P�Vo�\:<gU����C�5.!u�EVMt�\ЬK��Ei��<�]���DSMB�e\C
�80vu��-��Є�j@��c���� ��ғ���^|E�b�/_�b*��s��=�-]���,�SI4՘]c!eR#$�ڥT��Ģ�FSs�%��\��V�E}���ĩ�VӀ~����$�-%��3խ�`y>4��yx��{֣)�����ˤ�HX��E�I,�0��Mjy<_G�	�����ڨm�AT�==.	��"�iՒ��f�l$o�b����C]"�:����Ic��ݐ���]���XӾ=,��M܀u�pؓ9�B,Y���|V�C�t�K#�ٜ0� h��ɹ�~�����~�H���uhM  �IDATQ W���k��,<*��a�&DD�v�=��hh���i/��{բ�>��_�<q��&o��*��K8��ݟY��'W�N�2ͻ��dn�D�[��ژP� ��`<E&L���bU���D@q��
�s���Z��盛Jt�� CP\]�H��XZ]#''J���3�1�T͢$�".�*6jR)�Z��A��ץeT�����R2�I���d:-�]�y�n�B�EC�8��Sw��Mҩ�+\��%�5l5��^Z�r)��MQ�Pgh�$0j�(477�q�"��Ne��}=:���/���=Ԏ�Dm#�x}�,�+���f7D��Ne/+�Y��3�F��PWGm"�QԵm�C:�R��$h��zrE�
���q;�HgD�������G ����!S_�\��G�����R�H�nM̀EmQqrOYR���׍�㢯 ��[ȸ�4ݒ�V��V�+D$AyDz(�ݥ)��
K9�]�0���W�.W�����f�-��y9�ц�����fAa�U����\v�MMI�ȹ��4�jj�i��������k�|�mg�8�_�9��
o�[���C�;!��z����޾�Boˮ4�
0�<�&o�W��Q�D��Z�F�i�0S��t��<S�{�=C�����Ku[*��?̂���	j��P@cX�Xv0�b�s�B�"�b:�IS`�z��P
�-��`+L�v��Sr}���R�k� �z+T�g��Jcl�D��P����(������L�F�L��tIJ���H��h��ac���'�M��~T�z�۰R�1�|�+a!J"`]vؾDGmm�蹒K�wB�`xԜ-cӆ5�U���LW]m��|���a2C������Ae���=�Vڔ4��ٳ�cQ��ԥq�M	S��9Щ�K`�}a�?��?j�@2݈\ɕ̚�H�d��Rt{�)mb5�� �C����EdA�իb���q4��F������78�̄��kP����P�F�����	)��D���4��O�^�t�'u�O~p�g�����-�O �r�Ӌw����'�[&~�3j[�z�)3GOo'��|L��s�Q�d���{*�>MI�Q�)���#��T�~#W%�a����]N���ه<�PІi�a�6�f(����CuX$#�1T�'假|�(�H���?�!����;�T���p첤���L�IH�uu�ߋI.�P9I���'�nH�@^�\����gK�Z)'.ţ�.�ٚ5��3ٺ��J(��Jq�K�/�)�/����B"���҄^��)�T("�͢X�#v 0M1+%r����5aO��T��zQQ(�K	c���l0�,�m�c� ��k`�@�d�U$�^�t$���	�^�X�J�yJ�QVEbl�����Ӻ��E�����Չ^GZ���O՜���D�b��'&�H(VV�aFd5���i3�$YR'�N���\����x����ƻ����m�-��=^�ϞY�����Q���6��o��ME�Q}j|�#�PZ��B"P=ĝQL��V��R�>*�B�RI���i���W�Q5��.�IBN�C�F��C��bF��/"��4�*@V9d���T�6~��z��m)�@�⺐oc�.%�r�!��R~^��T��M��Q���^�<.�0����ku���&���G�G�\�K�)8D�K魐��EO�P��A���ӗ�
���r$]u�T��e���,�
�w�a���2l�ّ�*��AT-�(�!w�G����+.`XE.}�T���6�Ð\���j��{G�`P�-�"y��
�Uj�e�k��V�Y&�K�����K��T���;B�`Cs�\R\'�����]�@׼~֕�ݓ�i1�1�W�Z���L�GW^3s�q�
�_
/v�������?~p��S��v=��AK�AG���Yw��=t�Vz�T���WWT~"��|H�se��&���S�j���+ �|h�N§��.�=Jg5Lʇ��\2����YT;���Nd.Z�NK�
%@X�
���E�@vh�I��=Q�X���~�����;�r9e�q����A*��a�����tٖ��B܄0�@ғL��P���<���������!�@�@II��
�ʰq��(Rf�����ȽDmc%~�
"��T��P�F�UvD͗pDEmP�$m�0ҭR��"1��(]*����6�a�L4WF�)� �]�	�Vh��Eih���l!Ɇx\[,<�j碱6Y0J}�d���^��3�=m��cl+м�JtQ+� ~�7n?��%��h�8�Ȭ�1��H2#�bD#�D&_�2T?���r��#2���������C+���0^�����b	ؼ+\�Qj1�`R�|�2\�(�	��P�t��-q3�a��v��ڕ�i\�!�E,/�ݡV}��<.��S�|pտ�;�4 �>�aV�܊0P�8��Qx�甓�ą�S�����
��F�����J���`�u�]W�ܗ�)��H ��
F�����'�eE��S�i8F�TM�ʫ6�(Ū,U�<hy���,�R�h�yj�,Gp���z1VϽhÉD�e^�@]-ǡ�ڪ���qt�%~"�VC����b�*������b_�R����7�?�O�8bͶ����o^���A�������;�ɩd�-��5x���NY��L'ҏ��ѢV+���,3���J�@*D�ʎ^m/D�5l���\�Q��c��5�"GSYޠO]ya��ȃw�ȵP�@5�$�{�R�62>eWe�6ҍQ����<�\��d&uf"Cɣ.?c�9%�H�L�R�.4meYHp/�����'Z�T����"l��$��!�g��Pe����%�|	��g���(�ɦ�"I(1�@��L��Lb��跄��K�6K���#R	!XWeY(�-�4*�2Tx���=+1�D�my=�v�����u1ʲQi�� R������e�M�b����j��!��ru86��E�-J�&e���&gF1ax��r�/������s�/>}��+�o���m�]�o��e���@>�ݫ�?��Kc���Ƥi�+a�=�{>clZZ��d�Ax�p�@��QL�=�иP�*��0��=�Y�$�R���{�bUs��ZĄ�u]3�X��3 z8�zW��L�0u� G���E-ދ�)��X<Q ��M���e�����Y~'���0��-k�V�4�*S�d�r|Oc*�#�xɁz��Z,�.�%P���yI(y_e����ƌ1	�W�@)�q�	�WȄR�"�]W�:!F�9j+��/Z-&|�a T�dX-&��Bz(��%e��fSAƁxMXS}�yG1eO)�UJ�ZH�7��X	lQ�]m6aVXoT�"��b��t �q���K�����[�~0`�U/��i�+���N�O�}'˞��)I��fm���w`ug����s�	�\r�ǖ��ؖ����y�C/��A��/'����K���lϫuK��9I��)����z��i����� A�#�)��)�o�{����g����X��M���R���u������.���+���L�`�80|�H%�0 N��C�ahϫ�1����+�_���g�'��Z PhB�w����+�X�Dt�8~�j#+���@�^��	�]�/`	rh�h:����S4��H/ׯ�q�vO҄$z5��y=�W�д���>�G�Iԏ�_\��=n���~�������t]��d�Y�cc@Mg��i��k.�!���끯9�Q<<¦6��q�5�W��i~�It��d��e�����e�X8^/�b���z1_c��)��b�0D��dFQ���]��y�Lh��f��v�2�AM�Ø�� P�� K��oX��<������5>#Aj�	� ��L���s�O^�o�|������'�}F<���.�
I��h����k��7]��6��u[c+��?(#]#ײ������rD���N��S,��=KjD�@��!�Q���e*:�yM�5��]~]� ����3�R,��*��e���*�s���O�4Һ�4�_�
,9�:bPɡTP��BS��Ӂ���k�*����1��>���e�~ 5^m�Վ@P���f�4���B�kQ��V���Z��4�X!��gtM+�J��?���ۺ�eM+�=岦�y��|��?(���oV86�-T�\��%8��U��s��h���%QIw]3\�aL�w뺫y:��9��{EW+�nx���nۚ�{���ٶ	z�o�%�����m��s�0D��#Թ�<�����̀(Å�m�w��=݊���p��M��cZ��<M���\���4O����}׷|O���C�Q�;��%aN�E����N��p���?iZ��� pL4����]��<�e\�ui�j1�(%�xъ��I�	N���t:�Ӄ ��̾�����;o��n�� �; J�O�}���;0D�!�H�z�|O���w���\�O�P���~��#�4��?�ao���#�n��v@y�Gx������l������V����=�'~z��^��    IEND�B`�PK   :�-X�L�,� o� /   images/50816f02-2fca-41dc-8ce8-89c3cd37e619.pngl�s�%0�-zڶ�i۶��i{ڧm����m��}ڶ��}�֭���I�Vv*�T���ΎTV�F�Ǉ  H�2�  $  &�$�w��?�����f��  �J��{\t[�ٮ��<	�/�2�C��"G������C�@�Jb�*�ȱM'Mӽ�_&1�)�;dc��.0S�l�Q%ÆDE%�b�$g��?��=���W�����|潕x�)}���|})�;�ݺܺ���U�c�^����W��Xg��P�_h��1��8��q���/���F������Ai��������?VXdZ�����������u6���7���"��d��p�@�l-� ������9�r%,oM�?.L�)3�ͤh�L����!�H��iۜB�%|��D1�LH&I��e͑�qe��:�%�H{�%�W�Wz��ꙺ���**C�ɫ�~�T=wI-k��/7���Ì���e)?#)<_n+v�\n�j;�x������&����Z��~��mઑ)d��U��۝�И�ѳ�<-�x���]�hS]�-��J��zx>������T�H���K?�v��k=�{Up��p����S�����M�Ae�I5�ID���5
���4u�,h�G�uR)�?HQ˔O��<�n���4H.��l�����IbfZ �(4�R�*C]
��&2��*u��
x"3��M�o��}릊"_Xl����a�2����A������/]�/��M*Q����?���(I�WCD��� ���Ec�o��kr>�i�U��4��~Y��yެ�U�FCRE�S婱kI�_z:��k�mA]C=�\!�8o��mU��[�B�r9�Y�BQ:���	ċCT0�YJ�8�]�%f��f'��T+�j.B��A��h�q��-�ApL��Q�%c��d۬��@�7X�̈��D��e]\tp5���VխwV��+TdO���m��T�����0�N�=�4���4؄���bS�}R�ca����^��_[�:�V�_�:,�l������^��e��s��ڊ�#\Z�����{�Z�{��<�[����Ϯ�>�H��1�޸�Pf�d���S�R�-�ȱ�իhT'��� ���e�B�C���L�"��Ѧ
���2	��� �$	�XU��@guIץ$E�✒��*r�?��ֻ^�v�n�ȱ@B<�1�J=�� ���gn��)�Hq+��[RE"����q;A���w����O�YeT��n�5i�#�d�����{]���!>�� �v-�i�JP���F�BRH^��NTRDJ!��R[��<﮺�5�&����d1l��x"eq�2�iYK\}Rj���5*Eno��"����>�k$����2U�X�)�PY����m����#�OB��^���jUU��3������=�L��($�*+�����,�R���6a�7�9�b��/ӮG��"B�����ū\�v�z�-�Ӝ�q�4n�$���kMQ-�9��sz���V3�-%�ZjYE��1�A�kc�æ�:��Ovy��dko��N�#bP����1�>���+��	��?|�x���N���NeP�����u���4��c ��ף6�F����ݴ��+z =�%x���Y���L�а�+���^�\���G�0vЯE�1��`c����HP���2|�}NC����~g����� ���b��4�K������׵Z���[n��R���L��ETӗ��ЙN%���"8���u��t(�o�����7���J�}�����׊���p�8�]	M$�D�t҈&6ڰή`�#ިL#.����%�4���:�q����}�'E��d��qʜ��69�K�\�!�, :�6>O�?�|@��JGZCw�C�Ġvte��A5�C���v�����ۃ�W������������?#qW�{�]���>�[[�<բX���x7�ퟀ������t��؏�x�w�\�o��{O�S޾��w�(uϧ>Bv���6��`c�;8E)�N��Qɱ�X��}���OX377���,�Kn��zDZ-��P{&�aQ=�&6Zc/�c��q���9�Y��f�����_
��h�"������ۮ9�Pz���?L������V{WG�\�Kȗc�Ê�gc�aIdlS,H2��~�nw���v�a
$]�IJ���*yg�0F�j��p���=��lu5 ��������JA6;�-���$�ʵ�p,�,�b��&=���Z.�K�Z��*Ö�1��X+�Km�vRl砯`��Q5Îf�`�qY�5)�io9r�Mତ�>_�Z���N�D}�aC[�$���UÐ�M�͡��F�8G��[&sV��)lr� mJe�&-l��9I��b�ֺNV��]!�i�S�sml���%͚UY�չc/�L�b�lAos�9q�^s-E��MS9-�
X���i�0�U�	@<���6�d���L�s��F�{sŶ�i�tT�5��<>�"��V˲�Ȉ*M������Ql�^6&���0p�G,;m.��>EA����:�F��
����T'��������n��i�_�}nl�Ñ<�\�?�f��<��/54R�~�^ϴ<�P٘�Ud+���ũ�Y���q�۬Uw:^/�
�W���[^_�	_�=E����޽��|��L{�Ѝ�@U�R�J�BgQ�,1����f!�&��D�Y�h�F�MNc������;��������|F�&.#p�� �(*@X���0�a}��/y<i*�7�{>�z<�2gϜ9����&[�
./�B~��v[��T���`O�aac��H����R���$oHY~�(���#�뱈��i{�70`qrK�!��$��./bR�E��|����ndp$ؿˀi�����P�O{6@0+��(��iW�����x���D�w� 6�� �)��U�dl��e�c������_�F_��Ӆ|�gB�R�wx�@7�����Aϡ3����C��ځ"x��nE/�TҦ=%>Lf�X>��r�磍%9��F2F_�Cp��U4�zp�j~&�P	
peI-�^����ԑ�
B�����v����4�*��!��'�^*P�y{� @�8xxΤ?��ܷgMY8���v�G��?�����nyw���E2E/��p6ؖ��k�����D2�L��-��l�T\��6��3͙��g=��`Z�5cw��
[�<��pb��GB��?M�KaM�ڵ�@oeں�6s��\��EE^��V�:@�1��\T��òg'��v1�gt�d�m#eDx�>`h��k�;*l&����7�jL�LD#b��k��������ga�s�봘l�3��%z�U�`S��WSJu�_�&�F��F�q���{�'1��9k�/�����/K��}�y��?4E~��~J��ߵ\e.�E%:����r�W���։?���ڹ�2���v��N�-���g���?�V�gQ�.~QB��;9��ݎ���oUZ��
��8�� �<�g���!b�;����Qfq}�;�_n��w-�[	�9�r�&"�009ӂ�����~�	w
͐ma  @�vI�� ���+���1x��퍘M�������l��#"5��6�0����wj�H���ؾ��,Z?��}cF �P��qZ��Њ�]7����2����#�4-�?�!�WF"E|�S�f/���u�>$o���ieaZж� -[�ʸ�����D��l�@���F& �����Q��p��}P>�[���$�x�C.X��2;��96�N�
QQ�a��>�cpg��X:�a���W�d�XN�К]/#��/��:�>D��v�?y9�ZɋMsX��I"F�o��x@�e��\k'1uK�2��}		<������Y�x����:2� �p�JeG���s�<(=��a�!���a��΀�ߞ1��rGh#p������A��Ë\���\�d'&�b�OX���拳�ǓZG����J#�«r���©)W��X�?�<kQ��a+�V�U�m.u�"[a���p����UF,��/�;H��h�0��d��k�kAe�T+\˯�p�[�����,��<B�u<�՗Z�'�>������o���Մ��A��E��-�KG/�WA���$�K��~X��x)X����ʦơ`ϑϝ}x�Yc{��КZ Y�h�n�sE�҇s<�
�KU �
�D5����]#e�}�9#>5՜z<Wy��k5s�����ޯ]��u�Թ`�$��G%K�\QpO��!u�ִ��g��SA^�M�W��s�]���/[����~�wGs��^�=(�w(�+����R�)qP,�h���Z�͟�"�����
�٤�F�`��l�:�"8���lF��0	FP��7+�Y��>�[$̉��C���pJ���.`gF�R����n���s���l�|��]�u$��wt�6�ɘ+�NW�{ �|��߯�(?B��o��4L�<��;���͝��`�	 ��B��o`�-�V
�X�M!�oR,���$��D뤣,�5�_T�0����d���sy}�l�u.�>�'�Yd=��X��'��w�qШ�G�E?��L��
�}��4�Y�?�ά\�h	K��-���z�v�>pA+b�*H���n.�
l�F'�X�&.\�*��Yoo~�V���F�=?<�w3ǁ"0H��~�XR^t:��;��҅�$yc���Fn#�Q\,�~36c��k�n���\�H	� �ѡ3�1O:��W���ī�2�t䓒���V���K�b�� �ݮ [�t��������=N���4ʦ��'p�pw��&�+�}S� o���k����ɕ���܂��"e��!녻�і����P	�c�y�̐������,�:7��:{�O�ֽ�Ɯ5������L�~8JY�^�[��G��{ w\��7�ֵ�%�	 �_�w7�%.�y�ͽ�c�����W��f��n��V1(�o�|2$ʅ��M1�<���V�Q�v�.���>Ә�m;31��s<c��X�n���N{wE� �<3��TJw؎o*I��r�7sQ8
�]ߞ��B�/7���Nk�|�&����E�zߟ��r�.��E��Īb���a,_%g�Mh�ġ��JE��n�iϯ�Ks'�|Bx4$�������ml����J��$�ρk�l����ZT6�������k�Kg[�DBI��<=m�3SI���7�g��H����~h2��u�!7\��Ԃ�0qjY��X�̽��ɔ����EO�)�� �m�m�"��'�����,�;��)�Bބ���F =I��
}�,/?^TGh1*����"(Y~���˽�O���}�Z�xo��2A���=aO�=5����5l�m�}ƎZe-#kmS�3���'�ꀝ��d�� �5��,&��^j��5�@:5���f[�'
#	׶��0����T�!O�YUwe��y>��j�흩G ��4s�vY�F>p����������S�9���е#�An�bL h�9"�GR�`o�%%&ꇕ( �$i*Z�M�.H;H��B��7B��`��ӣ�U<%�"�WS0�A�d>k����X�Fs��D����z$!��LJG��@IL�9X*lU=xJa&0t�� 5+�tT�~_s�^�$�>��NUZ�q����Ӱ8��=�&�P������l�Y�/�H�Iy�:�i�� D���߁ف�Q�EVx&&*� �X�^�-�$sH'$i8˜99{�7�ɨ�����R�*�\C�(l��H*.�+�����e��1�	A�h/�S$΂,{��ޘ��|w@�э�̍���.D+�f�i,���+e��Α�X��ܸ��0嘶���to��v�v�`��AN"bVx�4}`��Or.���C��' �lú�5���QOGb)j2�
yN�ܨ����8�jB��j���̡�K�����s����C��e�^����1��L+���ؗ�澕a�w���gao�>L�kΩ�6^1:�
��cVRMA�5Q���x���5-z��𨿨,�j��՜x�)�G1I@��2>_�n=~ߖ��苷���/#�?�(#�&�r��|6��w]�4�w�܃~��О�.�KܮK�~�/g��hd�v	�*4��I���+T/Ȣg}�u��+U؜���a�=t�$�۲��MX�N��]M� ��A�H&F�0B��u�5K���6꽲96����xF��h&��>E�&�����f��N��c�l��t��a��r��������T�>RRҌvaHȣ�,��=�Ta�@���{2�#n���z�;�p�Q����'�Je6�XV��yC4���`�����~�|��3?�@i��k����I��WR;��`f>���f>��_Q_f�����_R���LNI�������ɕp��{���<�w����Ow���I��s��S���<�]��9�X�sh[�r�H8�6�[:�	G�U+C�mB/X����7j�puu,&�M��ʐ��x3%]���Ћ�^�f�r�� oS�T�D�|,(ٰ1�!r86Ҭ�1	'�4�N�g��r���҈Zj�!�^,,���[""�Pˇ� `�u,��61�����[и�5�����~Y*���Ime�'�B�߶\D��c�S��4xڜab��>b8G��l��j��&������e�#���6�tT�� y�aI(r�4�ۍ�g65�)dbS�;�>8qe�^������m�����~ 8^"^���>+�H7��/)0�Uy�˨��#\���:�D�щ�i�'F�C�ǿO� ��I6�!S9�O��T	zh�Ҝ+�m',;�q�,cCw��I�CC����@��7�L�tn�-��1����i���N;����D����]9��g� s{|3j��s����7��`瀱|C@���} ᮳�KW\\ܪ)�3`�nK2l�8M�\|b>�	%�R�&b�^��*����=���M��Ot�ʼ�n�(��Ƞc�.:�c2"v�L��#�Q;�!��`{a6FU���&;�tĪ�=�\�R����Q�﹕�7j�W��}C����� r�
L�F�(��v������z�7�.{�d["�%���I���6��y���m1�f�T��+�š�n�G��t���Nk��A��ټ� �r��MP���o�V����86X�Y��K�J����.�\
63��� �z�v��f<�Ƅ��ۏ$�|ΖK��US�F;����g(�#�^mz�J_i�E*����y��j�=�ژ&k^0#���X�u\��Lc��#�Z��o7�7wf����:�-8��B�B~X%~"��A��yΊ�/�"��8��{�ۋ��xO W�!	�ԑ�rϤ�s�SFu6R���b`x)W���ilT���V�c�c������A��޾��}�ߟBx'S
�Y�����Ǌy�ӿCx��*g�g���e���瞤��O���1&4p�m�r�}υ=ϯ�;��[W�O,U�K=>�_����l��V\�
�C.xG��5�H���s��㫻�n��%�0�H���ϋ�QD>�'���OB���`���}�b�޺�K��6U��<�I耒c��G\�o�\O�5��a�F��. w�#mL�����ݭ���(R�����V:Ȁ�.��ՠ���:c�d��8��ujȿQP8��t�6)�2+��S!,t}��c�Y��l��8�O�</84��X��m�z�z��W�?�9ݤPX�>�!/G"�$���}�ģ���^�y�1 B�B���Hn�NI5@5���aT�"p�)=�ǿ�G�������WK�f�l
S����|��y�T�����.�8+ C���M��c��#䰉��V�e��M�{���[�D�bC� ��+
KZg���H�S���%�3�b� ��XƐ{���߆��i��[�;��eÏ�@�=����/1��ՏQ2�N��Z����]���U2�;�D{M;=��	*KY-\.;�Gx��l��X������D�P�R���� ĨB��I��eø��y��f�j��p�	TNf�8:�O.�TP!ъ%�����z�2'��:������ľ�G���9�����B-�����>�a�Β�Q�N{o�_�mY�c9+�ư�PA��	$Q�-�tɀx =�Cb������Z�����g�����CǊ���L�9�#�O���^�O��|Ɍ�t�j{���m����8�]^���g���&z�u��!��HSƯ���G'��pv-�bqi�4�2�硫#PCP��)��ʘ#�Pf=k�����z�?	2Z��O�Z�d:�a��6ȱBf�NΓ'��P���)����@�5�O�p����|Ya�O�?�C*�xuLp��]{2^���UvN�}�[��A�pF�2r�E��y�4�0Ȭ�^<�%�BB��&��2=�і�앖Ҧ��%:��Y�aS\oo��Z�c���g��!\X[  ���3,:�{eK=�^�d�}j���Y��^�f!��?cL���*m}�B��O��l�`.v����O�1�
�"�H���j6������6���ԺԮ%2�-h�dI�A���%VM���`��a�����t4�VҎ��{ߐ3��oK�C��w�/�OC��n�?�&�w<N� ���lv|�E�v��^�BĻ��/��5x�DCl�!���$A��g+9�Ԡ�g�S���Wb��L���Y�v�5�7���<t���8w�¬
C�4��tG�GM
 ���bzP�JR_�Y���]�ˤ?$�o�2����%O�l���q��L{#]4���������ޕ�GI�����|�XpMg�z�^��k�u��r-k�/�'�q,�57��1�f���'�K"�V]0�ߙ=�n�KYRfG��Į���x͌��5M�K �e�C�K�g�Z���k�F1���+�{�׫?2a�W�\8ͨ�Y!�b��TcF)JadS��Cc��a��'��7r<n`�#=J��$؏�أ��K	��/8�b6 ~�?�|��n�ĵt����tY��������A��/��{���m�<j�5�I�tEpZ [��)T�o�����-1#]:U����_����Dm�C���7��t��i.?󼤙�)Q���+�~w�t�z�I?����U�.i��\:�o���v1?��d�[�m�� �5G�@�g�������ɭ+^�I��H�w?���;�y�$t	�ONR��X���j���=��)*��}�1���������5��C�����y�Q�!"�I�� VaL��C��OT���7�=&��~��yf�,�E˾>p��^�zyE�`�O�?C��'c"��P�q��A���,LCǇIq���ҳ��ic��#ݔt��t�_��93y�d�<g�[/�e��K8�ݳR��;V{��{v�Z���k���^(B�r���7���?S�_j�_��%d�#��q����#�<��|Sa�	�P�?��[B�5�a�E��~�ĽE鈚�6�;�I��b�̽��-��7?n�7!��<��`vI��۵E��]:FM1e��x&�>ϟ����������J�ϐ���2�aخ~~ɒv�P'���`zA^18�q���J�B�;Y0���1���6�Ȱ��{9-�%�k$;�sr*#��5�>KF��L�5?�|h�����	��ǃ��[�H��V��a%��h�-2Ō��߂����������C�+���i�8N0���e܀k|}C�Db�d<3�g�p<�Q+ I�� `�0bۧ}����A<�@��{t�8ࡔm>o��[@�5�9���_��^���}�=�Ad,\��	��l��d�����I�{���	�b����0|���e�|��.�}��*#7df�[*F���^�,7vӵ�������LV映A�,j~7IT��tX�$(B~TZ����Ƌ��9uǞ*ke���If�>��@�ҴUu��G&�PYR�Qw��]<j����	�����m���LC���7x�fk�u����8\������B�ݮ��kV��9L%�C6�<�=�;[��(_0�6��'|�E�"[q������C���ޯGLqM�*��B�/ �������gR��AJ��v!]�ɼ�	a��kn�Y@��SZ�JϑZ���� * "�Ӊ`00�j��'M��� '�~� ���?�6����6���6��t�sv�9'��	;+1��no�=��(�CUE�Gt	Irc�{~�ޝ$?�[X�zd�p��M�7e���u@�Ol�|�S�� ����U�����{8������gv�"y-���e�idT���h����`�M��{��[��F��W}9�,��@H��t����j׃��L!�Ǹ�F�%���pQ�L�/�n}H��<w�q-G�����[�4�7V>/:���z^�"`�k��z2�;�#�&Cn���q�%�����I��6�	�Y��;�c�!Z;������[$	�(��B�}��i��?Hm�x d�{�e����F�x��:膦D��;� z&I����Ƀk����~0�k�R��(�PV}���������i���d�@�������M(�M����4��_9���!4�Ş�t�#���dpȿ�����Z}�7�;:������FB,⟡
�~3�N�,a~gm*ZQ��_�����G/�$ѥ��:�v��F� X�0���a	-���H�T��<Pl}�F��b�1�M�h���z����|�Yek�M�Y�rm[�xNЃ~��uɲ��[I�� 6ۘ��1��T��kb���x����wtX2Z�y�}��bh���P�z�A���N���ӹnfrg��� ��g�Eʙo�Z�P3Tk:œ��[Rz2W��g5X���H�f,�'��f�(�d;*��5W��MG�{������箣+����ǇJl��͠?���wJ����u���?�7G������7>�Hq�Iv܉�Į�]� n=eb]�K������}Ut�w����<����|���;[���D��k/��V@�^����{:>���������y��
$����E������ �l�#�8C,
���t�p�����K�rQpS��<��! �Xi"��|n�<Ę�;d����s)���A�����)h6,Y�����$-
�%.<�*�4��)ę�t�$�Pw�ڌm�ｂQ��/Ɖ����tUbf��w��]�&�fܮ̦F��v���Wx^_�ǯ����^]�"��EcUA��#Q�8!ajj�-}���kޝ+�T��f禼��8���۟�.�����)�{ ��Ȟ�!��r��˰��������,�Ǔ�73)T?�:��E޸�):8��A]�SLy_�)��_;��y('E��wg�:�Jb�N=�A�*@�Ρsԕ�w��*	�d���Eύn�h�n��L�̏���^GC!�.���w�JY���\��h��K���Z#2�'�py��E���5���}1��g���cJ\d�?�0�1Z=`�g$V��|�~Pq�}x`��^�%���֢��=��S�P�v;O_���u��S�ʫY�Kw�
/��������w|����d4��W(�شV���5�ʭ�/ߔ��AǷr~���O*� �P�v~��7�Kz���D!t��H��z�z��8v~�tĕ=�¾;;�r%"�����ɟ�(�F�[�O����ԲB8]q��T���c�=3�!�Pb~�b�_�څuؓ<8(�d��&��o{ѿ�]�D`u��]��c�$U�9	B������?/W���P�U��OB9=NV@}���)�
=�|����]�<�q5��%�Ƕa�J,o�a��$��h�,���|�[�|o|��)��2�]�Z'���E��g��b��$�J��{�}�:�[�BWq!�55�H6����D��:P���3��)��6
� x���H�`B��<]0��/�կ����[Xfۭ.��;��ҝ�$��k}�r�n;�����~jXA�;��v�1V�"U���j������*��V�� ���A�8�9�	h%|@ã�O �5��Ob�4yMa鎦�=�3,EF�t3����w��e��iҨ�	k�!  �)�㡬,�+� ��r��� j��T(|lvN��=��E��l��5s���1��)�awE4���Fw��2YϫZ1gt���M���\/�
�9&��z%�W�gV�P�F���Y�>X�߀����
�����AZ�?i��z'�����en��Hf&�
�\f�M���i�U�$��*�/���|TF,�"$T�V�"�ڱOX�j"7_y�{,t(���z�J����?g����\�Au{!s	������+) #=Y�X%��=�佦�O��ջ�>#�GLGk:n_�:��z,�%񦲩7f=9$��HAOL���&��m4��-?�%�Gd�5x�oy�� X#�Z�>�n�y�C�h��*�<����8�0s��Ui2�j��z�c��R�?��a�z#���g�[g�l�+ �mLl�`h^lQ)�V,�x��eWp/F%����WxAD7��Y��ud�N�{�-����D�a�.�+;�ُ���u젃��>�ټ.󗉙�wo�E3����Î�9Kr~��q>�ݍ	x[7~��j}g}��BY���]��OW�։G��W�W+$����J58�4fK��N����ب�ɛ�J������Y�j��	����9g�u�Z�$�j���J��TT
2��5�3�-�ʤY�\�Z�n��n*�MF�Vx��Ul�qQ͌��uבc�K����qy�K�Vl7u~q���%I��E�%}��W>�hn�u4 7�j6I4�F����C���]���O�o��޳�:h^�oyK�oɎ�z���E_��$�/+�'���b�]�}�x���; L���.�]U^<��ǆO�{`Nb7��oc~O����;K<
�I�f<*M��u�;Ke7F�r���G:l�M[�$^��'�$>���`ɁTj�U�Yit?�lռ���|0�
�>8�-e
�	�xbA�� �S���W#i�;�"�� �,��� ����n�jH(0��^��y�=n��`Z�9n�`r8>�����[�c�W��L�nO�Gd�pH06`<4-Ȕ���8�/{*��ǀ%c}K9ܯ����j%���Ji�:�/X��G�4m���ABR)�_�U7Rþǜ}f�k)vz��p���3}�x�7�Zq�ew�U�c82�7�fy��$�;�M-.g�������jT5�ޖ\���|�,�2[��V�����dՎ�B�h(�ֻ$#�F����5���Љ�Ԕ��e��5_'�e�4�r�sĀt@�Mӏ��Rz+�Ty���^l�j=)��V�P3�%C�&؄��������d;��Z����yɼ|�6Yyz~i�����R}�U*�[}�xs1���C��e����`"�>v\��%}|%�2�@�6y��#A�Gѭ�2��2���4j���:�I�'�'�����J:�� �a�A�r�4m~�՞8��������9N|h�� ��1��Y�����g7a�sC�߿����c�Ѻ�X'|��R`#��{绖38����c���}��b��9�z�����,�2�!�?����R� �*�201�0�d� V��@��>oje�(��s�\�"��Px`�J�4C
\<koR����i$	����']a� � ��č���"|0���7v9��Xɮ�j���A���ɜX#͖�{4Jvz�5��y}��XM��fT�q�L!��z(�b�.k�����=.��V7�Țey�wr(N��ƒ/~�#3#{H�x��F�Z��ޖ�S�K�$T��Ş��t#n:��A@/$r���)�F�9�v���������2�,�j�f{Id������Km"K�r�:m�Wѓ�"_�!���W��ӊ�����=0\��@��*�r脗"�����4;I�L�P��\|��fь�6N���7j��%�ɨĕ6��N7�Z��rYWE㘹d�dTwgښݸ$.W�'L����o�A��2��0�_L���E�֠c��Z�B�B�W�@��y��F	4��>���|{�ҝ*����X2�P�����,oY��PSI&M'��_�Y�Ww
�r�VGhk�U5��B�ߖ���)4�ja�݅S(olKc V@1J�<���ZRS?��+	s����Gޚ`���u�Z�Npbx`�Zs�ȨezcEc�c�0�|�����kJ�q>�X�=b~b�Y4�:Q੊>�q��~a\k��Qc���u?'ga�|�c��5i��qLj�����V��U��`nJ�Ҳ)r��X�@\���f�L-�l���+,0�Nr��|o���������|�ǎcY�*i�	f{(�
g�KQ��O@�IsxQ��nYw&���]�mჅp�d"�Sl�C�W�Ǻ�0�8Q�-��g�^�GZ7�!�M�UXi}��`Vq�6�!(?;�eʣXyc�	t�/�X!�r0�u���g>����o�� }ɓ��ްSG���:����	� h�eH�k�c�6��2lkRɡb(k�5�,�ᬾ��,l�Ϝ������D��^�&��l՝x�y��>9D��J|ӘT���r �Ƃ��̽�[�}:Ӝ��7���F�� D�A-[[��K
ʈ ���}q����%�9c�ׅ��2� ~p?ʺ6�G�) ���o�V0Ӭz��P;�q�/���O'�C}p�09��8)��R�܎��n�]0�=��|įF�}-�C�"����4���.�Q~�{Z�D�m�i��>2�v���CS����i�g%�*��(<�M�&��@}�@�B)H9��l
�9���S�l��\1��F�Q0*	y9Xlr�χ������Qbx�y w��Ve�l��
'&�E�������Y�fYF"aR�?:��� �4	\��'>]���y���!����oTՒ�':���y�|���ݡ�"]�C��T����U>� �]��Y��^O�2`W���s�k~��Ӫ��w�7��0�v'*&L�m�<,�tb�<�O*�h�$�i�X�{�#'�d��/��ig�<j��Z_1x��Ǻ�����
<t�Y�RK	�
�B����F4%���z3��a��	o�y�r��6d�O®1s$Oy�R$�_���7*�����$�<�%O5<���+�ϛ���J�_�V'��5��#ϴ�qcޫ��d}�2�X��XT�f=R,���A��0��6����<iƱ_�+�T��(����{��"��	��䤂�ʨt���2��#�{pz�����A2Z��Z��`�G�
*��2�2���%�s�a@d����p���Li�!��A�71��U8ր������
�����i�p(��?k�e��D�@wSRRѸ擫e�qH^H�Y�m���o�c��[��y�����Zw*^]���ت �Q�ЪJ�3�SX�q~*����O���E���[oz�X�����h��'�$Ȑ��e�[f��PSr�����2����"S��Cf���]���ە����b]�PO�!Sm���ڑS}��L�=D��qAs��5��5��ɔ�9��3����,=n�ٟh�����k�@`l�gR���wh���?�Ǖ������l�>��ާ�<Ⴏ�.T�����I!���3:s$욆�iA���TD��ʾ�{�Ӆj�9������"q�M��ͽ�B�۔p�,��8�sw*MO~��a!9ES����p�t:P6��� >@Lm�pAY�=&�Zft���# �k�(J�E`n��x%g�K����Bbd�Y�FjLԘBj���T�U���0�Ǎ�$vSX#ƃ�ݔ���ҜȘF����M�;�z3?�>��G����'����Ҍ���b����`��?f		��ܟS[�;d��U��^��4�VՖ�D��$57#�-;vy�x�k���;����+٘��O��훧��h�8>9xp-r eLvm&�f��=����0�!���狞K���TO�<�WY��mQ�6-�9��Y6����X�^�������U%'�9�{!� ��%�`z��Rf�r�
�|��� &���n���\ �]�D�%��Z� ,P���(�*!q�
��(�r�x��:�'�^��܉Z�4!:����[#DD��e�6�}��O�
�Yf�����f�lUl��:j�f��jTrt�Ҩa��$�Y����,u�JF���_T���<����7�n^�3���B��@����3B��.�;r�V�B��c�Z��'R�%�'瓬�]����!n���g�	R o������lP�E��e�rF�
m �f�)��X���YX�%Փ���%txp@�1IF.�0��0�LQ�=(p�,���p����O��C횔�~��a��A�c��u�R0���-�f:^�X������LJ� c�>^�+Z�b�s*z	�EB�;��֭�N��dlx:�� ��ƖlB�m�y�����:�s<����3/c��w�d���2���oX/d\��>�/�c��~�DQ�Qǘ�����=9[�v�b��Y�8�y�:״!�B�8R"s���1���xko�� ܷ�졨w���d-|�_W��r��}qA�C�<���}���v<�P3�W)C����y��k�^��$ԅI ]�4���6�i�Ϲ^�ĺp2$6Iz�0��1�6�8�26P��H��/ �(����(����3Ħ���HӔD�n��AA�~ϝ��Rw]8O���^:��Iyө�u��\�Ѱ�Ӣ���!����콡���Θ-��NbM弡�����3OPC-�kz��-���O��{wsoq�(w�b�E�k�m�D6�3�!V��#O�t�8�lc��DD�Бr1䉶�q�A�P�Tڵe��^���_~�;?�����x����z�	��/?��������#�{0�8M�,�lب��Nǡh���Y ӂ�E���ل�\������7���ȉ��1��gEHӂ�J�z9=���B�����Α�V���sJ�$�¤]���X���9/TX�1��
y���D1R�ETk�>�т��4	�b�uz=q̙{!�(^�<F���V�����j�7|G��u��껰�{7;W����~A�@޼��4xm�nehB�+8�U��C���V�`i���o��yس���&]�����i
+��N��
qv$9>�	��b�Y��cZ�!K�bJmY�1g#���bB�w_����來S۔)�Â�\�J׮^��W}��I��r���o�bt�� �.�B[w_bm�k���\<I$r`} �] ) ky�2�$"=��\t2u�Kr{�b B l ��k�DD��Kp�z~̇M X�%U�#�D��|��-	��p� ��X�B���)�q(r��Sl�A�!�;�\�J���.�-^��YTP��˃�`H�8椀^!@]Ѝ~�U��26d4i�^@����˸�.��8�	y��EپZ��K?wǺ�ܓ�@@
�3җr�F gh;�R�dV�Gq�]��!�u|�0/Ej��0}t����Լ�(�����;�~��䞥_@6���b���i���1tC%�\���C��X��_d)�����Ue� m�P9������%Q�X�qbX�|"<b��4q0>�W&��g�k�΁[ק�%�c�GQ�Po4�b8b�N3m ��Y>�/J6�s!����Dn�g�K��"&����9�׶r��A/�(�t��C���V-o��`8B�w쏘�0�ixwB��-���g��d��}��`�	�q<� �Ή��ᾏ�Ր9�|�X��~jѰ�B�V!.{�����1�I!���Z��1���5d� θa���9�ܣ�Ϥ��q�3������'��H� O K�T��h��d�>;?|:t����F!��׆��nz��_A�~۷�w������|�*��4%S5��0��IK ��G�s��|!P�8�.��CT�9U�	�2�i�/]<CgϞ�5������SO��{4��TS� ���:��ݑ��BZ���1Xk@�00?�} ��4�Q���3����0�3�ktv{����q�4�s�%���9Z�q�]����e�;��8f N{{{t��u~��ic}�F�u��$���R�"�ƨ���tN_x�+�ȓ���/?M7v�6���Q���؛C����@��)��k=�Dا���(�x�-���5���4ۿ���������}�G?����~_rB�7>�����>�u�`��E
F0�^�R��Ȋ��ؒ��O������ɕs:�%�=��M���t� �v&d���iʋ>Q��M�1q��S7���������JS�Q9� =xR�bb�6����`��8,~��Vm��[���A*�f��"\�U���7���l��+&	h}HQ�'���F�u-7��hi�2�D�TX�|��T��e`2��Ӱ^�D�8���A{���	4ZRQd4��c2!���nx���ɲ�� ��~)T#�?�g�1����{���Ƶ��{�:YΌ�?OZV<�T�'��T���c�������s��g���[�Ԍ6�<K��=�A�/���h@�h@O|�Iz���|�H�� ��(�CZ�Y����.H���s+���%p��	������ґ2Po`�v\z�dd���
��bߝZ�����p��B0F0����)��Z�ER����mC�b���Ĝ�;YZ�;��EB�$!H�xK�{�1���S�lyo��B��N�]�]�=[�N�/��v�r�� 0�CPê��|�-�	B�J��ȧ$v�-Xw��t=1|� �ʀ�:��~�G ���v%Z/FTOy�#]����1��O�d˒k�����$�br0k���Gbb�Cpr>�G�Kλ�O�ɨۉ��cl��͒g��}��ҶB��״]�B���>�O6i��3K���l.@�d#������.��C �)����n\y��	���7b_M^\��ڐ���i�1�!a�&��Lx��f%��:�Lh:��Y �_K��~�T��Y�A��s�=�Ȁ�/!>
/6t�������Dx!k��Yxލ�i^!yDNk#::�gC
s �}��W�&&/ �a>�D�	P�*�����4���� x2H�����<��&�n��D���q\��e�s6�=�뺱	=�!�8X�CF)I�,k�����?q�R'�P�8�2W�X�� ���_^}�?)�"���1��oK8Ѵ�OPB�a��4eq��c���5M���aoH�.�[<K�{�k��s[��D������?�ǟ}�667�-���iNv�lr�x$J�jN\U��fo@�V������}��O����҅�b�[D���g���)z��}ڙ֔�=�)���U�9$�>�/H��!�����/h��Ҵ>�Vv~Dq[��SCz�+�w��Az�+�;�l�3-�ᆐ5�	����iw��n�i�`�IM@�ٻWW���G�nޠ[;{,??s�:w�Z���E`�7iP�TD��c���.>?DѻG5=��ez��k��S���2�KJ��T!&�G�K��c=��� Y�L�F�x�<`�PY��
��vB������t��������G�r�/���o��#o��_��?{�~c���x��cR���^�
�kG�-��re�$���)�㜴�i)���<H�ַ�9�:@��9sn��P�%)M�g�x�>�[��ݱ&�SKY���"���q6!L��:~q!�B6^, ���@�?�H���6XU!MLR& \iªy���`b�\�8����k6��E}��;�ã]^�Ξ9��݃��eEA�ۧi^���@7n��x��8M��O֣�����o� h[�= zl^�ꭒX-���$d�g�����V Vd�(K&X ��zt��5�y�:�ءvQzw����D� ��S�z����d�,^���nHT;e�,T�56���i��s�������Ӿ0�&f�G�����V���=	z��C>��%�fbs�ݿ0���v,����y%�P��),�b�|1O�.�Y��e��V��u��,2>��Y����S�.���ĐG^��m��,�!K�Xq���Q����K� �ˠU�J���/�z�s	���c�ޅ ������Ɏ#cT���?��dł�c�)@��y��%0Q4�́��6�����w�{=��6��^9�[C��6��9	��9��\�s�c��J�Y��*k��޵�{}����%'I��gm���S�a	���['����`�$AH��� (������B
� k㾉F��X�y�ܐa#p��	�������x疯BI��5���y�vk�E�N�>́�oث��f� /쇸o�s������ߣ[7whr�1B
 G�u�m�Bb$��4�Gi���2��I���s�"�tb��钨{O������hkk��#RR�p> �G@���km퓍��a��]JJ찞�y��p�s&0��{8��ձ��K�����G��x-���W��X /X�!s%ǅD��hg����
`w�A/�``2�rގ���������Pl��^���>v���1.�ťd(�+@�@ X����h"A
H�v�Ջ�C�1u��!}�;���tn�8F��=�,��?�i����[��V�ѿ�#t�sH��$FQ`N����*J��"����=��c�g�gt��e�#K���|�w��wn1��b�DtX��<J?��E�<u�����Krr:�iYq%n��:����U̗�!c4o��܌6��x����7Лx%���Ktv�g�:<Z���!���'�'��_y��\�Ee�Т	� nHR�v�⢵T�Yc�b��%cSQ�*z�;�F���ҝw^����
?��3C=�8�٣�ӓWn2�r0��yCM�Qel0#���J�OP�+��'ƇWq ��=s�NomSY���gh�}�-�����_~�������4�_��%���o�]?��?�3G�{஻��͂k x�T5U���,x�,,�����v�%�QJ�`�־~���oz#}������4�xNY"�d!@ʶÊ�w?�}�c���)^��Fl�iLI���eI~��/>l�q�"*�Mܖ�� ��w�1��Ŕ����vT���CS�T�3j�9-JE��"EiQ?˩���&��.?�4]��<M�3f}���>E�.\���5"h^[:8���tΕ-5�MQF�l̓	�6*X��b�e�Zq{�,� *p):��=! `Ɇ_����3���s��7Xp�{��v�
5�Sjf�wq�}��,C�&��DtA�2S
�A@?�^�1/�� ዘ�Մ�.�2G��@���w���u��sj`������ <yò-�ʎ�̋.=�M㹄B~F--��! 'A�H�����! P>� �9��� Bֽ��,-�'�ju=B>�L�%w��r���t�������aC��R�O ���!�N�J.�G�1?��/&�A��٩��ϗ��;�u���sK�mG;��ba��_~W��� U0$6H�'D͒؅�� �,#8Q)Y��������4�l�.��N�� +�c1
 �s���Jb�}���{�uw�.=)ᠥGF,���LAÒM,�a(P&������ϫ�[� y���C��g*>V<8ȟ/�k�XQe.t���&	��(	R B ـx� =A�w�.��I��E���!��l��� �m�`dr�τ���h6�����⥔���-Nz���A�.��� �&��0R�:t�'��ɓ�"-��Bk���[3��_̽wp��}.���q:@ {�$J�dI�-7Wٱ�8�'Nb�nO6�7s���&���l�Ȗ��b�rdY��e�.Rb'A��~pz/;��/ �z����� �9����W��3%�+Hnn1�z!��,�J"�Չx"���>}	G�a(��fQ0�@XA�5�S�jq��҃ό��>vdjJx(}M���ܜ
~�]pݲ��`��F-o m/�i\�f��:h^�nx*�1�e�C�7x���z][�0ӠQc�]7�����R�v�'a��z-��1�T�A$4���'i�	Ѳ��6ձ8�t���q*ڎ�ug�Cys����l�L~v\-�ߺ��ʢ
���!7��g����+b��9>!B�Uq��;8��>�;T��66�4����
u�{���w���C�����F�J,(�G�4c6��w�5k�?�h9;1�'o�u ݝ	����qގ-HE�z��
5 �����,��އq���hh����F�A��D0J/�P�V�?A���j�r�zmO�������g�F�ٲ�{��c��X���xo<���yL�;���9u/���&~��A��JھA��c���z�e��j��J��R.�Pȃի��ߕ����صmvn۬d>�c.SÑ�)�|�8^:|���#]n>Ԫ��H���\�!��F�T��5v{L�)~f��b�]�������cx��>wr�ͫ���?�����%����~��S4ٽ��.Þ� �m �EǶa�(�Ј�Ag����_��o��v�`ƺ	\�w/nz������d�j7Z���#�-��|?~�����t"ڱ�vPYr$F�e���J&�Z���wgpl;�X0�7�%��zٴ�k��3P!�nToPP>OS�lJd�*�Ky�i�3�j�vD#X5؋��AU�'Ξ���3�Uʘ��B���AG�
�NmP�)���/���>��"�3 (�IY�6Qap��iA����A�LE��ʩ�O~�����:��h���F-g	BDU�zM	I?t[�C?{gN���TC5_D�R7	�HS&�pd�`��0��-2yLTf� ����"`��B�9�q�6z֯¾��BW��STj�fL@Ņj$}:���*V~��n�K�6lۊv��/K\���`忣C��5�3q��A�99���M$\����@�܆��w���,	z�Lje��3��=��ҿ2�w$Y��J¯�^��mp��� ֋wE}�D�ARܳ]	���__y�+�s�VT�Wv����wH3!�J�\���%K�Yj��G<�圸���Dp)p'I>��w���W�	C�\�Kq����
������ݼ[�3�_9�~���Dj�/�7V����0kz�ߛ��T��5���XQ�zg�b��������GBPk�K�X	u	�f�J~�6-[��9,8�;����;Z��9���=}M�L�T`���VӘ�Y��@�T�db�+HB��xϪ>��[���"��-r0e��: U|�5�̷�֫"!N�&�4h�(�N�ҕD�B�
��_�������P�����^%�8;�B"١����G3�VP��Z��:�w!o��`H<�� <j|�2��)ty��*igF�?mV��!X�Ph������N��V�%La��\��"n��!|g��g&��?��v�0�`��E(�)�2��+;�,�1	 $��J���AC�V[�A�V�Pzz�B�\D�8ʵ�&��2���)@����NO>����ќ�9�W�B�xN�O&����I�;����O���r����0��������}���җ�� �}�O�{����3�����/�1�u��o�f�-4˸-YV��J�ɩAމ�3���-�5WQ(Vqzb���\�����`:SF��17Wk�C8�D��}d��j �i"�i�VȠU+#�c��Q�{ׅ�x�6��I!�"m���Gq��)=6������ؙ�N�2�2�'�?�z�\PJ'��f�Ĺ�j![.�ή �lIpnӜ�PO�Y�>�Ԛ�d�'�YF�[�Po{/؍�����۷�w���86Y����ŷ���I�gȗ�1a���6�6E9_�A�
�|��R�H�\}�mۂ�x��_��3;���Oܶ��_��2#��?��+����O�x�������7�r޽w-�?d�A���d2W����?�o��C4�1��Q����w]��/��R!��%��5IZr0���`�<��!��'ϡ��@$>���ļ �=d!C<�\f�$�	.c�Ȉ��nA�"�����6(�3��MUD�A�� qg�2���E��yx<54*%�s������n�F��<~���̴���BI�~2���Bv�"%�B��w�w���I
����"    IDATIt!O"�ę��#��cl��2mJ��r	�ad[FUK�9�47T���Ȫ	�h�E,�i1���c'�xf�lA�87n)1�'i��]�r:\,֒�/�
��L��觀�I�j��!��2-%׽�twczvJ$��AW�R�$.�ҹ<��Ym���Z֮����j�w*��j����0��k����X\1Xq��*��	�J�y8oo�sfxo�p)�/��گ�נ/�T!^��k_�<\U���b��̱D�^�����_x:�A#��5@l��.�|��_�A}DE��Ļ�w�7ᷫD��!Pm��/uf�ׂd��,���s���(��2�{}�,��x�qj��\��;��g�y���H�.����I��^�ڴ�_�ߓ������R���������		��U�Z�ad�n�~�Z���+;z�?���r�l6��N�����B~��G\ �J(?�zK]��"3�g���t�����O���'I��Ƌ|-�ZS��]<gR����X@����ٌ��B:��ܜȓ]�$�����Eg��+�1r�X���L�AX�G{�l�+�f��B�N��<f�&�P�B� ��5�C����4f�^\D1�C J�ZL :�{�9�@�ܢ�� 1!0P[�rF�K{�t����b�H�֭�b�KϿ�N�:V|��5�&�$[����!�k(`:�ũZ/� �	r�� K
Z���T�*�%����4��"�,�ݝ��	����H��HX�=����l�F_�b�S���F0G�&P����gǁI ����u	�zo�������P�;r 4��Š!�2��3�\�ʏ�k��d���S�]<���.+ׁ�"jo�<A��,�GN���(#�(᢭[���W12���8�u�w1�0��/���̧�k�J�*�&� �bx� �(fq��YD"1���Q����5�F	�)fpz�,�?���������<*M/�7nC��>�"'�e8�V0�J�:�h�Y) �:B�*J�9�$�سs>���{�ZtG��r�N�A%���O<�7^ۏ|��b��Z˃�� �y70$�/	��xP�V�-Qn�Q�7��V4��z�ZEB�H}!�,B��'�@:�Wǫ�(#�[�h�0�ߍm�7�]W^����80����๗_�Ͼ�����}���C�/��/���<2��y�y�z��� ���ء��?:�{��W���+���}����������o���Sg���n� .8ob�&bl�0��ߐv���|z��\�?�����q4�>����q��c�7O��f���*\(�p�(�*�c�ď|	�FB�h�C@��!�Y�7�gS�1���nx�2A��m���Oh����׊���Z�~o>V��y��i,��^��%�C�F��A?�*[����<�3�L��02|�ή�� �x��Qk�-�7�@(��?G,օ��at�E+�o(���H�n�W�h����B�<7nHt����d'�洕Jă�H�'�M�Q����dB��ݭgƄ`�3/��-��h�=eR�C���['�@ΰ&!X
nY!vf1V���R]b��hPثUT��o�����u���Y�,�����S.y&�j��ʠr)�uxj�q\�O���`�ݟ}}zg���
fx	�j1+���[ɺ�%�qm��|�ex-N��(3(����b-�g�m����%׽�\E��c*Ӂ%<�6S�I���۪�Z�"׵�kc+�.! ���Ҭ'��Z�T��Q���D�ni���V��4�lR��r�<+�U��ߙ���ǲ����0�<^��!���<
7s~�iu�)1`�O�� �V�F�w�k�N��D�����G0�����Z� H&�	��XԘ=;_̼p�� ^��s��C^+���m����I-Ã��ip�vM(R5sS��k�$�J*���I�f��	���K�� �s�^.�����"����(�"	�;ܼ��#���診�l�O��xƣ�'�.qf����W����Mɟ���b:���Uv�\�������:�q�z�^�U���p����oFc*�*/�7L2q(,�b7	vy���(gq��+IpI<��n�����|r��8���/ޑT��{&ć"����3|�/�f]�+U�R�ཻ3��7!=;�g�yF/
hpn��G9#�@4F�ZV"���$�����$��Pz�)8��U}��W�[�v�S�|&��ǜI]*���8t!��Q����(�s��!��GЙLi��;�	�013��^��N�����l!I��&����AK֧���
|��;;�u����A(���c�/�P*V$R���£<X(���IX]�^��1���	*d]���7�=�5�>2 �W�?3���t�pZ*El�W��q���8|�4��ޝ8t�0.��|�S�Ɩ��xk�1<��#"�_w�5�������O�M��}Wc�y;13��$��؝��S��Co������019�3��X̔���h��(��hE:�
DPg"f�°��"�&��ڕ�ߺ��&\�qF��-,�6?�o��Zf�G�P̗04�����'(�҅�d��:8,2�d�T����͢P-#W� S(`!��\6��LN�B�!S�r��l��\�"�"qd�9u��s��
�����p��ׁ�G�$��N��o��_��|�'�SB�Z��&U�
3��ٿٍ�2W�#������,��g/ٶ�/>wӥ���K���g������ppͺukї�#�E*�@2G4��UCW"���A��c.��/���'O!��B��@.W�ڑ�8��]�Ivjc-䲠c#�]8��|��S�q�C���'܏���u~��V�)�F��M��i��Zx����C�Bh�.T������R1�z��Z��z)_%����|!���
�b!��&P+g�!�0�QՁ�W^y	��4��L�%�����#�CzqYV�8���K>�����5��$:�=0����m��0�v��
&�"��͕)�CK&����P�++v��X�!P27e��
*�p�e0�M���/��7_z���ޫV�9���*�
��X���A���LB�T2T�
6��ÊR�K��
�``�(n��&D�b�MσF��G]e�\m�^��v�ו�ʯ��ː�Q@f��qwPSq[V����8/%���d������3�)֌�k�I���,���P0�7s���@����Y4��8930�O���*��� 4�%r���6 Jx<�:�+�"]�hx���DQ
�X��#�x�ҽ]�9�R�"�3�?�C�P2h�[���e�;q��Hu���]'��u��͆���ф��b��`O?�-��u���Y�y`�`a;Kl'9(SR��͍�G�5߶�X��6�v~�޼��
�M������e����C���I�ҐMH<m���9��;s�I�3
i. �j[����μ�R�1�� VKɧMd9^"��(1Au���.e���(���"9I+(`�^K�w�1��7LZō"&���A�#�;�c�9t����i�`>^���T6/�J�V���5I���z�T��j4|~]��':0;5�.1�><b��*��F�C`�_�D�TCde|��4*U�6i6F_{��"޶|m�y�~3�$�l��S�a��N�ԅB�K7�~�u/	%cXI���'W����(�Z�*1�}MNN��-H$"�م��!�T��L��Պ ,�/={M
�@��ȢS�^����P�����Т
��-��?�52dANґ�:Z��: ����p��{�g�Vv'Ѫ���;2dW����D�v��k�rUr�)
z��(�S��������VG��]�v����E11�ų���?��8:D:Ht"_��� ��㔙��j ��VDe|��}�����@*��!�~�~dE��s���p_�g�M���	��P��1cµ��d��=��Bѐ)Z"�#�0����l��Hg��� y��?u�zE��/����}�Jg�ϟ�9�{��Ţ��oæ�k��/������?�
��[���[��?}���w�N�q�m���[oUru��I�b�Y3*��'p��	A����R�3�b��C�&��������x�	�Y���m��9�PEg���m��k�e�0PΠ�Y@{!���$r��"
/��W)^X��xB2�{�L�#��v�����B蘩Ri?*���U�(��(q�PF��Ʊ�q���~8~���D"]��y��_g��5Q(����[�����`����*f�|�����+G�&P��P��W*�MO%��LY�%4�Z�[m��]H_�q�/?��������zu��C�}���>67����v� �ѶT���Z"��VB?�����|�3�Huw!�J��<3�`ڱ-�Ѭs�-+ �?TB������@�cH�Cd�S�2\t�:<M���!?H�����9s��k6��Zt'�ڐ*�4rS(��\ *y�B^$��o+Ȩkf�,�!��d�H�O�^�jE�l�d�b	_�Rֽ�C��F���`�_����DiV%�w�D��#X�q.�{9�mہBӃ�s3Ȗ*hQS�c�*�_p!TM{2�ep�GA�,�me�k��t��N����_�th6�a��~:�&����o%~ߙx�j�H������θ@�U|M{�%"��`������RBp�-7!�����������^�eq-���AȚJ������vMlB������T�J��]7��V#-��7 �=?��*��Xղ�2��T��}3�bgȨo���#�J��l��Ir0<V&]�@d,�t�c����$0�#MG���*oL,t!\��|5�pQ'>�ڬ�lF��FU-{����� VA�#�Ѝ�Au��S �b޶��;� ����J8���~�� ���Z��2��`��u7�ҬgU�9^L���P6n�����~T �P�.�^b������U��2,A�ͭ�lӡ��Ս�<p�flAK���6����I�)s�H3������r��3�3a�oeB��v@��Ѩ���2�% �1(�d`��$��n%LB;�VV|���6	����O�@�! n�td�cI�-�Q�	[S8��h}i-؎�2*�_��sNΔ/W�dy���[35��`�<�X(
Z�f	�X}=��1Д�G�9U���K����:H��G6�E�X��S�呞�E>�E�#)�p�3��U�"�P��/r���VrA\"� ^xoJ/��.�c�g��q�@���8������Ln�߇���I����Z�H��78 &|f�F]I�f	j8^�ȱ���uV)��B>/֬��/^{�eL��1�k��NX$Ԗ�f�HTѮ��،���^\q�&�l�Ƨk�i�z���@`-����9eJ^.�g�yw���YY�O�;j٨��'i]�E�����?�2����8<>�H��`TYo�K�5{1;V���F��������7��2�i�;ͺf�`~nOC�7��B�Y���Jf���"Dl�3���pU���_Yj�^l�ǟ�#�>�#i~����-7}�>�
u;�&���a۶mX�n�{�E��?�?*��Ƨ�w��c�?�o�q��������jt����:!�`!Q�!�0�Ο�?�<<����'x�WQ���O����ƫ�9��QDeq�VW�ކO�|.޹�F	�����<�
:�~���Dc����1/��j�e��m(v�!&�"i�}$�ý����ڰ�ܖt/�+�ް�;�����4�x�U�]�����MT|��J	��s�>}�2�1\��qۭ7`Ϯu�xK����^9x�h
�ҥ
�ݨ�����1Z%߁�̞:jS�nW�����n�������#��ï]���~��3��j�Q�@��T�I�X؃����^�wm�&wZ*1��8��q;\����ԼA��L%�	A"C<F/`�<��|�G����E8�J	A��l��4ʁ����w����J��uL�{������+hיT4Ѭ�[�F97�v��-h�R���"��J��[D">�c�L��[jʕ�Yͬ�5[�S� 2���g9t$ސ�Y��ڑf�{�a9'3�+�Z@�6���v�ً-;� �H��2��%��X��$ܶ�2���!H	X]t�o�1�����E�"T��N�b&��'N��+�#I�:�1���؂�Ky.�2n��&n��Z��KL%��Q�&A����:�o��T33�tc�T���7���/+��L��`=���0��j:-�������d魐���Vvڴ�Q��!/�N�B���3ash�."���	�2�5��d�,J
��ŐNB�C&4Kɞ��aaF
�D�RW�kMs#���IV2�0dp���ҬWѕ�𴦅nA4��Ye�aƉ����)׺�L.���v�,I�-w�J��׳5�!)�����-CԖaΗ�[+�o��(�g ea7K�dU=˷K��@�ڎs�v�%O0r�L�Y�6	2��m
.).���t1�<��t����t�򚨁Oe*cH
�8�R��ΑU&����2o[�3�y[�+\�uEe��f��L:8�Y!6��Ց�\3/�DMV�U�5�-Wp��F��5���i�b�=��HH^<C̼�uj�9E*;&@����,��b7j��M�������kv�:�b F1V�	��z�:�
����#K��٬�WJt!.���bf✤�׎���uk�>�\3�$���P���|=�C���B�X?�ISٰ<\���\wN���>�s��U.�07=���iq����.�����l� �P��H���,�*9Ƅ�r��1�7 ���c������t�?+ۂ���Kч�|��Y=M\y�����n�e�C��:/Y�[�k��f9�5��|H����-�����ߪ� ��� ��)I�۵I��X��WO�������W�������_���;`j�bA����}�6���b$e�\����<�*�
�'�5ǋs_?o!�=����w��ּ
*&��kr=(	["se�z�g[pōOfp���kwܩ��?�">�������R/7��8�5�n�3�?���D�q|��Ob��]x����;��1��cþ}�FwWR0p���v� F�x9i�ZφJ��ߞǽ?|S�|�n��^T5��_�h�sH۸x�z|�kq��;�Աx���Shf3TH�H�B�X0)�U�Z�JE�$�sMG�q��uͽb�B0�h�'J�,����ɇJU�H�D1��1�^,�#�x��i�J#Wc���o-�XT,P.,b׎M��-7��W�E2
<���{��819�L�^xC�u����a��>xCDoTD�Jhff�m^����=�{߾}oo�-��o��W�!��^�����f���e�4X��P+���o����>tûq�17>��o�y;w`͚5p1��ӧ΢Zm"O��d��x4�v�Y-����Ӈ����l-o���	�=�1���:2����=L5�A8�xe��J�ê�D�'hPzn3�c�ΟC�݁v�vٙI�|�%��b>�ba�RA_K� ���KRTGO�D��>��bk�/����l���i�l������ڋ�T�p{�B�<ۭ,�%1zޅص�2$�EV�Y� �/"ޑ����r]lZ}iI���	�������Ot���r.�srܜ<{s��A��JMʖ͛�9`����	BV�
)P��9oڊ�	�����Z����5���Ϣ���#�����!�gq	��C��w\�rh���XrKfpo	�a��Ӽ�$�DUR�nW`�MU��4-{%Fݶ�e�D�Z�vl]�<�B�_6�!K5{]D�8H�Q0נ`_�|��8�����^����B6�AC�s�u��8N��t'\�k K���t/�ī�U2���5�K��)7�v�\;����DR��5(r`�6�C��V+�I7�YZ·�Vf��������籙P���R;P&0\�x��4�A����N+���C[9��)w�T��z�1 5�����    IDAT�ָH����d�u'����b-Ui��ej���r��f&���|�����Ӷ���sLE��n���bCX_n���
�����̾�=�R!�|�~$Ti37�N��`-Ͻ��d��p}��t�h�5�.�8s�-u(�I��l3XRUۨ��9� *@տ�:IX�{�p�x0xf �qd��u����;�1_���s:�]���,��:	�60!i��Q�Ǜ�`��&=�?��%�[�o�1���3�2�R&j�~	r	�k��%����(Q5WĩS���f"�?�
�7n@G*�t6c�&c���֒�bR���3G��Ǒ�19~Zɀq�6��*蒫�"
�^kH��Y/#�8��+���o~�\�szha���T���<���4m`���e��@�L]{�LQM��oQ����}��mE ���-�݁B�{��¿�y7�{m?��$"������_���:%t�|��O�W]��}��غ������"z��Ou��J�	[�w]_��.Z�n����&�v���"�l�UM��U'��������G����u%3_��qۭ�U��z^䌁q>���q�]w!�H�c���܁g�}߸�N�9|����믕QeB��Atv&���i!��h��ٶ���8�{��:>��'��T��� ȳ���6�*�q������4Z���<�����,�QX��3��nkr���NXL��$�ٮW�*dr�۔4��4�;����4�PYT��ĺ�ѳqH����px*�W������<�m��$��]�ɟ97���p�V���[pյ�� ��ٓ815�v8��B�&]�)y�H�>�4Z5ʙP^,^u��/^��?��o<���� �}_��v�z�;����^��,j���
�D#�c�;��p5�ٹ'�<���86oۊ�n��*��~���uشi�	b0���H9Ħ�՞k���(�}ߋH���'���	�&~BnĐ���a�sS�;�!&įS���*����*��8��3'09~��<Ъ!��!4�]�O�XXB��E�VDoO
Ѱ`;̠�\|	�٣��?D�R���H)Q��h�ݡ����ge�a�K������1P,�
��i��.ր`���u�E�y�%Ȕ*���7���#��\mV�e�`�kӴ���R�ȯq���`=�^�b��)���їH��ͣ\,b����8urLwڔY���V�]�@1M�̸�M�X Kҵ�����
z7�ƍ�����ŜƓ�(iH��WXr*�>�r0m�M�7��`86 Y�t�A��p���,��@[�J�pӖ@�Pђ7I�d ��]�z����[	�=(������%I�G�ƃT$TV���%2��Ms�4���{z-�[��\b���V_��;e�e��J��+�%F,��yZ<+��̸2�p���I;v�P�$9�䏁�8&�6c��t
�������8G���-Mpv�l�$�w,)�Sֵ�`�9,���]���=&rp�LŪr!50O����ɱ|f�1�6�$�h;�-� 3@f�j�TPl��1�|^&@1္fC UR�"��7�ҥ��k�r�f�ױ���W�o���8^�Y���j	��R��ƵՌ9����C�y]u���[#T�`*��א�]�ŭ�L�nI����j=߇��*2�`jX���;t���3�)-u
;�/��$OL�L�����_�� �f�2'�g��c���A���b��/T2���vE)Bx8'	%b0� �&�م4�S���� �Xyg�J_YI93�\��ĸnq�"�V*:��;���:7�J=]�K�M��҇�l�Jy��EB_�������V�8~�8Ξ�T�BO�u�ף��W�b����N�M�PdSA7E�#hˠ2½������z��ob�M"����TV��F�|�VQ���ĭ�₍�d�.̹NOL�E��h\�L3��[���-���{��[�d�f::���lAG��qGV��K$B����b/�qO>�"N��F�ƛ��9��hI-��x1�c�{p�%{�q݈����Y� ���in�N�=����O�+�`G��1A��ipn�+,?��6�G��� b�{I���b������q�=��|�w>�+.�Lq�$�QtĢ�N>���p��D�>��ؼy3�x�	�˿|]	���8.�p7�Eͧ��Y�)���,��G�`����	)��O_=4���y ��?��/*�-�_�b!OGz�}{��.�h��gQMg�.�� ��C�vҾu����x�D��Eaw�|�tFIǉj`��>H^6�F��̹ �'�0��<^��J�E�p �nt��El�Z4�]H�|x��$�}�M�9>�s�"��I�}4 � ��Q;�����#زm=h����/�Ǐ�S�22�M/j� |�*������,�B��J>Oq��o��/>�����J��_.����'_}���~��-�?D�,���|N-}�
1�����	�����;p��q<���l���!e�?���;y;w���/ޫ�/�b��i�2S���X{���y�jI�{���iA��K8N _����$_V��˙,�t�:�C��F9����4
����;����y��5�bn��,��W�f�jQ�W_��4:2�v�������_��~�"�Tj^��q)�Y�W��yF�ITT���2��&��T�%�H�j��� j���ـ=�^��[v`&[D��@�ڄ/G0�6��������tu�+�V�M��3�[��J��N 7�FG'g�073k\���F�w.bf.r%���pMA�	�yo�d���0�>���l�x���4�A��Krft��B1��q|9�#��%;���`	+� k)X֢3;�g^c��|�¦jf!Ive��v� ��iC���� ~����5�H��y����n8B�����l3�,KRTG��\%R�����E�b�q�S��A^l5O|�d�׼�U�w$	�΀q 5��. fE�����@M�V�M��i�s��Dݭws��u@:���zNrrt�4q�5���بJ��J��W9�I�����;��C&q2��|�$���V?��?&�Z@K��%�}
n9�L�m�u���,��5�ƕ4M�O�p���#h���@]�&�A�!a`L���J��3�GH�_Lt%�h 5����re��r�YL�8�uг�ʄ�ٲZ�+����2$oY�W�c�^�"�d��o�7抦+�D�A�a+~����{ɀ���Z�Cbp�E����%�9gڭ��E�-�Z��T-�D-�-�%�zf� �q](U:3=-��t]�j�~���dD����>�7�ȡ�UgF?_�������Y�_h�y0���J���N�F��2�Cuu�Q���8��-���g1=7����p����ST�r}DR����+��*�R�Pa��'O`�̸$7�z���~�}J���DF	�<|��2ػ{+>���ʋ�#�B��+��_<�?�3d���]�c���X���7�3�\	g�F�#��ML����H ���OglGGJ�q�K._�B.�*�<_��EL�g�h�JTd@�D�X@ Boo?������ٹ�� Z�<֮Į��4w��[�Ց#���q	���l�ZX�bw�	�(>+)�5e�f`�AT�U��:J�%��z�vh �׎`hU��ګ�~��e|��㟿�m�Z�_��?�����1����2�ڹs'.ۻ�H�<�4z�!͍�ƓO=���###x��އ��^=t�������� fffp��1���P��]���oņkPn ���~�<�Г8>6�)}%x��J��
�}�^����"l��'���P�PFu1�]�g�aanV��J��&�����1�5Р�x:�������URvމ�`�6�L9P��Lg%ǌJ\���=���"ܳ
��UH�ـv2��3s��z�%�Y@��T?�&��J�ʅ9\s�.�Ƨ?�-�m��l��)<��a,�}H���x�:DyS&%�*�^.�k�F�
j���˶}鲿��7~�:~��|�G�S��g`���0ғ��YG1�I��k��������ә����`&�X�v�R%��{�ǩSgq��Waυ{uP��EL"C$�/�d����w?�\-����J��k�
�~�i�����;n�����
XUxZU<ĕ�P��`~�ʙ��'P�͢]��4' x�����Uf#T^i��ҷu�F���|�׭!���ڵ����/���"�F(���E�D`f�VI��_���n�i��Y��F-[�m���n���VP%~� |1�ۄ��}-��^d*u����~DS=��Ƹ�V�]����\|��x"��#��cqa�r�BQ�!蚥�������@A���
T�[  �9�E���
{"���xQMm[��?x#b]���[�k�j�j\*=���4*�8|�r�pڢ*��p��@�q��� �*U�8c=(;Y3K:���
�S�Q j!TQ"t�e�>��Y��j#LHxi�����d�FL���n�%�1�v]S�3w`����dX��;��S++�Rlj����O��E�);n�ȧ��:�q�������������1
b����Ʈ�<���wMS�3I!CF�_*�;�=�Q���$Dz/M:3V��0)�	����ov�̼���4�5�(J�aBOB�W�53F��e%E�OZ�������޴���o8��7^�:>46��R�:�ۦ2�H���=b㍳����{�"����򐴿,�ʤ^�DI+�,�[�e*0�5�X�XFn���|�0�|ZO̳�z���	��r$(�5�9��q��5�:r��b����٩k����h��.$��5�ﳤr�]2��k���pȯj(�K���L��~�s���O��ՙ����s����Z*����@oo��)�T��p~��b'�IL��S��o�5[�\k��Brε�v&��ަ.���{a����@	Yp1����Թ����{��r�q�|Z��7J삁)���#f]��Q��R����^�u�p��~��ҋ�Dp�����׋��8z���h&���"Y,��/^+��g�|��U{�C����o|���}��,w��hĈô[��X}5�K�i,V��c����!MD#���-��U�)t';�����WG���9�:3.߆��U�P��3��Ű�k��YuRXt$8M`frS���7b�M��<���sҥOuu���Cx��7p�ܔ<�z��DE)�\.�䧠�ʞ%�1Q�QY��r�:Ĭs_��k/���u����ޏ�^wS����������@�� ���S�_�/>�<��>L��UW]���������S�q��Dc�޽�d=����o �m�&���3gp��a%�?3�s����'0;7�����~�38o�6�����ϼ�W����YJ,b,����n����lH�4�3��O�!��U��\X���4ʥ�ᇶ���C��DWG(�Q�d��kv6'�Z�P�`��L�ǂ�1��1�-�:�斗>G>��X(ew���x
�~t�[�Ъ~�#1<s�z�����ɳ����	`��)�3c���>n��m(6��^}�?��fJ�T�(����\
uL�bT�O���6Q�?��t�?��y_��#��z�C����W�!��x���z������÷} �F{Ů��I.6:����q.�cH]W>hW��]���Ӹz�u8＝�X�)W�c;�CWi{���p���a�G�sTrج��EI� ����UvV��n�̨k�<��,�R�Gf�,��T��(-N�V���>�*<͊�Y���S�TT���^TC�y�Vlڸ^U$��ذq�|�i��������yD;�$q�/�u��d
�`D�kW��&�D(׆\э۪�a�<6:���]�����=�a�y�ETI�(6�H��B$�R��V�T��L��M�ٔ.��p@����TK%ɷu�b8}�0N=!'�v�h�7�l��`��a̉o�Lpf0�GkTvX54�!I�5J��Ї`��M���� �bfaVs��j�p��.*!`��%��GWS��?�
w�&�w	-S��B�x����-��b��m�s�<)��0�j������-m4��LB@�G�8��JH��R�~��eV��aBm�n<�l���s�t���eN��u��i��y�LP˟�Y���J�I2���!����z��BlTlx�.蕴�%�

�6e��:�	tww
�0unF�:O���@��V��3.�:�g�劬�>�:�ҏg"nȶ�NyI�٪���
���{`����Ӓ��0жr�L��y�?��hҗ�2�$�R֒��ȅUەR feu?��sD�9�
u��<Q��J��$�T=�z<��YUeM��`�
9�>�O�pwXc��%>�D2�	��,ɫڠQ��%\!1s�&�������NV�KV�;v~���&6�Sj:�ـRN2T2g�����ʃRu�ҵ�j��U2�������g��0%�	G�(����3j>�4o�4k43�]E���ӫ�K��P�T���Ic^[��x��<�5țb`])��	g�:��o�ǚ�k�#f:���@��s�%��;�da�]pI�SR����XH�a	�)ؙ�f~��n�4~�Ҫ�6jǳ��Y̩*�jd{��QB@YI�v��w0)
��"��r��0��	���x���T���]�a��*�;�cG��D(@�L�,v)X�$j��.ڵ��qͥ;�!@�%�����q���Ȥ.�WƔժ:[�$�I>l&�{��	��6mڄ���j,�ϡVXDw'��Wc��(��T�e2p��qIx���o �Q��)��@0��e1��_*U�Q-�0v��z�5|�C��ګ/E49J�`IA��������#�}�lٶMEV֙̜�B&��|wɹKh�G)a��m�ڊ_���I�k���}�b�P��O�}��lNyhjf���G�ڷ�����տ�k����'��?�1榦q�7�K�Et���V���A��E�V�U�\!���i^?�wzf�<�({�	$S=��>�իG���?��O=��c��j����i���9�Zq������?�ʘ;vD݁��Bu����E�i�3�H=����)rS��E(ͧQL�ѪVA�'��*{�$Kp�o!E�������&8X��`>�mb�u�E\�y���GD,���ѷm+<}8��a���\o����c�(T<�T�8|�E�������+h�x�W�!8q.�l#�\��"�_�X�8Y���5R��j(�'�n���{w�Zu���������c���W\�/���݆-�0\�٘�ŦQ-\��&�4�v��q ��N��{��Թ9\z����Ke��:��d�����7�����^��2�`k�]�P���rW$��"X�6~WY��"ul�S�� ={
��g�eQ�L����t-�iVU.��$�7�U�;:���f�n��:lߺo��*f�&��1s]��s:�z������ÿ@"�'�P$�\�dZ�0�a|�R�7V��̢`U��!vho^j�տ�?
�t���b��~�^��k6+�],���E ���aݶ��8��L�T�W�oL�
1�ԋ�j` �N��ēx�����d�O$,��0���˶��եo1�u]�[m�#AaQ����2���Xr� ����s�E8�0�s��j�졂Zu��1Ն�P�E�����S`Zւì8,���$=�*C��$z	��l�J���΍9�I�ɑ�M���v	MP{���!X
7�b6�d �l����r�r�*��ꄢ`H�`�bQB5�ë����EB�t�h#�]��4��:􅩧�[k׍����T����,j�*t~��Ãr�4R�jUt�m��ݬ��M��744���6�^x�����b�3��Y� յ�Le*b�?��{��'��|m��%OG��B^�cQB��H�;�*�    IDAT��1=;g�R@cC�N�'J�2�T�'�S�8�kv�,��c�D(@*�!����I%�D�[�!Ke��䰼�WX�+ԡ e���Tu���J����z�s��Ԥ�\�Ŵs�6
�� ¡$;����y 9Knd1ZUS&Ԥ$�uW�S��]1&��Uu���be��Q�,�=��¢QNa��j����J�}����I�ϫₓ��ڪ H�*���Kn:�"�«j>[ε�	�YP$����H(�R� S*v��0IfL/춗]戂u�5�b��w��d��K�?	��p3(pZ&�TJA1�R��.�tE�R�Pt&~^��}t�z�gV5�� Y�➃�s� �noֺh�����DJp �]1�0�Tl�Ȭoǘ��g@�P�4a���23=���oٲE��=3΂��Ĭ�pɟ�/��2��ǋ���C���H<���:;P.�8��B��\B�t��$̋\v��$vnY�?���㚽��A�D(�K����<�ؓ&R�Yo(�̂�6ދ�^���ܸ.��Q�X�z5.�{6�[����O>���	�iui��T�!���̴L�z���7�X"����r�%�htdH{gz!�`~��Y]Knq=])��u�p�9��fҒ��yw��1�g2��ʫq�%#�	%q��aLNLH@��+X��lm6���kC�L��
�܆�DJ� ��峨W�ش���ć�ћ�^R8R�5;���s7�}��X�a����L���{?y��s%��}�����o�+�I.���Ԫn�?�X���,�p~�hB�7c v3yj��,���^����i���?|���Pg �G�E�҂��@w4 #��n�W]��F��)�seDZ~��U�J��<�p$V��#&(rL;�����jTG���1���&l0���0�>ST$얜'#A�������8�KDX�x����8�jU������n��=��MJ$~��?ro�D�Mi����������?������s�A��b��|��
P>v �j��n�KA��
�g��\�������z%��۾����~�gϿ��7���y����&��d(j���D ۷��/�G�VA:���'�씋���?�3����s�X��b-���<��I�u�k�ʒ�1O0j������Ȁ�%�9�P��#J<=I�^�e�s��Ο���	,Μ���G��`�B�2�P�k��R�A[�H2���E{�Ǧ��%pj���E�H7nٌ��!�ݰ}�Cx��G��܏l�s��$��:N�9+Vn�ܜy�<��o�FpblL�O��"�6P)T	���uË�?�Vۏ�t��l�u�nۅ�JS]�v �*!U:�,,A��VR���C��#/rh��GY�dq��0s����$	�b�B|�$�9��r:`�y��+���97.r(�/[ ����O~{�� s�N��R�"���_U�
��E�l3�0������@S�kw��!4VR���%iϺ���N�$� ���U���ʜ$��h�ٜLK
��6%���ؠ���[��b6����X؏D$����(+��(U*�6�|����
�*��]���i8���>��̼<0(=����ֵ��}=qaw����аEY�FGW���KL:�Az!�r��B��R�*;w����2tnL3Bk*<X�v5v��.�ӫ��,c$J���(�
:8Ox0* �T��11�c��ɷ��[����ЮT�C��E�,������ ���qr�,�9B���M卡>7p�j] Eȑr2>��U�a�Ĭ���ݝ"�ML��R/��vp`Ͷ3�i���њT�D��뙖[�&d$&��/[QG�I�Z�'H*Eժ�U��1�oV+�HF��I�Gϖ��<�=���IP07�N��E�²D���++��Qs���th2	c�Q7]
�m|-�!<�:%��h�ZHD��U����I��ڣ챗�"?��e�U��p��~�$�k
sU����Wa�谔�H��»��e�-���C�;/옄�q��[ց���*j)hq�ۺ�=�5�G�o0�`���e�E%h�I�<��r���-�,�e�űfw��Tg���20�&���s�b�����@�(��Q9QşpD������ʰ�$X�4u�Fy��/��܁���AP�	H��>��@�#KsP�Ѻ���`��.$+��Z���R�;r� �:(rf*n���1�.sS�ٰ�ş�P1���Ů�k�'_�,��h�|~�D����w����ѧ�E��X�}B�^y�Ed�V1�>gu�B!�Z�͛7j�P���s<��A=v�Sf^�BH$S*4P�	g�d���mD��� �&},:��fm�C�:11v���\��(	�M
f�#��g+q��=�^MD���p����ȐG뻯�G?����81�R��3�f>��	t$ztمY���X?܅�~�#����Wr�N����,��|�;ߓ��W��㑟�?���t���+���oG<��;�1��$�a��ܓ��T��vr���<yRs��/���*%���x������;zә�e*��b��5��V[�
�p���a�ӏ��1D�E��'ʗ�g���r>Oǂ��b��WJC��	�3y�g��)�@��f��_u#��-x|5|�Z���,'L�ZA���S,��	��CD(�¢T�@:cq4�~���ѱf5:7nBǎݘ-6p�/�GO���/�@���Nc�����?�S9�����Cc(y¨y��7�����m"��Ga�j���@����k�������_����s���O��}�կF:���@jEx���$��kcˆ~�x�ؾe=�="�ٚիq��kQ*��o}�'q�W��/��	��#��BްI}��y`?�Q��=��������omB��7{[�%���ڵ<fϝ���q���d�Ъ�ѮЬ���6s4�l.�̸xDuv%�aݨZ����Vadd[�n����A�a��c�LϤ��K/���lQ�c@S3�:�x0����X��}��>;�*1ߗ�Z�m:;:��w��=*�������v\���}-�� ��Uԩ8I��,�:t�5U.��M%"�bRA �K�wavG�Gaj�%7���2�2 1�e���.�u0��gd�\�����9��C��F� D<����} ��=���ɹ"��?;��tFcvd:gM��w�0�|�:7\����V�}��)S�3� �Ã=X7܅T�A��HPr�M��պ6��+�r������@;���>�ZmUg֮]�M�Q-���Gܚ�u&�HD"�c�rU�Īa�#��q���LLby�.�Nn��T���<�D�Ġ҃U�������Q/Z�r�B�*�Ц�x$��e��U��t&�!���T��z|^BŖ	ܵfMJ_�u���ۉ�k�d��@I�,�[�OgEl\Hg�>G�q3D��Y^@�NV�9/�&�֮����Hă(�2�V��û��mp��4&&�U�����,M~�F�GJ���5�ke���p }���09^\L��kadt5��V�ٳ�16v
�si��\��*/'�\��+Ф�q�@�&���nqK�v��Vfi�G��J#}��ӝ@�`J�,� �����#c�x��֚d8���̀�R+[�X���d��K"N�_*b\{I�/W�(��̽g�\�y.�t��s��f0`� QIQ�L�"eYT��lKZY��ڵ�U�]׭����]_�V����"� �"�$r � �L��=�s���}ޯ�]���u�0�����{��IV.� Zt�!�/����m�0�߇d<���%qo�� Gf$s%�5�!�9��sU	��`�h��/]D5ή�K�,�w ���B�	�t��
.���p8&��
ϝ�A�&Y$)�u74;�Zڳ�z*�'���$�B�T�U������J&���w��!�Ic��s���kU�4��p\��EATl��}54Ԓ~��(D$_�5dc7KC��Dr
��^eq��Vm� �����M���m��׎��ݡ��u�Fץq��4y���p�D����-��������N�b�͇\�ҁ�MdMKQd�B:����R������y���yRBd]43��QM�2j�h�L�K�v�n�W>�Gؿk*��2R������o��7Ԍ�-[�������\D�(b�~yyY
���hmk�s�� +�I��pv�m��hnk�u��ōX��)�0s��hW��9�K�*/H(����~ШȠ�3�s)�Z�5���P_�3o�@CH�[~N��������%9Ft���@t��d��J�-z�;\H��.�#M�l� �@:FO������ć6�J�e�[^Y���+��g?GߦA|��_q����ӟ��/_FOOFGF��"G��!24�����!9�`���uhQ��x==p�;�GF_o?X",�%���W��ˇ���A��NX�������ܷ��-H��a�d`�d蓋r&�X"xt�Pd��������byjH�Q�d��03�{�܋bW]��Ӆ�n��� w�MP�l�j�D���V��d$�Ǆ�h��kZ��5`�;�����k���k'1.��sG�������f*[4!�� E�Mkh����Κ����[$Փ���х�;w}�s���ߩ������_����g��������i�f�Sď&��:�ݵ���^�w�������~���w�S����$~��"MattFG�˂U�TпX�T�Yp��,~��5�'u�� *&]�#d�G�!k���G�fE�����*<N;����E�M^Cb}Fn���|0�bAZ.f%g�v.�pJ+�:8�*�MmF���𹐈Ep`�<����*_���d�+R�8t7^�4^}�(���$��O왬�N���L����_��y�P��"��b��H��C��v��y����}��ܴ��TN��Mf]&��w�6��ʄ`�E%�r��
�ܺC��K�K�y�<̹,L���?�k\��hK�Ŝ����NC ԏz�S��u�_Ra��E�BJ9����k��<��|�c�l�#����F,	��i���#*����)�\��k�U�:��ZCP�����R����*R`QOUk��}�h
:`5U�r�t�/K��F��*"_&��
�ׅtXX�brvs+a�x;�����,�`)�:]3����H ��TL���*�(05��+WǱN���E�Y��2E'��r��n̈́��.l���ce��l�ܼ�"}�Ȇ��L&u[�̩rNb�p&2E\�1�p�3�j�T,�$����@_o|n;�.+l��5�=!��R
�SX^Y���"l��b?g�;A`����"��.�N���ׁ��f�4Y�P���s��l�t��lX�Hcni�k��'��X_QDbJ��!�#�Ci��s����q:��s*�	���;<.y�t���X,#��E$3IA1ı��Z!������./JU6�7������h4f)��N�\W�\;F��u����I�i6]E\h]�L��e�������k��p����w;�U�ky�\$�O�l�"�em-�L�M}4i�����l.���¶���6�c�L�B�$����r8�l��\��dI� �[��x�:��D�A-��L��NWR��݆m�G�ب!�_���KcB��:�K��,���01yK(՚�0]gQ��eF9/�P����f^�e���&�Z������q�8� b�����(���r%�Kf�p��3R<���s765I�µ�Be������3��z�!�8��-*��:=�_�kNtwL�Q	�k��5� _��ªU)Z� ���3|�l��0]�5�-Sj���h�˿_�&�!P�*�&�L#��9_���/cq�PkC� ��]"�|=
E� [PT<3ѩB
�T��Ɨ?�	��5���gAR�����������݉w��طg�����B�H�����	�(��x�'&o�
�uyϤ}੧�mtb�8.^������`�犡V���2���
AJJ#C�<�C.��p��D��5f�r]�@@ht�2�	R�L29�,�ɍc8�m����yvzN��x��r,h�I��q��9]�N�Ϗ;����8�V���3�r�z��=��>���5�(����~����_�����~��-�F8y�8�]�&���V�K��$-��tʱ��:����+Q����4��y�&�V����x�G��ׅ\�6v/���{�5��1%[��5;:�n<z`���#�G>��Rf�DT�v��@��]��')ƚ:ݨ�눐��JC+QL%`���$���m�@�Wj��u��HA�*$u�%⏢���d-�۫��
��-ҊH%ͺZA�fC��V�7#���7����qu1��A�R���	f�j�t�h
��4vR-IC�K`�U�7��k�w����F������Ums��_<t��ߘ]~���G�����UD�7�xػs�{����p��	���!���~��H�3x��aww�`����j�Fm`�C�-N\Z�O_���u�4��-E�t�r�Ň²�n�n�X�M�_���e�(��82�%hU�?(��Ş���9���v�Ae�_
�m[�����n��s��1:,!,"c��2xE���k�y�K+R���!������0{kJ���lA
���u�9{KK��L�ŋ?�vz�'Dw�)�A^�F�*;�B�@��6<���زc���"(W���D*�d:]�6-p{=*�����j�`azs�7�d(�0�U�5FQ*!�Q��]��'+�ޱn��I�$:�bLꫢPʠ��N���_�,|MA�l�����A6Oh�<_�D�b3.شw��5_���5(�uשh�ת���dUZ�Z P�ǜ�_m�V��Vty���$����S���i=��=#F�$r%��n����:Ƨ�qk~U`F
"}^7��[�:�T�W�D~�M���$�,X0,:" �.anv/�!�(��IQC�I��*!y�j�.���ϋ��F465���#�M���%Q�C@�䄓���N�+:A���;�)���q�/E����; HW&�hGmM�����"6x��9���,���ǡ�Wo��ʵG�(U5�+�X�B����J�A,6]�h ॰��n�ϫ?����x�h��٥5,�EK��>d�öM�(f�*!��2%��o�uu �w��q
���Te(W���5@����łJ��5L�ܢQʊ;����G8�ĩ�13�����	�E��k�ڢ�&i�ⴛ��s`�mho�I�`����c���ِ���(U��hrz�K�hl���n�f�.q�1�Y��0 ���Ui�6�LL��9�� ��{�M�L�����48-%�����nR�r%�El$2X^	cyuUh��m-�hnF{[ҩ(ʥ�V��VKR�1f1��G��%ss��2��� �6|7:�;��9pkfW��#��U�]PR�x���8�&i�|^�^�8�,ܺ���F�2d� �@���I�K�Dc9Ѿ��V�(�uhDM��'�h�f��S���]]VU(E|,����\]]�-�����$'R����[祖Se�Y�ܭ�k2�b�:�^�fq�g�A�"O~�_[Y\�b��M�6������A�
�`+��C�W��T4���f�m6�,LO� �秷�S~orr�*�I��� �3hi�M"]Ɓ�������n��,�b`n~���gq��ҩ<�����>�Q�ܱ����� A"��bA��լHB�uko���_8'HB{[���?Ǟ�� W*���'����旖eO%݋���\V&�%���[aC��㤄�E)��9���ڋtFB޸��1��e����|�8]v��,���Ӹv������� ������~��G���)P��XR�s���q|��C,Y�����O����x����ӏ�J��|�!��/��['����c�|Th�<�|����\�#���G���|�b㣄���̒�F��h4�\�x@���ۏ��V�%=z��o�T��a��Ό�RmN��S�    IDATp`t�n��a�V琎�I(%��B�l���ٗ�xq����a5�A�(�b�+D�ё�����:�<�;��b�j��I��VA�����jF*��T��[�3�X�¢I^l�Z���Z��0�1g#~u�*�?�6�e8�:�� 9͊*�ܬLV	B;뚅��ɢ52.���i-&#�w� 1@ο��'?p�7?�g�����.C�W���ݏ>�������	56����8�g����/��9���`;�x�!t6�q��e�&}����߃�,ί��������%��`����f�8�׀�c	|�'gq}.���Rjz����SX��O��%����8et"^��3o`��E���0�J6Ji/�#��ڬ���l��|*�]_*�7���~[�$���^l^�GĠ�$�f;���5+&�o���M�OL
��C�����4�XD*��Qd@�K+��r�*W�~��l 6K�k����)���rE��V���odĊt�����C�l��U�R����R6���Ħ��p���ag��"�:�b�I������@�!�Q��\��X)�&�J�!�c-�8��D�k�Y�s�Ć����ub�B�@��W���-��V�U��f�py����w�e4dR�E��)�A�(7�Z��b�QNN�X�ӷ:'Wg8�%�M���2�6C%@��Kh�Y�us:��w�����Y�s�)Q6D�߆BU���"t��2�9=�+7&N�����Zk3W��@o{36�7J��W7��3��$�!E;AҢ���6������ylD�H�J�X�"�+?��TN;
����GK�*ނ^��A9E[Y]��{(�$�cޣ��inl'"����L)(������I���<�'��ʖ��6�T�z�,���55H�N�EK�	;-��+��Ԡ8��G���'�q��%,.��������f��alD9����pІ�ǎ�� �[p�+ph%x�:<䱓���"�6������9DY�(�� ����>5�K�:,pZ5i�N�m��c�Ù��3OC�!R=T�u1[�57&RR�YZ�~0�
���߬��co��ۗo�l��y����2:�cK*���
���
vl݌�-�B�`���9�orj�c�KowXa�PC �EJ���ǟ�^Z+r�&#�p����u��ee�Ir��h&���I�;�
�.7z����
����j��1��O�4R��sBis�XX.��Ĕ8ٰ���E{s�>3�$���]eh �.�,l � **T��X�t^�_R���m�����X�D��"Kcf1��5��X��*��7bSo+l�
6|.�|Nq%�,/�e��*y�TB4[@�PBQ����vc��IA��=�ZIZ��zD��'݂�Z�r��:��6� ����'Տ��@)y�O��o��p� ��i��YHmq5��]Ì:eH�ȚK��8����y��_��֖We���P���)��*�Z���o���J
3)�)������ݎ�g�`qv�MV�:���NL����X�>�X@5�Bvc�߅/��a��-R��-f�FV���~ׯ���-a����G� C[zn�;B�=�J����>'��0���d~��y8\n|�����HAx��9|���%7����b��E��`4ABU3H��7�M��pe^R�H�85@a3Ž��)������֓�n���L�:u
�ؽ{������C�&�zx������f��7��������Y+%���Gw#>���ç�+E+�F,.����5�_��w=�(�����%������k_Gs�T�z�Gr���IZ�ִv.��9�417oL���e��A�n��ߍ��s��~�7�����m��3����;�����S6�|l�dDr*Xs@B*��j������:�L��%�qI+.�(�H�-	
Zo�����f����	❤�za,~�Y�/Y)�0Lf
�a�1�Ps��G�+�ք�Q�H�t�z�Ѹ� f�v���%�~ueW�\y��@҂h^@ڠF�؆	�!�)Ww.�v��M߷��/��ǿ�ށ.L���jCP�V���_�ѯ��?�-�yx |��ؽm ��v���w�򮵥�:�{�����5>.�������x��ް����B����V	�
^w���ۀ�72�������$to��F�0�g��YmR��6R���o ��l�X�õs�����B�[JJ;P��7�I�;�2de�%�"�%}AQX@���Ǉ�|?>����S1��1�-�p:��K�e���!���xSK"�C|����SBUU�~�%$�9�I����5'������:u�/\��僦{O(䪀#������F��G��LN�iU�e�E^w�aw9�&�'�����Ɍ�,�-"��"���Ysb,�Pm��M���ŧ���$��
s�G_��i
7�*<P��*^�ɳ�i��`�=�{�|����ani^uN,I��] 29N��Y�"H''�=:)�h�X��u'?�~���+�Z�M�ӕ�������9��� ���1�Ӊf�6���S���Q�M�B46�ZJ��	\��)t*��'�3���8�c���2p�x,�bٙʗd�0s�l���^��7�U;|�f8t�Xyr��܃"h��.47z��K}��6�@��ۂ�~-ȥK�D����1@cS>��f���a�+�v���	�Ss�z})X�~:�K�	�k�.��g��M�2 ��"�̋K�ةga$y��n�B4��������m��z�f	�ǩ	Q���ƀ���ft��ఔ��m�%�T�1�ű�a���W/�����N������j!�q�D���R\t�H*9��
؈ƐHa�t�%A��:v:�Bw�2LV3Lv)����Y��t��6��~�i!�ϥ٨�?��`O'6�ke�v`ۖ>�mBn'I��-�J#�P^It�r�D��D��&eڹu� ZZ�V��*"@7��xO�_K��L�:p��U�<s�}��-ފ�Z1��8�6���W+�Z*���h��pe즈����&�9�GW�nU:�5>bkȂ��rR㤼�u���|	��-~�&�1��nf�H�gb�2.]�� �h6Q�n����n�1��@K�.M$J(��h��i�Ն2��U �7�64	:q�2W���U��U���0׭�F+�2%�"����&�������=�9��~��<��/���|Φ��_r	ja�B�ʬ�TO"����.v�^G��ʽKi��+�I��Ƭ�L*{�!���r�ҰH@��QhʪZ3KC^]Ew�BΝ8�%fq��L"�����7dz�h�5'*r�9���!Ż�ߏ?��Ǳg�4�l��kx��g1qu^��� ������%ҠB�h�(/�oJ�&�oU�Kr���>5uK��V������������^x�~�U����~@h�Z���8N�>K5��i�*֬���sq{҄v�	?���"Q�+_����Ōp$��'N�P�'��7l��\LI b-��>�֨~��P�<u��&���LD�)S�����<�?x�aqv$��<���<��_���O
}���?ڻ�P��J�4�BSs��]�8X�],�6A��:�)s�8���\���\8��%�@A&�+�x�
����c��4������l���VX2I���QI�`6
�z��iQ����`s:�`��*Ӽ�a$�ð��I�[,�]�����c��pf"̄Z�3C9Rcx�ȽSӬ���H�j�yIa^6P.����v�j׋K�Y�ح��XsZ�Ь(5��y�A8w��~t�,�.D�59�#���@�C �5<����V�CZEH��D�����4��WR����3��۟|�W�}����Ԇ���/�����G���lx����A%���~�^~�e8t/�/�Z�����C8r����:>���8x`/�\�N\��"�!���S�T��B��w#m.�g��9�k�x����³1���S��PM6=6�ukZ%;�X]����U��+(&�Q�FᲒs�D��P�X*ʐ���<�Z�`�gϛ�X�b#����>����W�����L:)�}^��d�SS��$3)8��<p�����i׮8p��hm��S=ͮ6^��/��I"$�N.�=xz�z��7����_A<C/p;L� �+���ك��$��pZC��*�U�.Z���!�06q�ষ:��TxH��BF�x���f�wGT��*�Hl}TP���G˯��������e�wy&��	C���~�#�zt�/͋�!���dZ���l��8�:�jx�(?��QRة	�F�*1�|�W\křp	%��LB�k��,E��#�����$�N�����-:$�,��qk�����&�ځlM�:���v�ʉ��$���d��2-H�N5~��7�ڱ3�Z��І�� l˱�*����5:����2�S��Ť�㚬X��b-���r��8������Z�s������3������2�:�X�[ZC"U�f�"�50��.<tIc6JH���wZ��{����A�.6���j�N���"���5Z��{�6����ŉ�0qkmD=��b�(�a1���Ղ�C�z̰kU8��5�
%�aa���z2��/t!�k�Q�b�2	��vw`���|��U1�7w.�]��a���.^C*Y���|�C�6����%�ښŐA �T�Aa:V"I��t]tF�	��UF�eY��\XD4�⾔���f���v�b��W�O/u�r�8��<n��#�t�9�� �/N��g�J�m�0v��u��o-��_�p�W�;"	�.N���q0^���DcK��~{��zBpZIǣ�M-��jC���d�`9�����!(�ȶa�t�%䂩��('�<��D��Ŗ	[�"� �d��������:��)E>��6'�-����j�F��S�cz.M�8��[�`��[�W��B�G�F䋳r�YP�¸JՒ	E��biÂ��(~��Y��SB�"�kG<��|*#bP
L����(��I-E�����۩��uu-�Lj�=;*A��+���=�S}@��U4(5dS�bc����\���x��P��*I����,LcqAHR�z�z�	�';CBk��|"���z[��[p��c��uK���LP6�|=��m��hҩ�F�4h&n�%��C���<�];7IA�.������K�t�������A�B�Z�4��E���@,�y~"����-C�XX����cضm��G,��4Ν����G�C�9	G֑���]��	����Fd�D]H<��<Ɋ0kJ;R�J�@'����k�b���?�m���[�Ù3g���Ol
��ء����v����#��SqU�Ĳ8ya����+�,�&���F	�!;>�����O�K�*N�٠q�|��W���/�#MO��:d����4Ї��n9_#�ƨ �kvuU�33��(4���=�]�����	��}ۆTPX�Yh�b��;՜�[ǳ��>ν�&lv���ž�>��,H�,���V�kt�TP6���n�ƒf*��i�	�s�*��Pցp8)�|��a73�E!�l���Ux��gn757J�������P�Lc>�uQ��>4ː��.5DꙥSfl�������u�_:��z%"ž �N/r�	E6��!����ƺLC�(�L����ZՊtx9}�涿����懶ne��~��7��w~��ߜ<��7?������	�L������,*U�>54|���Ͻ�
~�ӟ��o ����:`�h4��@��7/�"�Uq�c��5Ͽ6�g��� \�M�h.��j"�5�h&����a�
�-pj%d�k���6�o��XF9�]RV9�O��$�A1������	�*	���#������~��x�?$ԆHtU�+�+�qMn*6�WEN8t�8Y����ohp3z{����!�iR@k������z�*�S7.�[��	Wo��V�Z�}�:�����a�f`@��a���ix
p"��d�#�ֆ��Y2�"�1�Nʤ��� Cv�kX��U���PbB1�j�ڒ���f�`61E��,�n�=ʵn�BBm���\�$�L�;�	��)�RA��m��?oȇ��yq��R�S+6C�r�aW]#@!h�iD�_5� 7���nt�..�=}�q��O^nE,B�VS���ؿ}��,ԯ��ۓ�"g��M.���[H��Ȗ����p8N��Jk��b�rqA.��)�:�V��,�;t�n̈^���Ic�t�(22�:؅ݣhkp���d�zd��tyE$9����sW��G��T8'.W��da��ڀ᭛��݌��������#Ҵ���E��=��D�3��^^���F��A*��=�?Z�����l��ldo/!����Yi�x\�̸:���Gޒ:l��35�bM[N����x��uª���T+lv/`�`n)�߾y�q�y�^U���%�h
�9�Ek�)FM>�iQH���n٤!g�JX�D165�����:����o˩M0�AO_+��[����xE���1�f\��Ǎ�Y��6�J�����^�,ત��T�V6��REw;�`��~�����Keu��"�H��qz����vwv`S_v�lŦM~Anx��I����n�3V�~��L̮�br���fq��M�K���c��SvSE��4��UD2e\�1���q��d�1�C��#�M�m��M+éSԭ()�Ë|�
��s�x|k6�T�T�8��ͧ�-$H)'q<WԜD�9�u�2��X��� �it�}Vtu�0�݄�'�L�� ��� ������WQ�Hϳ�����uN�+j�t�K	.���L'�X_[����իrX\0Q�dxI�-��]R\��iy�u����x�����S�kw���<���sJ�P[�����ӄ��2���dH�eKڐ8�V�acCD�j�(��",#�D��s����籶�,A�Z�7�X:���`/�
#�Sʦ��XŽ;����ǱwǠ���*Kf����-�9�p�o���U����+�`=+��cJw�{8�}�"v�L&��E��}����j�#W����S����+��^J��͉q�U�}7Cػw�8��!�Â��<��ዛ7o�fu=��%�hmi���{�3��$���-���+�XZZ��褱��`":�]%�K�
Ai��aF<c������K��P�#G�U6/aoA��~�>|�=�JK`nՙb�}�M�p���/�ɤf�1�~at���۔�B�YDFI�(�^Y���1�=+�����:"�7���Q�un
�2���,�<z'^}-&�1�C�!��ad�W�%�4�R9��0�*�v�;G���q:p.��$���5��wa�.�-�&����_�Bf.�y�(>�0Ѳ���h/>q��3(�ƺP}!��94�N� ��N�l
�J�Jۜ�x�(��з���^��N㯿�,T-��	���b�!3�_��܂�*���(3��(
�;�XK<�}�k{��?���T0/Կ|��ϼ��[�}�=�>����o��B��X�N/�P�2t�˹"�]����Y,���hᔵ��x��{�}����]g �ZLy�����~�L��]�~~I# �o&��t�H�ݟJ���&b���"M(��[{�$���d7�r�%�t��bwH�oHRi�'��ȌT6#c0��N�߳S�z�7�7�ӟ�#Y�J���]����!�"�y����Y� ��c�֌؋�#G$�X�.���ŀ_\h�,�8x��-�M���*����������~�#o���� C�d�c`h'��� ��V\�YD�bÖ�[~�sO2�P|Hzh�('#���$��Y���X�Y��U mHd�=Ey�+ꄺiH��� =���&`*#BM0��N��VT�"�
���HC�kJCMf����*�>I>e�B-m��3����ԂZۄ�ɪ�2�ޔ�P8���-�72i ��6S	[�[q`�ft6�`)P��.�M�f;9`baק���!���I�
��a�]    IDAT��T��V�asW�ݹ=�~8,��P�U��F��D����~�"�x�,���ymZM�X4\�>ԃ��F�\R��U}���M"m�쥛8r��oV75��"7�\�B�T���GGk=]����PpL_q�G01$�c6\����I����e/s�X��`GH��}�pjE���8��3�C�	���Åp2�sWn���+(t�hE�i��k$E<�Ex�:6�����d�Y���'��O����o����f�.���h�J[6�`��t6pZ`3�-̡��!��	��7�p��,G�0����f�o{ؗJ�)L���D__+�6w"�g�H�y�{ND�E�q�*�ߜ����铜	>���c&�1�$��"��PF�������F�v�;E�+�sGa�I�I�pkn��]����\�>�vwb��0Z�9���!}��	���=�T�6��.(nD%#���-�س}P]���S ^4�-�qe|�/�@4U�ߓi15`�:�B�æ�f�6���V��t	t:�'���.�ss+z���Me�](�����\�J�M-3�]��� �` �C,E+�,R�vܿg+�t ��D�*|$"4\�9���X�,�޹��M����̴��2i�!@B��&�������'N3�lFʐU�b�̉��T�=��s��u��kR�	�7	����,����瓺�s]? �TC!u�H6)C,`i��d_��`��4���[���n�����
�(�n�43�Ks�����t��aҋ��:hl$"��uu	b�]�#�4���>��Ǳ�ͽ��XY������k�%w4����(�|w ��p�Z_GE2��B���l�166&nDx��ڜ��Zd�9����oavv{���'?�ii:�9��G� �}��8~���d��G�8{�,�9"ַO?�����u��-�G_��/S6R##[�/}	{v�������`�B,vAPD[�3]�z<�!g���M���e���I�ꕣ0Ln��S*�F��ؿ�w�v	x�s�5�;��;�C�yU��M��ep��G�Z�&�T��ƺ���0�iBt��@j�8í�#�IciyS�3X]\��
t����^�$�@ �P���l��/��/ ���[o_A��@�MGvi�D��*��)8,(�6W�eh3�Hm��eC {��J*+��DT�$D �t�b6��*A���X�d��At�Tr
���h�L���ᦲQ'�tPi\�w����b�� CB���C��� E�a�`��%��kJ��D�i����������G�.�ח�a"��a���o�j�j��P��z�x�m����
Y�8lK����������;���^y�Ͻ�#��i}�����@UDO8�������Jt	�?=�=LN�I���WՄw�����B1��,v[<Q�[%�8m���o.�'ϟA�������r�!੪7V���@�*,�$�Ƥ!H,N���
E|�:�EĂ�BH]��5	�X,�JC��7�Ê�e����;�=��l�y�U�-�����Qn�L6[����ĲkeiY<99�{Gww��&����^:O��)����.'>����F��������?�`�Q�Q5���ҋ�{D[�0�֢H����`T��	*I�������"b9�UG6����,6QN��Dڕ��}���7k�I�4+3C2����Ȇ@6!aQ���0/|ޥq31�&>���	�{G�?����L��#S��gY�&vѴ�#�Qi ���
����!���OP����:�~Gl��'�v��Uib��T���ׂ�;�r+��T3IfXuˑ������e���,��(�ch��,g1�݄������Z��.if̯$p��$N_��7B��/ݜ��bd��Ў�z��H����X\M���k8ui��_�LXY��Mr)A�3�~6��a�� B�TT�A���͋\фT8v��\�@��{T���!Hn���cþ��ؿ}nk	f#���%b9���AD��
�l��z'߾*(����ۈ�A'$L�&�g�V��lK��U�e_iG�lťks8}aL�74Zh9k���Fk���?�[�t� �A�P�*��`�9���i�tE���v8m>h�B�؅3K��x"����`P������%ߟ��B8a�ͳqkv��$,E<�q��C�/��䓲�*���2�m7a��#[���Hqj���,Xل�-��(���1�=��4]�&C��ؾ} ��_���
"fs�l����I���S��i�ɰ�
\��:��D�ژ�C��};EoU-ӫ��V�:�����g� _քf��xUs�I	:�Fb�H���{l2�+�2>'֥�d�\��زeɍ���D�.�E�[����	��\�9����X<�$�+0U3�=҇w�݆޶�&�n�))�9�+TNqi|�/�#B�*��/$Ǘ�"6p\ɹ�^U��V��*v�|�B��ͽ������R/��ڑ�'�u���̀4Luה'X��6��hV�������8eV����I����&�m��;��@B��ѱr(�@:ZB��	�Y� ��:t�&ǁ7�$�|�&��Ne���"�)>�N�	��[hphx���}�~�B�
����̹sغy#[E�����ZO&���A�b�(��:��ɤ�D2���E�vب|�������-�-�СC"^���z��/_����Ͽ����K���O}�����mH!Oz��=��^ý��+T$~0����C��(��<v�w������p`�>����,aiaQ��Ĥ�FG�j�Rr­���c�'&�L���D8|�"~���Z�(Rɸ���z����x���R��,��h/�r'N�D{{��Al߶��ZH�L�����+/��+b&1�u��މ��.�|�80���\�(��ff�<?�D8,�y6S��5����l�"��N��yud�x�b7n��ϣ��L�W�r�p����@�sq����Nd7��X#��*�9[D9EK�b�"�,C"~��1���B�j����=�t5݂��F���+{(k�P���Z���Er[�Z�^g�V䰎�*
�H��GQN�H�1�V6�;^٪#F�]g#\���e�Ø1l����א��Prd:H��4p4�͢���U%��(g���&���������o?��C���|��S���W������ں[w�܎���V�+�.�"�&�_�W3.ܸ��(�M���x��*��;:�v���n��+��� @��q�ˇdՄ�^�/_~�f['4�/�q	���yr����f� �2A�
H�Mcy�f�/#�>0w���k�4�Z��+�N&u�7K����2����ۆ���"Vzss��YܽwC�9>.�Ȏ�jqJ%���♓�NkO�|�af���Id��W.����*���$� �{{��jD'#��Qc�,I�V8�>���x�����ah>�B�:��bp���E$�E�q��Қ��4-��������s���H`zl�E%�Sr��8u�Ee�l�9�.�S�$.\8�a�ؔ�J�'�eH����U�ze�?������������'f��F�H�������zC@�`�!P�r�7 bz�����SmڂJ�8���L	�IY��<k5���f��Ak�	�]q��U���qƁ��"��uc��Q��ՃB����#ڠD�vs�;!h�Q �O[�n���"N�����e�,*E������h����t��	g��i6?E:�)
�ba%�k7�pki��]�,6�意��9�Lw���ɋ{vmFw�F.�Y�>X��r±"�^���c���F�@��T� ��c.c�`7��=
�����߭����Y�������q-�����6>�B�b�h,=���f�¯��j���1`C�G�/Is�����.�M���fA�\��e�H��	ފ�6l�*\6M<�I�sy��Z�k�Q�v�,��@�:�����6C/^e��G!Eow�nߊ��6iN� 3P���+�Y
�l�
B��Mx��AP��P�W~M�qR�.D�8�M�VŦ�fܻwTِ�+��� 1���0�&�'�t�O��AI ��@��-C����ǜ�����Ya�=(�-�X�o�<�\�.�G3a��f�aTs�x�`�A$c��u��@%3��p��k0@6;|^/��ҋt9��}��6���� �0���x��+8uaL�S���3\.7Z[PHe}Ld�(W
��jǁ�{���*V��Dc7�q�Ҹ؏����f���)�hp���waǖ^UT��Z���X�&������^����O�	&���F��Ų#�H��9%��p�Ά��hXf�e��Ÿ#���u���~���������X-��6�o�"(�*��մ
��c�sU%�������� /�|��2�b�*T��2O"�t�
,:���0rYh�B��=.�N�:>�m�z�d�\���!KAj*)ÜL6/\{� ��G�����'��][�� V��Ϝ�񓧱{�N�O�%{���C��������%`n~^����ߝ[\M�Sx{v푠���*^=�~����^��҄O��"�}�7���](*�'_�{y/���]���{���p��a)�yNZZZ��3�H�ꍛc�ɏ�����@�ğ�����\lɗ�ŝ�C����^�|Hvy��pe�Ia1�u�c%U�/��sGN��n4���4�~~������dkkzyϽ��_|����#=���EK63�X�f�����_;�x2�` ��"z��4(Z���.�+�lf16a�a,�*s �*՜)�C��P��-hkhA��D5�-��¹K�?�64�1e3p2�/����5���m�1e�E>G2�!�&ASY�2J�F���\����&����MS�T��5 S-��󠥳]���I��ӝ�3��"m8�����F������K�_��h+O&Y3���ќ"��6�� ��Mh��\#������C�c.�C�f|��#���Ͱ�^����z+�(�'"��#}��<�s����������[y�����P-gd�a1IN`WV����u/Vc	l$�By��r�����ڌ��Vl��@�Gx� ��<:MM�.D���ǯ��×-x`�Z`��n7u"E�\��p8Lh�2:���4s��0�@1��6�)�����+n�lv�ȝ�E}.�,悒J���P?z���Z��;/0#�ޞ�nI���?�p��1
)ٵ��b���Q��oD��������v�g'Z�1>~���hnlAg�KP&�����ݺK|����boC4Y~�"���3���M�ҹ�	u`������/�W$�C"[^9E��Q�]�Զ��	���#��:���"�ڀY6��N_,�*
ʍ�*n�/�(P|�ȁB1��QB^�ǩ�g�J�A
�Y曤!�ǘݻ��?�1�MN���)��(��@ؿ�-�C�������Vx񦾫ؿ3ySڎ�F}��,4 ѕ �ii8�e�ta� ��:\�?
��C���p����c�Hӝ���@:�,�D�~��x�v��Bw�_�	�)S'@��d����8{�nN����%lx�{FH�q��g6�%>�t�0'|j3+XK�!�&)�:�&sfW�nF���l��;7���MTH�To�@��N����_����h�0��
i�����Q��8��8ԐZ@��4ҙ�����d����(�ܘ��F.o�Ь≬y��P�z;[��ф�&7B~�Ej_�(V$R._����*L](L����;z�w�_lFy�r��c�N��X�څ��+�̕�876�X�+��ph� �A�B��f�qD7��Æc��<���*XZ�ҍI�-GP2�k��$�3]��ǸY9��T�4LP.�n�(�����[�r�JȺ�&T��Ao�ML^}�$�\��!�|o;08�*Bۀ���DFYZ�z-�.���061�������Q��yp��z��e
�"�4��|��Wq��5�"���ɱ�Ԅo[���^�����̈́â�KJ,a`f1����t�r�Q�`�Iʳ��ߌR5�|)����7�2�@-p��,ο}�\Y�W
�=l*E������v��]Є�S��jE&���Z4����qL.D��Z�\`�]�Ю��2��u��u7Q�KZ)����,��07/�_���wB��k��:�>�]m�����j�=�?Y�׬!�+���k�sR�b���"�BQR_h�-�i��fhMM�4H��Ƃ�(��k?�̭[2�ټe�;�TC�@8��D2)	�d�`���k0e6���_������B���ͷN�C�%,�]>���NY���F����c�H�0O� KKXXZT��\��By���'���m[}]X�ǡC��g?��؀S��/��q��|����l*�/|�x��GI�x�"�z�)l�:�cǎ�'?�	旄����~����������}\�zEb<�_����SO
�oea3���K�h	�j����2}Pī������P�F
������//�����i���!ې��j�����+��|�*���Q�^���Çq��u<���xp�A����hV��Jd�t'�>��gO��VW[;��~��n��0��bA����^���Z.#�-�4���0Hŧ�B�z�
�V],���
bӷ�~�&2��@4�B,*5���,��̡��	���SG1�B1�����gOf��RJN�"u��6�-(q�v鰺ݪ�-�%�(�ϣ������`��*�;���T�΁^� �~&�Bv���-�%��	ape�1�8AQ�@�"�[����-u	�ي�݊�߁|S��܇����t���|'.Oa&�D���@�6�f��q/`��Z�z��֪�Lt5�{�������_���!�Y������_9����U���+�Ų���ӁͰ0��N �wMfX\.YD)��koŖ�NV4:ut41|�S)�!�6Q���&�x��4�,Eo���H\+�F�B�S}FE�\Z�:*��\=���K����iX�?��;H��<|���u���y0�  "$� �"%K�hR�,˫��v�۽��=W���Y�뵵�h˲�`�E*�""g�`0���t��u���릱�������TM0��~��}�'��ȣR�A�3��(�	v����hvg��g�͂P��-ؽs;���#�3��%��k?����R�wtw���IFG�p9=F1�dׯ��������]2�(0��Ԇz���KF�!��\>	�al6ń��6S��1E���\�1�^�Ŀ��nN�J��B�l�Н��o�І���e1���@ʩ�`!Yg"9�HK㳈�,�M(�,lւl��bZ,�ذ����"�����H�[���	��)��a�+�˴٪I	(��Q	.$�؉g>�	��L�͊� hn
9�sL5DB}�T9�5��*e��x�[���M�Ws�m����� ȆM�OI��R��]=80H��Š�#'��1����y�N��$F���E�����L[���ף�����d�%~V�ŉD���\���RT�|��9�Un*��΃�;���݀��
��.�<p�&e9*&3�bx��U�.���T�<A+QҗY�F��sP�� ���j�bW_;�������	�l�ye֤[��m�xc�F'��X��X8�e�M[���6�-�źU��wy.�a�!D���6d�e$s�.m`=���S��f���<"�1�)���7d�B��ҼpaOf*�g0=��D�(��N�(=/Ԡ}�]����d=�6��[.j�d+�{1���Z�'Ocv-w]=T�"#�Y̛a5٥����}AB�,z^�ʇ��Ag{���ͯ�blj�k[����d�ߧ��cⶤjV�dEpωYɘ$����04�Mr	H-c��+L��iiZŊ�p
o�wK�Q��A0��8��������+"j6��eJ�X��F����)����P=A��I�v:�2h�p��~tw6�ZO�1���u�h�h��x�<�X� 3��Ϡ�k��n���    IDATFo���y��ͬ�)Hg-،�p����g�q�_x�tL��!��/#WLK�4�ͻ�;ѳmb�Μ���#���
��Rʕ��!���>�u�_�\I4KrV�" �9����u�F�(1���B�@�(��YK��y)�48������Y(D���1�ŵ��3��*^&���I��%6�����Iem�@���	����j���I�q��~�@�yH C@��&Re��� ?�K�IM%�r��uY{͜>�����5.�U�Fg�CJ&�D,,{Q�����4����4���2��Sh�a�[��`#]2á���o~���da��wN�����4Yy�CطsP�`iTĞ6#�ߠs$��O�D�ˆ��x<G"�#�&���ԇ���FN���ʞ���$�ߗ��e|�S���s���ߐ�ɧ^�$�����01>)+�����?{]�}�3��}��'��_|Q�ǆC`�������Z�Al��anj�tn��
\��U�B�u'4��}�I��:�k���-|��7�ʻ��U|��=Bq)�#���x����ǿ��&�y�=N�E��[�`qs�}�q��oC*
��-H�3:v�lE��Ib��Ǐ���6������2��0�u��Տ���B�L�;-���MFERA\
n[>5����O���%����G(]M��i���/B|���S(�ҰS�+����1��#��Ƥ�"3`x�p���
�B��SN���<�Z���i��. x	���dz2���ӊ\k�����z"-Bs�i�hh7M���j���d:-�i���
{���Of�V3N+�~�w��{aھ�^�+���scSȚ�0��`Ai��9݂����1�&��+��d8qx��������7M,�����_LMy���~�'g�f����2;;r�xA��'=c8���L8;^�1(���M(d�ho����@g;���p��\�]eqB�P�ۦb3U�{Wf��Ϯ`=e�2$(�I7�E܄�|r��58�
vq�>���k�GWyd�r���md��J�����OA0ř����s����g�N�u�a:<�Ӂt!�w���p%7�<5��ͭhhh��9�!�&+���Ȩ�ɻ<p`v���u���~��u?�ۘ�	��hٜxs����.F>��&��8�����x����k�`u3]���Ѕ�w܋m�ara�[q��n�T7lVC�hT�eTL%��t(&�	��-"�� D7a.�a�`V�(��m��+5�7Gx��*D�l����.��&S3�e
L�})�Y
�K(�!PM��?��?��43���f��@�>���E�l4V�����r��!�I1x���@���Do������IFIC&�����.��68�eT�� ;&�ɌQ�_���FEFN��ڄ�E���MA9�CGOk �-q,� �ת�P��`~-�K��1�F�bL�<.�k�6�1�ӌ�z'T+}�F�bw��eF�Q�-�\���\�V<�'��e��|At+���0�TF�931��,zZ���ӌ����i%�Hg��h(����V\���Vb)XL6���N�TH����߆F�CB�h-���5C*'y �o]Tt���D%�)"_�be=�KWF���	��'E&|�wbGOTGE삉�Db,�ű��o}6ʺ���)/Ͻ��G�v�(Y/��	�R��ݴ����W'��{�,�li�ٮ�� Q|�����.�4�[�L�#���*�6G��bh�\�c��>6��p6�q�ղ.��GWD�De��6q"�d��K��#��b��.��э�05�w��Ya����;?"�|��/�L:��5���h�[נ�H�U%���	[���Q�:%���#�1%Z�V
�m���{��+2���Y���k�@8Uƻ��F$��D�
���	��x�����"V�D���&�6$����UI�.Z��)QDS	�S�UL
KJ ^�L����f8��Wo@��$��au��IJC����[	��5��C;Q�J��$	�*���L�8<)ӮH��;��'�v��(UOr6����H���,E"A.�bE)��b�(E�L`oK�Mk��6���O)���S�k4��:���"�m-Ь���A��E0ς�v��S	)��Dt����l.W}βP0e��ײ4c�r�z|��o�KNk����361)_�z�ۤQb�'v�EL&
[>���z��gǑ�;�2��5�w���7�m�x�cOc��>��6;�I�ϭh�j��}�	�QD#�x܃A�� ��!�����w��7�|�hT�r_��o᳟���}��!-�/|w����2�eZ@0���o
���=��G�����6,<nԲ<��x�ÿ��ۍ�Ʀd6�8C�����0-�5x�&3Lv;��y|�>���E�Ã�s���+o��gG+��;Ĳ��CE�?u?���|
LF����ޭ�u���/1M�؉�j���1\8wׯ_���
t����&?q��P��-��ԣ���Q��'�b��A��8>����ni�$u��2W��L��STR9�Z���ΟG|j�H^���&�#�si|�_;�����DL�ي"	�G�I��=ё����(n��nCA]s#lM�@�G�ILR�ayz�Dݻw�]w���H�T40?�u6]��7]\AauӸoB8�~�L�.ag#T( ��Axj��!�a���bE�$m��������q��a2���8�w��D�k�
L%6����,�4jM@VS9K9;q���}�����3zc���>��������k��ڭ��s&#L"<2Rj��hV��kb�S��e��+�B�iV��{��]���"�d�4��P��3O\,�KC@Q�J�\�.�J|�瞣?jXܠ��ݮ�(2^����X�E97�q�&D�Q"�Œ��E�iw��eK,�uSs=:;�q���9~��R,������6<,����/X���x}��/���a�Ӷf�@d�TBsK#�]��p8,�Gc �fxS��8qP�V��r��(����$�D��?N�ngQ��/�|�EL̮CKW`u`����8���D�X�^+%	�2�2��.�TԄ۷������ڄ���՜�4���pť�b2&��B<�Y�#mM�R��Rj\����V)ƈ��BX��OXw��94��~��"T�Y���7q�TA��6%��?G�^uBPv�m��[�G-3��{�i��jn�R��J�T�bC@W��EcЉcw	���x�NjTΠ�8\�5>��K�S،��p.�6i�XPZl`9������Q���&�{m�U�].�KV�,*6"Y\�v7&�Y1!�q�5��z�7���
Ķ��p"W2c=��������� �fw�6'�n�l8!�n&%gt�Gw�{�ڤ����I����q��ȕ�ι��^��Z4��#��IF�2���A��7ë*0SP8=bG�U������v"ON<��y��ztbW��a}#
�נ�1Hl�`���)2�瓈���XX� �,��pI�Ŧ�뵉�ضF�꼒�@���~�t�ҭp���s�����$���
��p
����P]���h���(B� �Pȥ�K'd��mk���>٠nN�!�Z��jL�#8J(p�a2�G:{0��G��1U��v�w�;���3�&v�V�-.9��\���،�k��3Y�)o�p��B��t�H97�\M�*6+N_�z8.�L��N E��m�Ю>(
�FUI.V0���释�oL!���,��2J�,"�kh	9��Ç%�^&�"T�
�hFV�!�S���a�35�J�U�Jp;=�d9	*d��:�:���)v�`3���F��G�9��x�f*IC��َ� ؁���!,&xU����
.^����"re��q/���6�wp�fQD�ς/OJ��� ��[6R|��J��9�q�k�@MOR+�k~�RēҐ�!Y��y;��Fz�~V�Ԛ�?e-�m!����42��������ȟ�^4�G��ݧ��)`��̣M���WJ����'�fjnN�I���F3@*�b��!_{J���R81ԏ��q�&z>���7�g�����x쑇�P�C" �Ev�X� N�y�T�[&��C�_��1t�h�;֖�F<��#��c�1��w�F܂�<��}�w�>�����w����ٟ	�ǩ�=w�-����M|���{�w��������g�CGG^}��x���f�l��!b\N��^����A[Sr�	yR;�
E%��D���Ť���M흀�8��0���|��}mF�=b̑�/��ц��_���`a�h�{����K�������4tt�s,�Έ~� '�%-��w��/<��m=bLJ%�2�$��<�>;�ӗ�bzn��*v�u�3�x�;��ہ��5a5�Û���lhFС�Ò�!7?���'��[��PD��/�!���x�9�!}�a�'�'�E1�Fbe�Ur1\�&"&���}���ɤ��g�W��duM�`
�,�+(3G&Bѯ"NѲ8*��U8�d`�P=N�8]��y�:�Qt�� ;z>>ǢQ�@K6ln ���ld�\�dvN7��X,"C`�����:ǞX3���o]���	�狈��H�,J��,2�L��X�MF�!vߑ������������xC�_��㯝���͒+h���B7��I� A�[s���y��h�CA�B�*�&c�p���+�}-�mnB@��-T�nhm�310۝�$9�Z�_~�M\]G}�^iXd�a�,�bf(��2 ա���qi��3�RaiH���cwR,��p�l�;$ʼ��}�{����N%173�υ|�1<�����h��x��ױ�4��LNR��:����'�}�$F�]7�jZZea�C�D���8r����+H$�%vh����֌v�j�J�G�� 2!�Ƀ�LL�b+�BCk7z��`x"��������d�
���������+�|�depGg�۫��P�v�b���G�H��c��(]�͜A�EY�П i
��9 ;Om�œ@��,l%%��!ŖUX�V�
��CAC��3�;���~R�
זl:�h%ES���!�P���ZLP���x-�M(���>ݒ�I��*G��)����7^�%�f��p��9�-A:�~�'��I0��)|�h�dV�f�]Լ~��wc�8l%�u5�Cy�u~/�Ad�r����0��%���U����qذ��	C=�k�	'T�d��
(3}Ru!�W�����z���0��%V�F��r���H��11�@ո�J�,TKQ\�����~�Y��"x*(ea��qitF��k:MyP�g`�q���m��S�\��qv J�Z��'S c�E޵V6����VãS����# �0�w�]ی�R+eE���ƍ�3X^Kʤ�E���@c��]M����"���Q,��v���J�υ뷰��@*_���X�ՎR��1��`�i�¤XѨdPP�VB!��C1�Zĉh�X@���-vn��0k���RPh�&Tҙ�%3K(Ilko�m�uh�M�d����c��ZK[��ES9��.�����R�����ط�]��x���OB�����02���~yZ,~��z#m�jE��Į�64s���n� ���o6�ܚƹ+7���%N\�2�R�lm�!��ɇah�Kh�i#D�+t�p`t<��SX�$��	ba�ˉ>��NhI��xU�dsi)����&�Z�2ĬR*IR+�%�R��e�1�Y'>��!�49�(
5)lDs�^���s��ȗ�~Eq��i|-F;�/U֙�͈���N����o��C���TA��zJG����$���6<L�Th���NI�%F&#��n$��d���g���!Z�C��D�H�%������F�A[�~Wg�4460!�ڀP�$�F�T���&R�8Mgc,��ٴ����u��Hr��m��報7��������mB��x����3O���.��>{����	�N�B/�05=-��������:���EP,��퉈t� V�,�:ۛ���`�;T���ɛ���'���՗�(�⟽���/�B�Q��=����ocjbR4N�%t!���@Pd���cڃ���x�I'z��'pǞ=h�0;6��[c����X&-�A�I�45�d�����咯�P�� �n,n�/�~~a	�YC.�{L�$��|�G��c�¥�������?��WǱ��
5�H�&"PF��z1�;�8�/񷰧ǏD
����܂L�n��av3��H\�Xˢ�͏}��I�_<{
��⧈����܀{��CwE�b������k�9��5x���f��`�b��`^��N���4f�#��'�ͅ�H-@���AG1��l|�3�k��H��3O!�P��hW��̈́�^FN�_JQ���E�Mg;��G�68N�;{$�SDK[]�ׇt
��u�Ӏ�df�j?�u�8qw����@��q$<!�v�~z�
V�D4`#�GI�Ca�,M"H��2���+91H������+��o���]C���ɟ��{�h4��^�d���ĉ"W��33EX��RB!O���8�7�����@>�Svm�Ů�^�Ȑ�2� ��W���ؼ�o��[�xsCrt�[Dŵ"���T)����~Cp��[Hl�@c�V�!0��y�fp1Ul�	�⤣
�H��.�s�������������E]�!����~�㗑/dQ�� � [�L&+:���� /^��q�˩��$�D")j��:
:556�$�\D�P�F�����a���p��ゴ2����+8{�2|�-8������~�?��I�*��!4u�F��!�6��dSy�ilPU��BI���,�|Nڅ�N�a��5諳0�(<��R�eZ]�9��	�n R" #�dc����!/Q�Vl�*BN]�FǣA�����q�~<���pxT�//�S��4��X�0ʼ����J�������FvSx�O��ڄ����6���j�_���0L��.�CCh��a�+'+eC�N'f[�,��N`|v	�D6;��jp�D�g`5�"�mo����E�=��$E`p&E�JD���-�u������ց�V�DRR�1�6�ْ��2F'Wp��-$��m�$�0d\���MJ�i�vŠ>���f�{�۰��u.��w�`�� �T�y��<:���MY�d�@��ӊw�G{��� ��Py�S��/uA��Y!�ɰ8��l:�a+����
&g���{+�	R���9�F���jL�UK19�&������~�6���8Iᰉ����F:����qA�9f�6�K�$D�D'�Rt͒]u���~�,f�0� #%��mX-yL)��� uI�U3/�1���� �ƥ�%<Q��s���Q���`/��;Q�"G?)c<����h�	��v�dAha�6�F�s[����+$��R.�hd�dn��&q�9}�"�����C�PE�IZ
�ʒ�A�QU�������[�E!��FѸI6�|&�T2��?=�{�;��r�K7:R�ؔY1<��#Xڊ��&�j3�>x��I�Dx�������WdB��Qp�h�������ht-�������}t^��|Foj���ln�ob�֢�E����4U�Y��p!�ÄH8���MYc$���Ⓣ��S�3g)����r&�e@V���fQ��jr)�ǀ��'����}zdբ�F�	��܁��i��sJ$b���]]�g� 1A׋�x�Ō���ګS5r�(��')w��l��Kpi{�PT��ۼN$c��1,̪�����p����w⷟}w���A��/�Ͼ�q�;z�iF��193-4@������rQ��ghV�g�F�]55��}x�>:| �s�sb�������2Ƽ�'>�A���[��׾&������3�<#�13��k��8{����@�������^��$0��b��婧���}�r��~�n\���;U�8��ѭ&/TJ^?.�_�-��li��Ҏ��A�\K�ş��k�F�ѽ"*�DE���N�G=���q�hP%z,r    IDAT24צ��~�_�A���[Z�R/H[�lZ4!��]��>���{��ZJ����*�����5�.� 7a5�q��a|������k��#�L����G������@iq��X����&�`7)��6����V'�ȲPQL��x�"KKp�e��U,�ZIsn���[�p�S�fmWd����T�U+�P]n�%?�kr��V�,�Cm=����+E�2ӂ�����V�Kt�bj2Y�:<�~�S!/4:�7m��=b�bF�jA��B���h��!��o^��߿}7W�X����
3�Bk�@��؂�L5`J)�k��?���o~��W��h���~��^�Y�o�a��nǪ����U���Aie���F��,S��Fس���y���|�E���{���S6���̴cs��ZQ� ��Ƥ!�XοLƆ@lF͆�Q~A;M��ç�2!~��FC�	�� *tE��&�"M�tv�-�y���u�c+���c[o>��s�����5R���<^��Kk��܌B����M� ��y��{�ލ)�@�͆����X��'�w�^�n߸���7���K&���;��C�J�7�d,.�����d�r`p�1�r&��7q��,2,p��Zйc�,"���4�Q�l�+(������еfFưx���I(H�(P��bJ��e�O4���1�j�,�! �KA�b�b��2�Iڬ.�&� �n��8<b��9����T<�8�Lΰ4+��0J��,��o�2�O�	T�kH����ͷF�}Bp;��Y�|�Z���� �{w��=�������bC�d�����5�<ܞ����D����q��΍�ۊ�/z�\L�$=�h�re#��.�`|a.wP�h�Ә����u4��EL�~NY�L�r
.^���Ü��n�5(�m.�Ɔ@��P�x5W�E6v���ی��-2!h��ol2EH�4d�fl$��82���E�+�1"��9��]���%���av
�I�O����)wc���G���6;Q�Z�d��f�W0��%����{qh�Nt���Gg,���-��<��eR�hu�#T������kAO��&D��<��#cڕ-��\����'To6�[
%e�H
#���p95��mYoH� U��7�S|JN��J*+(�	�&���b#ː=&AKfVɠ���x�+�rPIÆ�4�݇z��J!c���]�;�q	����6�Q��`h�=���N�S�)�L����)�����[Z��i�A�>�BW[�dU��Y�f<���9ܚZ��V���U:�)EG������2�y螽��q:��`�m����Z�ijE�1�0QdN;\�5��@Wo�H�����8u����L�t�]����d�����3�"�֠����ݒM�����Q:_"S�T�+�T�`�q	:bآ�1��q�ɔ��t�!��t6RE�5!�^�Hv���-bm����$��j}���=��Z��f�?'������&0�ю��f7rj��l&%nr$�B��tZ>'�*�#�6���p�D+F��JYl�Im%}���F��	�)�Y#�xF�a1kx����ۿ���蒢2�/���+��������	�ǭ"��a=�eP�vI>&��|'^��H�tR�_"�}��@��z:q���{�	i~H?b�ط��[�'@�.��=��[�я~$I��|�s���� L��/�Ka<���x�t�N�>��#,`��<�����'����{�5+�~�.�:�R*��.�?K�";�I1��0�d�b���jES�LG�����s��*~8\~b�<��%|�ރ��'���:5M1�����^��g�#I����baZ��QD[��a����to�#됉��lN��� Y�T�t��A��1�Me\<w�t^����8<ЇG�A��Bdl��א��B%��5_�E�L�"�o�(}�І������H �����:z	n��QO���)Ф� �Dv�|Fv��W�
�WF�,�$UZ\��Y��
�M!��4H! Y"��ʀ49^uD�-
�ZIN+ٜ�f�r��Ow@���F�����`udt ��P���{��?t������?����Zi�,����D�d�1����*���=ۿ��?����Z5�?}��O���}j#��S�~Rmk���wɫ;+��E������ؘ(I1�E��{3S2Y�������X]�ՋQ����Νh��!"���
��ٌ7ޛ����$63*��>I*�!Q�+[�Y�O��knHC^��ȩ@|m��&�%�JJh ��2T���v�ai�G�.�Ć@�;R�ޱ�}�Y�n,�$��q��i�rC�f
2�'��ر��o�.�ꓓS�F⨫ɢǋ{hh�9�Â3g�㭷ޒ�Y��@K�O~�1l�ކ����el�#�/�[���&f��`pl$Q��̊�UO�:Ѿ}�d��M�&���+��UQ����]n�@,MLcs�ʛs0��E���H�uf�P|��ʎ,��"��11��V�6;�,F+f�L.Xl�?���p$��b	�RF�ѽ��ouM��]��*��y��1���%�¾TE�D�i����ܔ	��q�B�@&�(XUGp;�6t���^�qw[��wnÎ�:qB>c؏�aF0��)Mh��$ʠ�G�R����t�l��Hl��s�(x.��ؠ8�،��Oadr._ N�!�����h���4�-�)9(&M����9݅�x'���Ց)�s,
\$�R޿�w$��I�1��,���N`����w���A))*f�M���p��(��Z@��-
4UD�zd� ����
���czfN�A���G�]�]�*5D��d�Ε������6Sb��
�����v���MA���e\�X|���lp5�׹�s�{�;�2�TH�*�5���d�o��
C�&0�E��YQ*[��#ݑy,�t8�v)��|I�Ȧ2�ςR.'�i�U� &�,�����LDpǩ@��S
Aխ�u'97bJŝ� -�^L���mx�{P�t��e����U�.�g*�5+���T_:ښ$�E%��
f�y�%	�7��fq�ʰX��h���C�l�#�	���r`bnU�	+a�ͤY���)�$D�����u���C�򋑩���E(��q>֕�Jf$��0� e��J����n�DGG��-.o��L�.	N���$��,~��^���~1��� �D_gr�8L���ְL7e��KNx=��&�K�Ҷ$��[�Aw��.�x,)�)Z/�YF�/~YX�}M�*�RP�*M���p��T���W&�"�7����5����j� A����W?k���.�����Z+��K�}S�8��J���bX!Z�����pɒ&��M��
��'��Ϧ���L`��!Ј!/4Ҍ��z�����'�o=���!�O���3��᏾�Uq�ڽKlf���Pf�MI�T&+��Ԕ�X�)����#H�b�A� �*��u��=��C�eO%����/~�Ν����@��P��̌L>X�?t����a����N�<)�|����񜛛Õ+Wd�g0'�c��ă>�m]]p��ũI\<{+�3�|�I��n���Zb���M��ƚ���P<�}��������cЬ>X])賙-4�<����3O�M����f�������1~��I	6��]���~k�Z��V�e�%�Km���9�4��w�h����<�bZ(�A��{�BS}�Ъ�+�Cuh��ޢ��ㄿ\Ajv
�W�YX��"c]��j�@X9��"����]�>�E�VP�
C��O���&Db�e:D-!u>r��_�^��PrX��aR8�9��A����5��c7�"�4�P��~ev�jC�\@<���#Ќ��2��*�.�:\^����������.i��hn���~ J� �M��{o����ͪJ�&i��f�$�J�!�Y��������_�̯������m��Ͽ���x��/���qܱ�7.������azj&�P|�(}&�Γ�5�R���W��X>��G0?7���a�>ڳ�u��:U�|%h���*�<5���"�� `iEYq
�^K*�PkT�	^8-�4��N#�<�l�	��"o�QA>�p`m6��t�u������)<��	<�����B$� �1�R������<�@{{�L��,^�`����-\�tEf��&���I;t��~�ϟ7,�v���!�D���=w�=��F��aiaQD�MM-P=^(3�k��K�>tQw�3��RV����h����h4݊"}�eC�%��E*c�sy���-�ckn
���� J���3�&'Q�,��V��1J��Fl��Jż��|��=�t*[aW\PLv�M(��͆-�Z%tڅO}�shhm���*7ո���&I{[)��@m3����jeA��O�m����� �vn�j.C��4U����������V��Th!iA�l�}RZ��oV�:�ϗ��LA��6+��["�U3�|n�RȪ�8�X����Oalvv�GVA�ݱ]��e\����p���6��5a|~�/���rX]�3���� q�+�������	$I�3��S���F���!�F�[��)�L����K�42�L�,�� �z'�܋��(z��>#�)���8��� ��ߏ��>�U�o8��![/|�JNͯ�������C�����A�K�iW:1��+#ӈ���$ ��z'�����m��ʰrC�N�$��T7
��i��6���4�"p�9�D�ͩT"5��tyx*B�~���z�l��nA�"����0eچdQC�X�}n�)�Y�B=%:-�5�]6}�%�]+�ٰ^���Դ8LZ{��ăw��g��2łx� �����J�x���jhDoO�h.ZC>i�	��T'��4�bVqsb��\���.�)�Ю	�#-���lM˥�X�J�� =N�R6��~KC���kCW�>Ә3�Z}���z=����e�rE$�	�$R�P���^�_�����N�5׮�ĩ�W�/�P�Ԇ��E�wy� �c�n��#��K�`>�iA��t�ter1&��V\C��oj�D\��Q84��H%�K�c�A��dR����gI�g�,i�Db�\�ŧf1Z�*�&|�����6	�(cՑ�v��Rh\�մ�ꤏS,I�L���Oy�e�]�M9�,���c6Kc��$��K��g�N�h����Rƍ��X[[1�M"�l�t�&�%&��|kV�DO�&.-ӻ�~�����i%�Ű4>s�
~�+��X����nGGgv��#�pT���%l�����(#�B:����	0h�I���>�I4SP.f\�|���wp��e���yc�����>�s��.'�Լ�8a����v���k�J2�c��C���������jG2��ӧp����1����b(�J���x�u���'X�:����pk%�������YuIÕτ���_��OੇN�Z,���`jq���o��*R���rH1$�.�<g�sKe*A&��،r���EĽ� ���$d���.<�����'I�4vq�v��,��F�^YD�Պ�^Bx�
2�s�d��2g�6����X���t���8���"�����ȭm@���Z%���|^���CqA�%
������Z�P�Y�� c�� S�^�.�a���u)f�y�%���q�<2٭�5HfҒf�sA4>7��ꀛ�C�3#���>d��r�T_�����nt����ݸ4���~�oN A�9�f�,	�jeTh�O�m1g8饶�����w���������_�	�wϜ�����7��p����[Oݎ
S2�:%��F�,����)��f���*�W������=�k�/���5�vv���!��=n�0tB)��p'���h}u�C7�H���HS�D^#�����X*ii�ǯ!�<�tl�F�y�T�k0YHwQ`W��b�x��O[[S�p8*���1<��}�=�]��ٳ������"��o.����/�!�e���~����Y\�6,h������嬊�g$ҜE���
67V��hlb�P��������M.>���Ǧ�*����f��x��T��L�_]�w��l%rBI�IY�P�͛����V�P��@)�Ef3���[(E��n4�yf9de���g\���F��mٸ��v���O��B��?ʌ鶹���ì[�b �n7���n<��O��)�����o	�D�)_.JC��	��v̾���d
@�&�������Z�_���n�D����k�����B��:B���ok�iaqU���ņ�fE�#�)�sI"�A!jjg�5EA����"S�a�'<�2v�� �8甁��ő[X
�$�|�z�O���y�%��xQp�
�t6ܘZõ[��H���r��K�oI��J���b�.�!�R�Оmm�D�O.�B���V��ƍD�'16�&5��\*���G�C�-HǢ���T6���M\�>*��΁��j��c��e���㓦(�)�&6�Y\�5��5T�I�$��> �m,��j8���SH$)H-��e����у�Wu�i��:[q��$��M��y3�Q(6�.#���㢶`����W�u��{{o�`�(/1Z�!0ie�Ҫ/�� ��f4�l䰰���=����2=�y� B�/A�,IE(Oĕ���8v`@�Œ���&&�V8��Q4�Xي��w�`naIև��^������ȭg���{lJ����3�|uѭ���-�ދP���Hќ[�`xbK�a�4E�����P�(M��İ�.�CC;���m-�X ���I�L^G�Ӵl�2�
����u�A�2�e:�5��[����. �)p3���i*���\Gok O�{{w�����e�v�`R�Rk3��צ�E�*k'l�$g���]��<�w�g�,����	5���f�WD��5�&L�cٰC���5���.k�mf�C����I��-����L���ƅ�1>���� P6.�D��D��"[N�ʒ!n�f�����Y(r�Μ���<��r�t��v2٘YB�4r�au&��z^x�)��'���ES�O���?��W�Ʊ����ƾ�{�F����Uq����C4����u���E�=�H?��Ɔz=t��tw����<�^}�U�N����1�{���!'y<��ukQ��������d$횅<�26Y�M�˹���űc���`��vD�6��o�����M&$���&�R������|��9dR4��jF]� ��,�ۯ���zC�(��fSb�g�6|�+_��w��"<6fR s�Q|�{/���>R9j9-b	�����BOW'��L��[ayO4D��bU����=�T{eND˕v�o��>�;�R Y7U�4fcq��
f�\B����8����<�3���
�X����!�4�k���B{[����cH,-é��w:��5 �{���C1�5�,v��:��]�<q�z�8>���9he�ܗ��9�
J�"ss�2m��Hڝk��S����n��Kb�m&���`�<gZ�;y8��`�ƥ�e:�|'��Z�@0������}�)(݃�8����>��nLbK+#V(���I�+��Ć��R��E<�����8�������׋2��w����o~�
f�}�>��ك�S�����pcr?��{�69-"#3���^8aC��	�����N��s'q���܉����Gt��B��=�]bO�橛����HC�	���H@-��R�����Xa.�[��/M���0lGi�h��*A&D�dto���6�^�C����z7�����#��{�n���t��\�$c����pt�T^�tw�
-�7���{���%se+,)ih�{��%�N�LQ^[������2<."�n������v�i��[�s8s�:F�����J�~�^I{݊`qԡwp�4,��YUج�?�ÁU��F�.�@��l$�6�!�Da.G��rB�&VP�qR@n)on��-1N��0    IDATW}�A��9������&;�'J�
l�:�wl�{�d4pQw��86���������p�i3HZbě�.��Q��+�h �D�ǪkF���x;'���ZC��b����r#�2K��d��&%S�`zaE܆
NO� =6&aq4*�h҅TYd�~��@e����:�Vd�)�&gW$L.���`F1W�z��C܉��UiB	[G2�F��#��1����|�[Y��S�!�q�-�֌�fNY�� "df",i '@ؿE8L%�ؿ�C;:�%��t�,S���Z����֢L6�yW��hP�IC�o�Z..�$�����#���vw

H��eG��1��t-s�b�#�c���Els�:��gg/|~�ei���%\�>�~C�4�:;<��v?�E_YY���PkS�(�L/���W��J8��^�8�d�6��@�հ�"ݦ�яޮFt�7H��3�V�;`*���ʗ�x!�	�q��4,.G�ڒ͠�0،Z�����P%�.�O��&���L�J��E���pt�_�b��ٞb�p�h���p׮ݒ�Ng�}h�w��Ή��O��y�-X��Fz��\3�����2|v���A�
�ςH����G1<>�X� ����`D!L�}��
�t/�������e+��f���r#��,�Rv��̈ ��#)Ye8�N	��f�7����@�|�.����a	�S^��~y~!*VV
HF6��шG�>�����5x\4�6��j$�S��qyde�G(���Z'&�	��5r��TC��ɤ��,�Y,��QJ�Q�p�[�>��5q9��b��gm:p;0���4�:�kj�5��Ť�xG�-�@.5��hM��x�O���+i҈J<dCd�F�@�o�SDP*���I�cgN����l��1(��/ـs����*�__:F�Wŧ��0>����-$tԼ������ݿ���:��[p��c8q�=օ��5?����	��o���{6eZ1/�<Q�,mGu�A��5����8��Ȇd�>}Z>�[����ԟx]n���`"� A/�ך�_kv�<Gy
���4_�C8�/|����c�����?��_�*����S���!t���㢓�q���jj�A{�^ܘY�_��
�>se�UE��E6����~y�\��(�!�K݋�|�[�C�~��fQCKk>�O���E]�# P,�%��5Nɾ`p�@SC��}�-�������ׇ��f4Ndl-�c��i����r�`g:�hDjY����F��^��5���i"����!�Arn
��J��;�⎤�E��+��t�����e4�@���Z��O�b!�����6�	��sH��b���̭����TF�CE¯�R�U
ԏUPd�E����)^,�9q�yfsB`Z�����7�h^�!8v�F�cZ����E���e���Z&��d����#���4�_-�ȧ����{}��������_�EmG����������V����:���V�3�;{B��e:���I���Y\��Ս���Z�^�S1Q�?���8��^��֦f<x���4B^��<*D$-e9�,pN]���^����C����!��,"xB�:�E����&n����3o#�2	�� ��Q9�y �8��^����D[k3C!�4գ��G��¡C{DD4�0�x���w2?�!cL�0;v�X���đ�a/���,�
q��
n��D�!G��}�XtS��G:�siI�o�u����䩱Xf(��k����XZKb+Aj��f��$5i�����ӏH2+�+'"���S\�.d��t�b[K����@ۚ�j.H�EI"�5�TtUn".@��6�_:s��ǆ@�w�bL��܊��;`��s:�&�������yq�r4����觞��eǍ[�Pl*�����L���&f]☎(�!��M�p�\��V2��
�۹�5��f�����jb�Q�Ru�4׹$��|d�u3۰��p��hW�`����S�ÊT:+HBc��\
�t��-�nA�[Dk@>����������El�X4�r������ػ�]M����P͈gRиx[�X��06����5D"9��Ɔ,���i�*c�+%g����I-iy$�����ݞ4>���Q��Lg�<�b#�|6�E���`o3�W�+1�[���Fn��x�ǡ��YB��(LW�aX��@Ew7N[4�GF1?;���:��&��|�,�R��\�D&kԨ��k��Gv��QA!�����"���16�Y�'����Ī���&T"������*��	�at-�^�w��% 7�J��ur�s�M�3UԐ,�qk~c3��������<�E�={f��0�  ��"V5��$۲��qY��ز�z����NVrn~�fݛ����%��*�q/�U˲$��؉F�����^�z�o�������\K�9 f�������>�XNy�<]��UU�+G�j��ƺ���b�#h^qw�@6�hx����H��qu��Á�h[�4�ֱ��%`_:��8-�j���e�N?~N��8 �mau�'�0?� ��oQ25Y|&V�vqebs�Q��0՗֟��ZU�+f����R\.�1�ׁ�'G򐎙�K�VO&se9�9Xn���g�8=h:��-e��6��XO��^�4
���7,��Z&֊��\�<_�p�9:$.�Ԅy��r;6w�x��C`xZ���Pf^��|R*e
�Z���ޱ��t�{�I�!�1���NU��D��㿛�V$�����H����̈́�\������>|O,����X�s�M�$݇�r�z����ɜd�7�=���i,x�����=�GkSH�^:/r�ܟ
H&b@&I���
�X�F�:�*��]V���߉����a�'�2�"O<�,��/�;�V�܃���f�߇t*#V��s�H$�b@�����H#����b�X�e�x�o}��N��]f�����5��:�笀w�~誱4��n��6ߜ��۠��kED�Ik��y�	�����'1�/�F���Ǟ��¼�b<t�����9V��ft����q;�b_�)]sk;��}����o��x���(jttt"�ˈȷ�����r=�!`eP& 	���͇���p�Y)������g����7��,��׹��Tzz���<�T��(�wd7�W�i���_8�/}�2-�t��I�[+c/�r��y�ݰ�c�T-�VHWT@ �x�֫��P ����%�3i���#%��'���ȴ@��<Z�����҂�o�Fs36���۬�x`���KX����~�2l;I4���)�5T��)}��Z���J��Q�� ��M�M��9��M�>��M�~6&��6��>Ԛ��KG����w��^�xu������o`i'��WU�'V�E�A+U�(UU�1s��rz����O������0���׆��ϼ�����W���l�ۻ{�z��;p��w�#D��nn����Kx�Wg1����߰����䱛𶷽�'Fq��y47�q��M800(�˰� ��@�h��(~}q�,�e�O��%�5�Pr�u�6�X��.���^?��їPOn :��8v���yn��W�����EKs^��{�9�{�x
��~�|^x�y�}�<��a��1&����N��7�`(,�>��iJzo��3ʕ���L�䡠ƕ.q?X[ݐ��)���0*
�2I%�<v�P��.Ҷtjq��N`ayۉ<.�΢\�-�.�q,�9��7w�f�"ǿ��ȗ,� �Ak{n;Q��\6��97���*t-��44�O_���a�S<U�tLaS�1���]B40��`B���G8�	���$�Q�`�\�� ����pelR��8!�����H��MhD�\4F�\"fa+.!^mE5���W��(�#{S�g��9~f��m��^�����%�� �ӹq�l���?�d����FM#M��i�t�Z��_�u��Ў�{��!�m���)�&��x����u\_�v�&���&��D�8q` {��ඔ��6��b�C�⒆���2��-"������T�FV�&Xhv�����W�Y	M�i�����#��S��RPJz�1��zc�<{[�
�VE� G��Z��r:m �[䫯�������)$�8{{:1��=a�4�%4�AA���V���$"x8��:t��`���'c<S��j
�M
m�����$���-� *����Tkr���(�.#]Ա������X�J�fw�����")5� ��W�#�nG�BuN��7�Ǳ�0��L�� \�nE�X��m��_���k��G�=-s%�]<q�׬
/��Lɸ&Y��9e�Ih��ƽ㍷K�5QX�W��<�6iܘ[��VT����[$P/rK·�^����?�p��Y�[��-HS������hmk��D�-#͆���M΋n�y�]���p����:�~�t1�o���#8u|^��
�n�:jQ8� E�\���K�:��+�t�<�>���|�׸t}.�`��i��^R���X��JI�9y���KgPQJh$</�^3��L�^�:�WF�ETnp�@Ђ�1fO��IZV��W�be7�}�@a�7����녟��c�7�&��Z A�Y�H�(A����:>�B��4�����yfހ����JM��*���; ֤�ڴ'5ir�~I݀N1=��r	m-M"J�t��C�"�hwg�T6�Ns�M���@��\�2r�8�Z~�=���ɤ�9t�z�ٳ���"��MH���a��ǝg�H�)2�����҈e�9��c��4��>MN��`#��z-҅8��� ��T:��F�������(�L��I��2Ch6��� �a��4����'���&���3X]]�07��ׇ����N47�i�s!��}EZZ��aj~�����/���A��B1���Z�\x����g>��9�i�_�8��}�a���m����6���Ͼ��p�� ��.�CX�����U#@j.�t�v�_�!�f���bŹsW���_/�-���GO��SC�ni���F�ˎ`�WU��5��!�H�]-�cN��L�RA깞�Nx,:vQI%j��Yg-��{@@��X�ޫב&5��D�5��U�n<��J	��~��;e���mѱ;1��W�T!����\Ar�X�����cс��K� l�����Ks�
�
�S�n�TI�(��Z�(���w�ZN�;��%����0:/����!����4F�sW�V+�^L��>v�S���g~�����_��n�z&��&x_o'�Go[��vb�?BGU�y��-������!��`ycs�KȤ�hk�`��N�U�ae�w�5�'r00����_Y��lK%�u�$Y��:ڰz�al��2�t{�J�ޜ����ؘ��
�̉���אLa�Bn�>�Ve�����Ǜ�p
���x������ ��,ҶH�Ѕ2�"Ξ=/�E[����f���%�)v�E
�L�W�P��������s��cJ��6�V�nɦv���̗��+Xߊcbjk��6�X\��X�7{��Q8}-���ԎtcD_՜r���`s@�9�ÂB.�f�b�S�!(m��RM����������,@�fQ��B
㎩�hxY��!;�3��Цi�*t�`�>o�ע�&�&��}�Ň?� ��\�T\k���
�t1i4n���S�2֧�s^������n�&�'�LÆ�_�f@�p~g�E)Ď�Ş�&�]6T�(J�����v�=K�Hdi9HW{#D�"�ݰ��J�C���=�"���c��Q���|��x���6��p���ZEgK@������"5.�΂�RR�ay7���\�X��r��##]6��G�܀(8��W-����Fe_��=����ge���65��6P��2���^�Z����߃PRan�ž�6�_�(T*�n�191��5fl�u�-5D���#�fP�����ʼ�l�JȦw䙥�fu����(SK;�]�n*�L6�VDww�vC{[�Ҍꁝ��h+(5d�6l%˸:��˓�!����DGCTT��< lB%`3V+gE��е[�����
P�^I�E[?�H��kӸ��2qK�8��Y�&Q��E�t��@�q�X8x�7�X�ZM�Q���{1���a�Ņ��a+����9�^����p��4���xl�@���,J�2
�2��e����U�./"�A_/*�t:zխ�Y������9�l��,���#���S(zB��4n?1�7�>�N�ȜX�9],Bh�W�Zt�_�Jck;.c,�(f޿��Mp���B,V�K/_���)9Dm.����dY,viR'Q�Ġ׳��Λq|'�6.�h�`��2M8]JdK�\�F�F�<�2��]EDܻ�c�-��0��s�7p��4�m��k�J��c��g��e�G&�X%��ј�(����R��Q�6�?��攀A�����fC���ϯ���*NR���Ig�zM&��.._|�(l�M��9��'wQϧ���c��&�4�ɡ�W�NK�����>����6��ٓ�<���C���jj˴}_���/66�8[\Y��2�'�Ż��eym�aQ>���,���@� D-���˹�Hv�>).��~�d#��n�B���r�.����p� [5e+��E�@V#��Z+�P3@�(����6�pz������G��Iݹ|e_������kp���;���6���c����;��e�����}�a���!S(�v��N!�Ӊ�|�x��߉ps@���nLBN;Z��ȉ�E�ynGҀQS���kF�Zr��_�������ʵ1)ֹ�v:u������"Z	m�>;�ݵ&M4A�2A�_�Zxݻ:��'���bb�lv�I"u��!�m�&�A�"Y�J��Mg$՘���+{���@+�躵�%��ő���d�P���n�{>)���	Ҁt��/U�՚h^�^7JBu�>�7k������==�>
��c�[x��I����^���9P�(s��U���4��t�����ۏ�|�����VM��˳�������;i�E�6*��D^������#�+����Z̃�g�]�%ːd̩���tE��y� �e]��^�Z1��Ǔ�Oa|>���u�'Gk�=�+�="X4��UE9����/ �4�J�:3�6D�>r&��9h#"��M������ܧph����B����Ol>�$�)�"f����	���
8x�0N�|���L���RǾ}{���ӆ�v6qG {Î�ְ��+�F���*c��n�v��T�˫؎��-h����#�I�Ӎ�e�M���mA��Q�Z���HN���� �"/����Vo�*��-����l�Ϡ�D-�˨�a�P�o����VL�Z�H%��Q7Nk������M�o�
5B��C���P��anmDQ�����ӆ�ۏ��<A?F''��(v"��vc��c:��Eu�ǚ�!v��Ў�R�]��81(��OC��ڑ��$P�,��2�N.{��qpoZ��bZ��͎f ��bfq���	�����zV���R�Bv��ְ�m��@��6fD�X��p"_�19��_��RL|޹.9��l����nF��
'��Hȕ��nՂ�Tӫ��\��fV�)�h���{!�1����%���K���0�ۆc�a��^�[�����q��B��kbٹ�(�J]��e�59q�@?��D���i�g.���
&'�����B���'oFWG�L*�Ud���I�R��r1#�,�RjV�EsLd�_A<��(�R>)S��G�q��C��O�8�qʔK3�SG�jC�����y��:�D��/��P�sD�')6ጲ3��7��V?^w��K��Qc��i��V��ynEi��6�2�KT+',�6�i��y�a!�_< ��CV�d9�:������6�rdH&�*��X�H7���.2�w���p�ll�cn~Z��{���R(K�7m�3�2�����]���    IDATmB�����jŵK��^�n�"'�dUЫ�T��������x�-�s�W��I*G�U��el(���F'f���I��ʲ4o>y#���#������O#�,�v�WJ�-�%d�b�{�mG0��Ex���!�4`�|U v�9i��X��@wx�!�R&6�04�9�x��,�̉ ��Y��4���"� 4����{LD��͇i|�ߥ �TD���l~��Zy.�iKCXlNȁ�{
��r�8���6:�5���t��� �!������w�%��ڕK؍��n��dCP�e$k�Ω�P�y�Y��dP��nG|�=x��C__��N�~������T5�N�K�9Jf(d^�@�d���(Ia��d��GiH��/
h�Lq_u��*��HA=�X��<��DZL��2M��/H4MG��K��[���nX6�>p���SY1p�=�&Pc��ּ��y�Z�V��A5�x]2��{�x��@8Ԅ`�I�ǳs�x���cqm/Cr�;kh���~�x����)H�ʸ6:���oቧ����9B��G�X�[�}#��>���}����s�_���hdd��v"���19���zF�Xk(���x��w���W�L�?zO��E��9�S�W
Ջ�	�HW;��<\�-t��pW4X8)���������mB#�=cC���a���5$�W�<��(�`�v���D��"ת�B��@��$R��8goX��nC��S4�BQ 2�����xLjjd�4��)}�M����󒅿2`�V��=�!�Z�rU�E�p"�����#�Qh��X4�_����Ϗc7��bs!G�:m`I�yܘ��aC`���[����'����>�[�|�g{��_��ŝě���1-��j��ӊV�{�;1�ߏ�������D�Y.s�J�����F,���U�2t��#��΋�f�9ѝ�l���m���K�ߨ�ji��b��X�6�=����S�AGu�Cv�-EL��cP�]U��j:�f� �FÎpk�z:%�7�ؖ���������x�G������.=z�p�qp3&���h�$ǘylE㘙��B��⾁A�t�MH�bX^^D.��ͷ�"�0�6���)�#n��r�����>�N%�m���;N��j'����<����܁��v,,mblb�3�_ڀ��g��v�cm'%�x�P�D�+ڐe�IcP��-�V(ccf	s�^�P+%�٭�V�P�������g�*�Re���@>h�`����f�n'|�7MV$b	�<�� |��I���%�|n~^�Da�$=E!5��!�/sJ �3��PS|'E~�!0G����ޫ�-�D�j�uX�����n�i�5g���Eй�8k6�6��0��2q�R8�~��i��	�q��=�
�TnC�*�Nl�c3�x��E̬���ElJ�GgX
�}]ax�
L�6��dU�v�&	�W�汽C6�::4)[X
��Z�y�rC�I�T�RB��@O{��:��'���*A~l(�����0��0>'(y��hW�?:�+M�ӡڒ����&�S+�f�ߡS�D�a?���>4S�M�1��s���%�K��� 8C��F�7qe|NRk��Jꖒ���w�@[�)�������"L'А�/^���K�H�i��i&�tҫ��]��D��K�]�e=}�n9���Y0��,�kH�ʈ�s�_��ձ9l%
��-�D�`1LA<�2�@j�6�vHq��N'HWr�j��7��+���~7�>˰5�\��t��i7,�l���Ʌ,�.`jjRF�tu�n��&c<Q��iL-���psHh l��&titS��H�	򨃔��
�#�R�+��8�L
��8s��V��V���D(j�%�~3��׍�I�& ¦�����f�JE�fG2�����oLc'��4ךn:7�PS��കpx�G	���E��ҍ"K��o�R�<��k(Y�2!`�#����fI�nXx�{��	(�d�+�D�)�l
�יȼY��y�ŭ���ee{)Emc�mR�^�G�W���J
�FSi�G"��}Jօr12~?�5�m���yM�Ś�Թ:V+��(&�ǑL���Ag��G��J	:��Ւ8��:rP���$����|胿'�w�E�~�������%�(������/)���C�7�?�"�������sE�������NTR8iɼ�{l4mfC��3x��7�4���hU5aJ�&5�! ���/�j��72$�.��lP7����4�dC`��0;�[�^4Vl�4�Y*�D��\l��P,a#�Z�'��J����:�N|�#�?��b�AЈ�s�/�_��M<���p{<8q�A�nL�����/��7���O>��<��Ʈ�{=}�|�ӟ�������=�0&&&�ͧq���O>�_12t?�����o}�+Qq,$[í��.g��u�PG3ڬ54�3�p�`��0j�>/j��>&O����� ��+{ufc��0�tF#��֞@��l^%���݆���	U�6�s�r���,�l
;�Ԟ�$��1�4y]<��Ə{iT�z�	LЉR��4(i��eC A�bP���	��9*҆��}p�|��g����iL�&Pѽ��t�I���B`QQ�U�!R	��f�˷9�ɧ�����V5߽8��7��^�Z����M�NQ|sL�Hs�MG��B�ߋ��vq���+h�"�1ar�BMH�rXZ\�n���%�/� ju8\����1�p��
���������J�J<D��A$Sv�%N��#��߁�k���sO"�I���Y&
�u#%Gv�z�H�؝Q���@��n��>�[������]Sc�H�X�Q�J.�����/בL01>���5����;�o�>X���]	=��SBb����8��k7�H���ݐ<v��뫢O��w�[����M\�2���8��6q#�-�26���Mܘ^��N�@�����#�"Z-Rl�Ɏ�b�'�n��E8ɼ�b[s+X���VL��
�J�Fd� �F_�������a7��(��-����qRzȏ+����ڼZ��ΣN?d��.<s3������sc}s�ݴ|fA��;���e����@&Dj�U�]Ù��`4���@ ��?���l�4��)�:z�B88ЉވG8��V���o~�����݄��]å��YN��9qC!ǰX�o��Տ��fi�`�\v���Ai�$�{bn	Ϟ����� �llZ=mM8q`/��#8��X��`7`w���7��Wbx��$����E$�S-��Dv��4�,�*�,\�a?:���4)u�a�\��B���LO>	��k�\A�9Q\X)f�	�i��G�D���E,���n�qDc����'�B6KU��#��I3�Z�`��z�)�y)H�����M���Y)�-���W���h�]�8�mMAi�
��4#�jv�e=��5)L�t�;�G+�k��,��ͥP�{F.�^�mG�q����2}�����wMe��0�M�ܥq̮D��]p�!�S��8�<`���
�)N�x4��J�-�A\KF�����ێ�'Bs�#dD��?lt�kN}�%��m�I����L9[[�p��wc��KZ�<6��\�ݘxm��H��L�$=��+�XX��T#�����#6��t({�*Ŭ`����߆;����ఫ��\�#��#G�G����.\��	��NG�JG���t��	�Ҫ�P*�$tmfaۻ	.Z�e��烳�"*��:�i���0�6�$Es�l�X�/�O������V��؜�Ś]��p?`�b
~y̂�L�IGT���W]}���Wѿ�1�=Lj��b-S�BAM��2��kMj�9}�F�P9.B됴aUD�X"��i����1݅hy+�g#dޤxr͙{�4f�y�ei�Ѫ2���k��g���� �J���a%͌C!�+�<�lj���>�>����@gGg�=�������[1Y�<��PN>>;}�ϣ�&��7T���+Ey^)�e$׎�皲�pTM��L��F�rT����❮��ޱ ��V`��V�uI�j�t%gAǦ�ֹ���Uc��,��Q�J3FGU5���4M� �J�n(m'5�._Pi�i$��t�� ����Z��!x��g���~���%؝��u����=���B�^�?�~7�x�	|��_��R6���8���˿���0���/�����>��f��a�������W����!�@�\�>�������A/���x�&KF��n�F<4Q)fs{C�#�%b�e��ڂ��X�y�ז�\Z��iC�Z*�W������8�1�N�k0��j~�9#�BlЙ?�hЄ�W�#��	��M��H?���FѡE#kA�k��P6�V��ۅA�`��vt9	��l�]8;����M���b����ZP5�H �a/6�I���Ttu�ԑ�O=����5!��׍�<��{��د�>QӃVo EڼQtS+��[��ڊ�f	{��\�n|YP�hq뱛p�-7c'����G$����U��T�!�Q������V��</���#)�ұ�p%r�w,v8����~�]H,��쓿@tu
��3������H�z�w8��=ݰhl�lH��_~�s��ԭ��r�����˯�sA{W�x$�+�M��œ(x`�1uc7��UB�Mm�p���ر#�7��h?�0�]�.�5~"<��w�d����%"T�>t�{���L�����bl|�NOW旷���������2�ַ��=�=C�`�6��%Qk�2�<*L���8��^��@>G{C+�R;�kX��@-�K-�Z��S6��V�?9t�tZ��h�͑�]��-Ɔ��/O���Qm��y�#U����ێ�]�/</V7��y���;r���߀����Mᗊ����k�����(�Y�u&���Ex��(�5�]-������˶�,n<@se�܆�J���Wqybe�2KC�R�i�ǀ+�K�"�Y���$ٗ�,��I�U]Ǎ�U<aK�EI2�Zj�t�'���.�8Q�V�m�!�[VdJ���.^|�F'�asx_}�X��Ƃh��l1���ي�H3�ۚ�) բţ}��]�(]��?��EL-m#[�A��h��Z�¨gpdd��c�NY��\	kIܘY�v� �w�����8�pw˱�h	Zu�R� �//��&9դ�!�߈��+Ӹ4:+�Dr�lZ-!�8<��� �+|C�?Qu���"_�Å���dP'M7�!P4D�v+�$*EحUXk�me�rx?�8q�$������(kp|H��Ϗ���[�Ҭ�u�4�����P�aO)6���D�
��C�3��<5dQxlU?�_,p{ښ��(��ҝ�"I��ʘ��D`'�Ƶ�Q�|�Z�M�ݷ�C=]�K����ړ��l�yֹ�5L/l��$�J)@s���6�4�i��Ui>Ģ�T}C�e�ءh�<F�()',v���uDw��J������D^r�=>�ʖ��&a8Ծ�zĊ�����&v�)褫؝�w,����@%������!�dաiE�ҹ]v����rO�0�����L�H�`C�� �],֤�&�����M����4��NL����7�@5f�b
��I��T!�n�8�-�)L�[��I��\/.��:��Q��?e��o6��)2���5�����J�\�:�)+��鰢%B"��/����*<�І�h�!p2��-�4<�lT�%d�1��|������ކ��&�eaj�Kc���:&nL��16|$L+TS�mo�a28�e�����sr��{�}=��XR�I�cW�B�ٸol:vJ���5�����(?_5�j��h3MZcU�Kڤq&p�,�U5�}Z�Sc��!y�rOc�B@����dA���i�j�"V N�u	�$�A�>Ț����=����|��#0�-�g?����q�긤;H=A�5�������×��O�@/q��-����7���E|�k_S��l�����_`p`��?���}J�r���xum;w�#b�����Mm^�Ji��:$�F�\��t!w@&I�lJ�H�Zh�Nǝ\۫˨��� e���Uq253j�d��55�3^W��4q����=�F�RQ�:�9E����'j>%"��Qڨj�#\�8��	��n�Qa�
�����Ձ��~4��3�禗��i\Z^�B,�T����t��dt�f��iiOt4�ѥ��������G>�����/~�&|3_~f��_�֏��O�XCM�3���A*�����w�������W��6#�N~����r3�����򕋈nn��[O����*���ؗ>亠�u�钆��7���?�ո���|rh�����
ɃV�f)�)�����a���83�2�Ņ]X,E�ZI�Y�-S@jw�E�_*�%��}��.����uZeBp��E�n�<�p� �L��M��N�a6��p��(���`�4`��}����ؿP�l�/\�#�<"	%	����E:>>*���Ȱxs��74�w��]��f���1Vע��?�x�$��wX����Ģ�k�����ٱ��D��<u
���%��8%��l�jY�U$W6�6;�Rb(1��Թ�2�Pč�,&8�'�BgA��$�T!�\�,�fW^*�j� �)^cC�s�L<?旗��s3f3P%�&>�
��P/5��tܐ1��H��kx�e6�$l�O�k�y� 2�4�.�4tЉ��l��A��F�I�Pډ��:�勸1�&����E���p�t��b3tb_;F:�b#�i�$Hk��@��.m���l�V�!pU�\]���ώ��q�� �j�����t�1�ڎ��]���u�άBMg
�� �#�LU(����>t���n;��Y8݁B݊�DO�xI��d��C�dI�W3�i���'�N�H�I�K�6:���eѲ�Wh-:�����h�p����*5䎲�v�b����95/�ps�1<q3+QT,N9���M$�5��f�+�������y�,5�\�Ն�63+1L/mbq#�T���8�P<h1l��hrW�p��pZ��u�e���!�I~l��3��½�llϽt�O�uc���л�eb1��4�\�C6<��lT����Z�	�����]jz�B[�R"�R�F���E"�UD�el��������
���{��ގV�%gZ6iXe��*�G�t��\vqr�46+�m;tsх���*
���Ng����b�#�w��[nB_O@lS���=��R|�������z��)�l'�M��F�[�t��~���as�aw��f<��c�#]:*�3g�K��<�����80B5���b�g�*�\�#S�!��blnc3+�g�B�����#�HD,�/�8U�o�G���'� �����8�~������3E�f�n"Ȧ�P@��������6iD�qHM�UEI���B̀9Qc���L�M�	b��b�T��6�U��Ё��� ���t��J
�K/����:|?v��J��d��HgT*-�&��?�BS����~�=����]�^�4]�.]���
����Y����J��'��oUy�,5v�gΉ�餣��b���'I��(��s*�#��aeuKkt+ʡ�hE��t��� R�x�%�J\�j"��������)�kf��CuNYZӪ�SE��_�T�r	o@����&D9Ԫ����!���)6�k��i�������AW4 ����'�����.^E2��Ɠ�5Ҍ��y|����P�+_���|�n�;�/���q��!|�K_¿��6��)=y_�c��������1q��vڢ�V����ƙ#�WQ�X��N?��<R{i�L��Ep�,	�Lx��'i7���\n�=�0ܚ���ui6뜢p��^(�j��fJ:�F�����������I���׉�T�?� ��/�Pu@C��1�f��4l,�1(�B��Z g�z8���^Dat�a���G/\�������W��U�vN88��c���f�8iܕ,J���]'�|�ѿX㕆    IDAT���V5uǏ.�����g���)y��m(Y-�ۈ�%%?�^��Z~Álz�X����D���Gុ����+K˸�����$؇��<����T=�����[���~��Vw7O�x�s,Hq7�����GE	n��hqZ�4uӣ��:�vam��bo(�B��U8�DZ���Q.fqhd���qӁ!��yLN�!���L!�������'G-�.*��T������t� �����b5������g?}��կ$ ����-S 8@ǿ׮]���S����U��]xǻ~�]}x���pcf�`�ݏ����܋�����,�5�����'ʝtZB�(��9}e�x�*Z�l�0�kHml#�4���&jE�!`~CVh4�M��(�Ħa��͍O��PNJ%*�)?�+�Ft��+b���@���p���7������Ej��T\��h[�����%�!m�p��8��A�L�@н���~�^�5�ֈ�0B���#���_�?�V%�f�5���צ�x��_cv9
�p#��b�紆��r~�a{��oOA/زh(�bC�.U���Չ%̬f��KV��k���f�PVn=2�=s���P�L=�l�2BY�6��b�e�&�����æ�,�����=G���fw���h���R^l
Oi��ӓ���Zނf�
M�W���R�p�� <vH�͵H����^x�*��9��؈�j�bVɧ%���3�HS�pP>�V!u�ߋ�5qz`*3u��-`#����.*5�O{�ˀ�Z�,���49`��E�+;�`7[���2�O3�/SНFg���8)U��9�%qb:����~t���Պ(�7Ft�M/{&�����KX�eP�8��F���4t�j䨨S�dD<װ��T2f�ci��,e�u�����)���C&.���τz�X��*�$�Y����YL�O������N쉰P��Vd�f�EA�j`�̮��\�����
�w�H�JpR���O틙�M
F��fPͧ�����'�o�v�(�\��ܦ�+�f���UL/mIA*�Q9�Ȥ�cA2ʞ�JڌM��L.&��JwC�5h0QD)CG��y�=�0e��t|K�dyH}~Tk���u\����9q�bv�R�!�} (�2a;'��q2�v�3b�K���ߤ���5����|=���t�p7��r^i�̟e����6��q���#?\4h�� �,�ޤ�Q%Vf����)n;kWixh�)�V�ü:�1���cm���f��1�*��	�>����8�Z.�b:-|mK�*�!B���8��wߋ�ϛ�o_JE�qJ�US�*��L�kO��<Hh��P����W���'�'?'��j��Ns��3��rQ���R�MyՂ��(�~�9<��_c;���*wFN��h��k�Y1r�*��f� �#�$�: �e��J&�#J��ƃ,
[�3W-׃I��A}������&|���9a"�q�P�J�BA7�t�����!�P>4�8w�e|�1��"{O�Z���ui�~�wކO|�c21x衇��g#�����7���$G��������~]�7>[��~>�'��޽���W��Ǐ�~�&]�`�
�{:�޷�	LBڝ��+EĮ#d�Ò/�V$�a�M-�]�A�OѾ�%��1	$����B�x\�Qg�"\�oj�_�+�g��V�Z��2<L�v���2Ǆ� �	���Ȓ�� C�Y*l�${��↽*ݷd��u�;��R�ӭ��Bٰ"л��6��"�ׇ���_��O_���|i݁Dł����BɪK�	�#�MNK̆@�VQ%�]L��s��O��/>��oUC��K[��������܇�@+���퉬)g��t��%5��9�� �#���؁�����𝇿���9���o�]����i;��_cq0Ά�ŁsW�񝟞�����U��Ƀ'\ݐ	A]����O�^��V?v7�1;qk�㨥��������ZXD߬��m
�r؅����+���p Kk�x��XY]���D�[��˘��~�+X]��Pd�x�,=�Q�����D	�s��fp��9�'�h��>��X�@?y򸈏�6@~���n��4�tϽ�[X�<����t#����؊����>�مuqL9|�F�Sy$���p�K�kkHAme��K:��n��2�m��΢��!�T�q:���h�T����D*�8���R�����(7c�%}I�>>Pr��a![`�f}�o�{?��2�0'q����ϗ��/6f�Xc�ȵ h?��|�t^c��?��!S�g����p���O�HW�#䴢�Ń�Mhy% �16,.b�*�7�=?���<�͝(�X�1�Ԟ��I�����v<�Z^R �q�.D�z;�ù�70�D1��LJ9%|N]�GO�<�����">�tk`�U(հ��J͕�u$�5�K�,'G�.8BZ�QTO=��^]�.�vrma�P�X��ᔰ���D���3˘Y�#]Ԡ^u��ޗ3�Z����0��袡Id<��[;i\�6����%#C��_'hK�RNp�݂H��}=�ӥ2*YA���ށxU�R4�W�永�@"S�]��5����ky��r*y:;Zdr �Rp�*�Uo���x� ���p�°'��Ws�9���ΰ�N@W$((!7tRlt��L	�N�0|7W���s`�B�L���|v� k�X��:-�Pʧa��?���C�D��1���~�P�2ټh���QḼ`|f
��$::[q��C��B�n�VIK"��j�ՠ���f��__��/\DZ��~T�6�Dq�� B�ڐ��H��\^CC�Ê�8<�%�"m:s�����ƕ9��i�ZG��u_��l��U���h�7]�8��	��r"�L��as�a� [GG�o}�)�4b~�A�`B!/�gn�v��dY4$g/�a7WS9jq�<p��϶)��,�Mߜ*�}l� AĽ�@�����#�M�l"���6��@MT�*�Hi*����������	 �҂$� +�
�y�8S�����uռ�!P?�a����!�2d�'x+�ɮ���ͦ<㤔�x�Υ�.J�������?�t$��ӥ���߉�}�hk�K�@�=9�<ӕY�o>Ol�mB�20'W�PJd��x��S {�*ֈ6��HR��Z��D��^	�g�
�;����=�09Y ]��y,"y���_�lB î�f���w�w��V�v�&��T�g�M�q2��ƫqޑ���
��MGcm����4����Ib6S�%^� CNI������!4(^�n [.���x��"��I A�K�.�X(�ԩSx�����!��O~(@���Ɖ�O���CϞ^|��ÿ����w�)�p�uw�����>���9|�arz�\A�Hs��to���mV��L��4�Ztz&�Ӗ|Nr�+e�6���j��ކ��[ص:�6.�u(�3rVqz@	s.x�����RVV��	����f5%��$�f�ƎBB��Ui��tZA�5A&�R6�fSF�U�7j��T���%���	ks3����<4��˃+K[�����E����V_3
�U�u�K��=T�觨�e�q��v��s��G����?�[�|�����o}mv#q�'�{ $�,�t�kL��x:=�keAuY@��u��-G�7�?��c}mw��N�r���!:��NrS5i�_�Q��Vg�:�u��Xl���'c� �7\�vK�
�����q�\��bb�Զ$��,8�mxN��Hʩ8�~�gn;����N<4�xb3���*^������"l}m�|^OH��D*�d:���i:8�e3�hPPu�����+X_ߔ��)5##C8xhmA����Ii<����#�܆��y/_Gk�^���nkN|��O�W/\@Mw�gϠ4	8ϕ�+�Q���ؐU�8mJ��p;�}ri�U�$�7�>;�r**(�P��3k�lŝYPz6
�'/��pM�ł����#��(�R6p�,4�Ҵ�q���ɂ�3��w?p��WV��j��@��!��b�!��k��X�MC�j�������B��W��Xԑ/f�s[%Dlog3��=�tx�M@�����`']�j4���Mcqm��XA��ڑy�r����12؅&�Ulp��+�t�܌e��+c�^J���R	���X�ED�n������<<H�R|s�N�~rg��Y\^\��N�,���ȁ5�ቨ[��D��;�t�����C{��2�|j�y��Hayc�Ӌ�Y�F�b���*"D����8yx?�"!xi&������D���$m��*�u8�)���˹Z��a��`x��Mn�(��%����6vp}v�+Q��5XXR�I�F�"J)��铤^�׀æheb\�)AM��z�L`bz��怲Ŭq_S��]g\`��X�lǑ�>�%��Yy��=�h�0�:6���%��^���CRl�aP��Z��&E%��U�x��$3�ɮ����G�(�ZHȄ��B�n�L�R���Ņ��<^�>���9q���4�v����8��.+��,z6�Sh	5z��NIs~���y�22e�l���<Z�卜:Q|,.PE&ǔ��e�4���(.�:�sb7\�Cr2�K!�Ս�ՐÙf���M����<�ץ���}px��Mdd߭�֐��|W}�!��t����F��LZ��,��N��.���kS���B���?	�X�ˁ|A�)T��M34)C�w���?��Q�Wh�IR�&��`����q tN=���*�	T��B�mR�(�������-g�#N@�
�bE}i��`b62;%�B��w;���4b��vv�uy��g������t�).�4J�4G04\���I�/�U��-�����{���،��@]���8%�I�;�il
��C�Ah"|6%����2t�ө��Ԑ)���*�A������B�������#��M�����|��QW?KC(�(�8vt��ԃ���M��)�$�*i^Ho�{4�i��F���{5�2�Vnz԰�ɛo�#�'�'k�H�f�Jn]�(�t
K+�H%3X67������2R��ؚ��/뉍��䤸%B{W�����5\}��ͧ��ۍ�G��#Ҏh4�������fg�J�1��z���M���mkkׯ#:=�*S���3Z���nB�	�-�X`��+��А���"vE���J�PR#)�e%����<!��gE96��ƓBa	��������7Y$܏9!P?Z�$%Y�����I��S���Uؐqbn�wO�FB�`lu�����-"g� ���	�d� ]��hs��� �h�x�{+!��45�}�:�sw�z����O�V5��ԯ���?�[۹ʭVw�K%�L����:��e졂�*r�݆!�z1�3��ě�p^|�E�<p {��"�P�rN�$؜t�HƎWƢx��g1���v8|-���K�&`"��T�.����||��W�]��q8�T���0S�x:#�͆�Ca���7�o}�.��.n�N���+p{t��KwLG!���N/�B-�y��pƒ)\�zW�^��N��`�'����șT� ����G$��������������҉�=�_���r�@=���-|��?��nvw�{�o�F���I�2�jN����M�U]���J*���l�Ϣ�	a*6����*gI {
��P�X�s�B�"J0�࡭d;R���Do�.�?}oyϻD���C�.�!�07~D�v�ߏ�� ��Ϧ6]���!��	���!�D��'���j�=�
iq��׉{;�t�C>�]m6,`8!���2!�2���h��.T*TA�1FE�������� �7���Q��dS�X�"H^���s/^��|n_+<D��y�V��8��u�8�{{#"�#�;�)��2&6v���I,�F�����KN݁V)	��7ľ��Z=�j����g��C��y�$V7��ϖQ�y��"�FJ �S���8rp��1���#��cay�&f��̣��D�*����Rϒ�%�Imi��	M~�n�"�3�;hyL���\ܐ@>�;�1iv�P��4:���i.����r�ŔnКӅ�TW��qy|ۻXlXlnE�euK�b
�\�=-��u'��ύ�vFP{N�2���]����]���4N6gP���b�����k��2�J��[��BnY5�YY5,�8M����C��P�'`�I��0�?�~�����^�2���(Ju��'e�rbd �OD$d�d�T-���H�s���0��Q��g��s�>9W���չ[�j����`K6� ��af���,00s����{��� <���`��IN�,Y9��
-u��r����<���e���./���������{��IҾ�=<��e<w����䀸�}v�v@ �o�3����v��za��w��E���	�"��3�O1����K�?� ��c2j`�!�p8�N�-������/=��OPÌӧ.bu5�f�&����D�����A�~�L��!`�.'~^_ =w�bS9t9�z#����P8,'50���C��4��Ʊ�+�/m����S�8��&�v0"���g�︡��hQo�s&�W�Ҵ����Q�kh��*P����F�4g[v�g�6�ݬG6����v۸�Ps���Obm}E�3��t���V��^��v��>��݀������8pp>����n�P��~��I� �u��Jl�a�D���E��y�b�F�6t���	ٰ�h �kȔ\�����s�o�<��2=��W�ß�"f���`E�2Ma1�{�Ɣ3H~�f���o;�����[��فs�I���W�&�P#;+�����{40u�&����}B����H�8v�#i)���~al���T��/j-�l;0����ќ��L;6uRu����2(�Ij�Z���'5�R�����������_�/���8��Ѓ�51�N�w��P�y�y�~��X m�B�V�&�t�#��te�J�X�-���b0יV�����G{8?��x�����ә�k� +D.��x�ɪ�bb�"��P��0�E���@MNj��)�`}ɫA���5>R�c���"�{bӻ��u������=�".�7�I���8��#������%��a6=��,�Z��\4���ӭ��sd�o��������Ϟ|r������s߼������jx���::����<�T�I��B4�0�m\�/<�Ks3X_�ʫ?Ob���Vø.�\�Sk1����[����#/��\m�����+E�G�4�hUj�ynO>&�z[�*�����+e��KOc���@�����06��;�P0�D,�V��;n;�_��q��.�庶���_~�/��Б1�۷����6����z@��u�L2�+��SO�@��䤦?\�[�N��8���O�B�V�D����X,���\�<'����)M+0��p����-���ć`���#�:�\}4�mM��w󡡘'�����H�/���f�:3�vfID�.Ć���c	IA���f��� pG�ſ6����,�-�(�;	���c������R�?Z�	ǆ�5����r�q��!pE�.d�kop�(��Z�����z;kU"@�ნKV�ty�<m�ݶG�Ė���qr�����a�E� U�ӗ��Z@�o�c�4�"=�Kk�^AOcCQ��9���iD�}Yű)�)F�k��ŕ�%<��I�,�T��C�Ĵ�\Й��ȴ.=��G`��-Z@�I��T��\�]^�~��r+W3���u�#1����`L9 ;0�u� �mK|\��ౢ(Vk8s�2�:}�����-��tX1�׬bl0���7�vZ�l��3�.cfq]�7���#Y-rzi(�b��A,�H*�S���F,�}%{�R���~u���^?�s3Kz��4�A�)�*��Ɔ�طg;vL�(�V+H�L3+A����R���0��C��@���s#��G7��\lH�z�1=G%W�¨Rkb�PW0}�O��E��/��%*?+�!$�p�    IDAT͆@�W�kClH54�|U��d�L��T!Kw�z�Gѭg���[��X4���Jm�����3Q�vᥕc�<�n߂����D�n:� 
Q�����Z/��ř�%Ѽ���iLUk z�C����J;�\�FA���{�kkޞ��d�@�ւ��1.������E̯�s	Ei��C�CD�������f�%��HЇ��al�:�x:�Fx���xaV�%����9�+a�DJ�t[��!h�kBؔ5:���x�7q����!`SI"�P�N�5� �'n
�R3g_��v
�,�A_���Hn�9�E�=��D[�F��G���I�uQfA�ZJ��j}�����r�>Â�_tk�L��_�4>�׵ڰ�D�?�T,�����E���rHz2�{DHv��h��hW���xF����J���vރɉ�����S�L��j��[a�tj3p��d �=��t�_s�HC%�ۧ��X��y��J�M���X�� �{��+�q�����w�����-O#��IĊ������P�R�b|�����{�혞Jh��}Go"/�NK`LG!�N��.c1I��s�C���Kp�S�I6u�v�1�Q�+̉�!�	ʫ"�J!�4:���xF�}'�/�ZJ�ak3x&��?��Ԁ1������Em6�!O>����G������!ٷ�VŅE��\9�:ξ�
�kX��W�hW�
u��H�FB��Q�Bc���}��ͨ^.�Q.�����@kv�wDH���0�O�?ۮ���p�����؈��2�d��FB�<���tI�	E�Ə����\p�H��#22�ԶiDw��Cxkq�<�"�8��V�Ӹ�λE"Z;��G��B�DZ�����n_�~}W-/�{{��Vssw���G��o�x��������S{#��?�kš��@�E�ih���	�C	�p3����U�³^ɨ_;)�/]�5����`bH�"�==���ҵ���KU�÷^ƙ��4����05z�
ʖ�"�mvC@���c�h
;�GQX�����:.�xE�!�C����g�dC�D�ʥ5$�!��}������b��1=o�����㨕˸���|�&ټɝ���imH�P�zI�����*���66"S�;DbwJ>���H!�t"�?R�:��(�#����y.�?���x�Y��	"cHn�)/��P���+�A�a�l"�0"���/n
���=�T�X�p˗/����)�Nd�l�S(O��/��&gq&�*�3�s�����o&�ȶ�c�����~��Ҏ�{ 6���Q|���Ɖ���M6l9:�q،ln G��tNSO9�$��ݫK���-Ca���TxK;+�Zۍ��x��斳h�9�6��F�f�6[z�]ۇ1�#���i��':Pot�����ˋx��re�X��L�d�`&��F~_��'��&�%f�a�֐���D�Y\er�,��7W�+y��j�&Ǳ��c���x���Xoci�.z��Wf�/W%���:����&g�nI�=zxұ :�:���G����WpavA�
���a@}6���Ω$�������Ug$C,��A.-���
R}N��E��E(�Ԕ����v�~��s��߳�i�h3G�L^�LCmt�-50�����e����hv�&U�V�9��d؏�Q�MOP�ܓ�'�28+mTi�:��������欓bh�8e�k(���y��+����'����n�M)��x����~GN�!��k�`���s�y�v�
N_����|p"�>�n�������5:� :=?�W�8q�
^>5�R�����'�����²T)�T���hY�:#���[0=���T3
�^����t\xC���St��pˣb��Dg ݎ�C��L�chh}��kE�__�t�VW�L#���jd (jގ�q��p���P��k1�ǟ?�+�Y�cC�y�Fh4�\��q�q��5Q�>&d�F��nsa�4	N���8wh(Π�A�d�i�~;C�k��Jw�!`q+'�m�k�������L�{�QbgO41<FOf6J�H9�-l::D�A	�k�2�y�)ds�GtRx M>�	#=�RF�J)ò�	u�C�v�L|t�|n�g��i�j�jقF�P���$����1�y-��f�b��q(9B�]����<][�6�,��������g:|&[���38�(���9��x���v�>T��m��n������C�ݍ#��KP]�TЪ�Œ ����ءrBM[_0ͥfҮ�\�tXG���&^c;J�D:�I!kJ���XM��md29Q��ȼs�.�޽Cף'3�>��6¡ F��߀�,��A��S�z�Á.B�����i���~5��k�S0�g�{O<����n����Pb����
UW��<W��0���UTYu:�z���14����B��A-�����F��Ok.��o�usYt�#���Oq~��R./t҇IՒ��X�6�-�'��An�L�G�o�E\[�ZSk��Q�_��LDy�������[�"�SHON"26���R��7���ko����x�g���_G��ħ��Kx���(�=�F���Ā���v��^�Z�����&��w��[���>��M���	T�g����g�z����'�x8K����?�ƽ����MA�DS�dd�i�߆����S:3�P�z���,f��h2�����D�-&h�U��ZƗ�y�g�hb@7L�c�)EŜ
�v���@�݂7�Ŷ�lIE�*dq���p�سX�9��]|��fA��@��^A̤�Ѓ�XZ���Q����z�~��4��fV�E[Q4'^��x��9j^?je�E����ӧ�o}�/_���68p��c�a��#ڐN3|���O6yq�]& ���C�|����?�,�כ�&���I ��@<9�������A�zN*Z�"�R�����1��M̝9��gO��@M W����pP ��n�&�B_��	`�����k���P��?�1_Q�8x0q�ux�?�P,�"T�n�}#��{'�٣��h�9��N�b{�4����C���*]�gC�5�MatdÃIAÞ^M����� ���!��'ܞ Z=�ke,,�Eʗ����Z׃ɔ�ϡD[�bt�"�,OS�x�9ג��enA�J�f�pqv	kk%���=m���z�x0�19>���wb��V}@�ҒƁ��?�Z9��&G���]^s؉H�hĤo�aȋ�Uf���N_�����le�I����x���.RQ�pp7�m�E*7� \��F˫���C��u�ɳ}r�� �=Z�����I#�617&�RL�9�����`����,�Փ�E��Y��A�����Vp7ѪD�ڹ}vMbd(����c&\�I��\�w��p��P7Q攳�E��>�Ncz�(vNcb0��.,T�-��}t���WKu	��Vr(䉦�Thp��|]��^��% �r��ܰ�4�/%ɵr�@o�� n;�.N�˴S�$�Ax!^�]�s��ą�EcI�����Q�d2��n=�]�)��eT��`a艠��cvn�^;�7/�#���V�9�4n)���FE��pc(�R�r������w�q�M�)!V
��ƻ��Z����\�ɳ�(�u��`�;-DCA�S1��-u8G�!�1�N`p0���|��ӧgx�������&�b'�o!���C�qp�V9��+U��-x��]k���g�)�J�*	�G��n�|b;�p�m���V�� �1�Po����wc߱o��v�$�	p�=c-���h��wRm7��&���=�������~�~���c��4J�n�7��D<���4���}�i��Y�~�Ay[t��E��6�P��AD͚����.�PXBmmѨe�,�C�ȅ�ڲ]�((fdk�L�e�A������m~��E���5��ϔ��_+d�tQ稤[��-y�MN�}A$�i���j�dR)�lʤ�Y����GċF�h��� 또衵bYg	�$�$�g����t�ph�I�u6��|�{�R�'v��s�PX��;�T�����1a���t##CI#����_��v���������'��c�=�3o߾=��۱cz�\�?�8.���F��ӻ�qǝw�=q��9d2Y�KU\��E�VŖ-cL&ЪT�_\���<<�&��>�Z��ɠ��(g��V+H�����81>$�x~m��e�YQ�R��RI$�Q�Q��+�g�ٲ�>bXl<��ˣ^%��\7R���w���&S�~� l0��r���Ve�D\%5�b��޶���Y�LF`KDeF��(�5}n)��ky�[-୙E\-V0�g/~�����^Ժ������سX�4P�yP�V�%V�P��R@]���>"4�,e������������?}868t��?���3�a>�����FQ]M�^����΀��o,����)0�k�P�e�T��\�U����n/^=���������*��7҄����{]n�|6e��)�C~�-�
+8��8�Ƌ���ş��1�>'Ђ��Pb!᣺
��;�q�������C�pÑ��y#/���X$d
-{b�iD�\��N�_���믿��~�{�K޶���	��Ƌ��U>X�'�L��1�	.^:1�Z\]Z��/-��g^ų�N�4��!=�ՖO�!�?nh
n7Ztm�[9����F�~M�Zj���`��\>�&�ͨ!ཥ{�l��^�>�l��#�3��J�{0��������Z�X@��w��O�
 ��d��aG$H�n���M����؎�̵�&�rz_��Ά�p���o����mc�|�ۜ��0�"匱)hfL���s�Q�[JÅ�\+��lh����[��2�S[0�"u��b�U��Հ�G��	�aC����	t��8��)h��@�͉�s�Ӆ��J%��3"w�ϗ��S��i	�D��X�R��֟d�A۶�#��ϭ7 ,�v��W$$�0�!/�tJɎ���D�HX�!��XtO��`yh�i����QC�аfe�@V[��_��ª��VH0~~�͑��ST[F$l�W3��h��M\^Z�[�g������LD�i��裎V���4���q��>�t,��DD� ZO��������ui~^�%��R$cH���u�Ɩ�ۖa�Q�2��r�X��q���2f��(0��O.���{���`�f�7V�b�Ԅx�\Ԉ���8�E�ܰ
�^?-�P�V��C��'�r8}�*�:�2�҃H��B㪹$=-�{�a<t�~ԫ*z=_��Wf�����TI���B�6�ۑ#��f��F�"�d<"�F���Pԋw�u��"ȩ0�9��Q����N_�Õ�����^��,ko!�A<yŹ^���H���D���\Z]��W�`-���X(�@����*�%��]�:OO��e�gE�\��m���)/���+�:�V͞[�!�&Ҷ8E��	�r��"�LeM��Ї��i
�}�G�q���_��ۺ��h�ӌ�$�{��蝜�o�{���� 9e��|���ޝ�B`S07^��?e�L��f�0��8
�,^~�%Y�Fcaqۙ���9A�P0�����?�
G��y0�Qk���A�h�`��Y)E�t���u@ɱ����9�O�u)@m���=ƵK�R��{��f� �<��U��d���L�_T�P��k6�D[R��]��i�����ф��H��db�!��-J�}r�e����G���ߩ�P��*cSʟw� ���1br��I��>��q#j�AP��x��Z�� ҵ�]o�����_���|���_}�/T���a<��;�K���J~����~�RQ�mw܊���oK���>�'�|Z{q&W�`V�N����D}&��H������z�/�y��~���	=$�5�_}�6*+k�-]ՠ#�em�p:�8'����Dq�J��j�2�N��D�\A�Rٸf\��R�>pݐ�f�:6�2����y,Fl.�*��+h��#6�T#�aJ4�p2	w$��7�+�".�q~%��L�H�o������=۰���׾���ԋ�t=(�,�Tj���rh�#���Y�a�y�f~��>�����'�w�����'��ԁ���?��@"q讻ߦM��z�^nBl�ItQ'���� �
���$��Pz �N�W3�}�.��y-rf]]%�z��4�hy�8v*���.\m�g�L	~e��9Tp���5�v���������dv(�^%�%�qh��[@�.q�oP�����ӂaC���-�����D�[�p���p���e�N�16:��dRi�T�+y��f�+g�Bh.�)E�/��j��}�~\�����(�,�����0�������|���Ɨ�>.�f��$�M 9�Go��u$t�S(G��b�g�'�*�맩�ϭ�>NK9���j.��P�jg�3�6S`��������m�����96F�AKZ664�Y7aV
�zmxRQ��F��=�Z���w����l��L�K��	!Dȃդ�f�Nt ~����g
�;>��JEל4��;�c�/�5z�W	���Zp�i�Ǣ���69�a��-��XY+`��Uܲ�طk��\W���c��%��ioIj�������)����%��0�l��6}�e�kփ��Us�uQ�����(�L�@<A��{��H�RC���M[_=ģ1]C¥�JK�P+@�M����̕�87��r�I�9!���=�G�H&��twL�3%�@�S���g[]
y��E�b�]��uhW��(�Z��v��F3/�Ͼ�;096��D�<��.�-bna�
� |� �tQbz�b����TZr�aS��ae#)��:��'�6�	���ԑ3S�RG ��@Tk�K
 �Lϔղ	"�P�t�.�����X`�V��l����oB|�wnv�b�%�0�֕v�F���6Q6p�z���F8�g�wO��eH�g���#�k����![i"�Ji��*g��p��}x�}7�R)�֨�����%���v��?�N����m���F��T��mY����ØJ��7ioK��ۥ!��zA��:��.�\����*�u1��Y��#a�¤K@���p\�[ę��X[���F��'04��֩A,̝��oz���F�����Z&�'1���O*��֧��!�A�
I�%�����9��3�yS���Q������	�)6-�]���;�e���4D�6֎��d7�_VS��&�tc�#��L����@���oTJ��H�Q���ꫯ��N���U=�S8�,�N��@9�ux6���b���Q�ca�8]�_D.W��m ���D��B96=ܧX�K{�1�K� [StҕE�2�q�N��r��{�5E���t��vP�Yu�1���Rp�a�K_�Q�@*����DC*��k��>K�a��]dz��k�g�3�rG��P�t�-��)�L��)j��p��!��dd�9��ٷ*n�): QN�k���?���×���_�;�m��A|�#����ӟ�|�_Ԛ����7�!�s�_���x���f��y���r!߿�h!��b<��x$��hq�;�-x:R*��L�RC�c���^��c��$,ҟ�Σ�YA�Z���Ha�f+��h'�n�R)��=���B�B��d����e@��@=�=�j�z���Q6����<Ȧ�B0ArhHZ�e!����,)"XA�X�vG��bǍ��6.�P�������w"0���������K_}�fVPuQ�%"�}���-RBe�n�M��iVμ�mw|���ÿ}�Ǫ!��o<s�>������C����g��`����=��6�Pf߃H,��h�jc�~�}���m�x���a��
n��NL�ڃj��D�N*MX����1�y�u|��Oaf�Wxnz���Fٷ�6/��yhq.N=8��|�I�$3��ma��[���q�� U�-M�h�����%�������?���j
c[�1<���p
{�Mc��-H�⽱�S�+�I�-S&�u�a�z�5|�������;��7�`�mX��P47uN.����6��'��4X    IDATTZ(W��Ǟ���gp�r#<�c�7`xb��c9��
��X��}��-&�Rsa͘���k�أ�����ʅ,�;���f�I��^C�Q�e�)�v<0�va'q7��'0�&8�um���ڦ�=�ƽ�y7�!�4|����
؜Iq_�Zl�w�ɺM`��6�mذճ5LT��j: m��ٜ������@��͇�`d�!��,�C�IwO�:���]�Ut{�Z-+�b��ٙ��/jJ��I뱡!��E��GC���{M<�A���IAy:��(�\XX�ayuM�'�� &@ٿ(��n|xiy��:��ϩU:����qL� �-R-�p��QA�h�������OJJ�RM:���dJ��^�ciPS�\,J���nI�s�v�@*a��]6�nS�(n�B�.Ԥ��u,g
�_\G&_TC�X�	Q"
��秸�S�����7>2���&�J�f��x�Ξ��B8�'/֍�/**���DpP���G
(,H�0>6��-CH����d�n�g�C����
����tx
�u�U���U�E�t�r���ǩ3qu5��7��N�7�Y����gv&�δ���J�f�´�9��ZJ�C�����A�|dF�Ӂ�8�s�gq��<.���"�����γ� ��3���8�~�!�E8E�����Wp��U\],��
ˉ�SNY"�a��R���-Q��D�~9ME"^��:��T��@݀�.�\����f��9������z��^D!�K���30;��z��'����
Z�>�� �I�x�>��X^�E�	���m)Q8N}����X"�/-�����Zn?����p�%��@���8zg�QaB������k��k�nNc���O�^���%;��h�F#a#��k� �k��db�V�|��׆��C51�C��c�'H�B��(J�eC�u�8J�"�?�\!o���4j�>��B��6��\�\}�EQ>ʭ�'�~v�[�m�ԶI�o���ŲN�9Q7<y��d$�@ ��6���B��dêtk�F�^0I�ױ�|Ea�	�s�x�ו�?��Dar�;�l�'p�����m�>s����fq2N:#�1���|���&bFiNb
S�Ƙ��T`~��:�����h�,W��s���Z�����E�UD*��J�v���!��+��:4*i�P̮�C�����������#_{DV�|��r~�~S��������zDZ�R����}>���\�̧�Ǐ���pS�I�VU��#�c�\�>?��I�'�HG��z�f)��ׅ^��z� 7�+�n�h������ j�
k+X[�*w!�p�5��azjB��B�R�rE�/��#��A�׋�*-ݙ��4�����Õ3�[���	��a�щ\DХM�!�@�D�݇;D�ӗ���!G���r����?��]���ƣ�L������b_}�	{��V�
&�7�h�k�e�Yc�b��tZ�YJ�f��{�~�G��{���UC�'�z���٧����u��qT�}UJ����?�Dr&�I��L
L-�e�I�߾�'qh�.��O���9:|7�t�����v��{GѴ�'^Z�_~�	\�zJm��1�������B����4
�YI�`sb�-�+���P �R��9��y,�K	�^R��E���⮹i�c,4B:��ō�E��Ci$RQ'059������G02�@�]f��"u��F<`n��]8�8z��޳S�~���sgRc��B7T×��A�_;�?����ﾈ��^����SX��Piӥ)��,���/�M�t����&0��Jh�藩{������Ϡ8;��zP�0��ף�6U0,�9qv@(�Y	��&��ZC`����٥�u���;[����<D_4���jL3p�!��p?g�ƢcA�����h�bY�1�����D�|(��,���EG�@79(���g�ɮ
꥾�ORAX���nB1�-R �r�,�j:Rq���<jx~��O�A�TR�p?�K%mb�r����=�g!&������ghQ�I�:m;q��A�%È�L�'T>+&`��2�9c��'<�+U�|�es(U�H���ġk�6nN����i��&��`�t2�F��:q�>D�1��1��b���]͉�_op��7<��_p�iA��p��FØ���萊h'�:�����[Q�Q�{��5L��:t�`�g� C��~K�
x�X®�ea�	�I�Ɔ���8�˩�@���.\ҫ�E��fQ��� �Ei*������|��A��M��Xtj!T��LC���gq�ڔ���p7^��'R���^�3%�y�D�ي+�RO�?�h��,��16ǭ�^�T�..,��(�8u�<�\YB�B���\�L1y�z�9)��:��w߾HDج呈�1��b(`Ic�s�U���x.W�*$t�����r�����<2�ZI�,n|�F�!������
�z�����o�#=91��w�+�V��i5�s�U�Z3D}��P�UW�֔��7��4��L�,ę_D&�Y%2dx"�lr��^dL���iL��â��Ź��q����Z8E���� ��Ҵ+!��6��ͦ�*;��S�;(���M�a��|]5�N�gGtFx]��݅����g�U�Z�s���EMq��H�(ѭ7E�3	�&o��e��Bj0.�7�˗/��P�0��nCNF�줍y��*�;J��--�I��i�p3.�.�5����I����z8��#�/���
`�z	I�١bB8��^Ϥ�6�H�����.6l�ȳo�yZ��~t[]9�M��_�Qw(�L�)�.Rgi�KD����lv�D]x��SC�� ��Pc��YB�,B�y
��w5��(��p�������m�x�|�S��׿�u�c<�n��V|����(C���G���R}����w�w~��5t���k����WDVI�k)�Y
���m��X���H�����tЏ0�z-�uk��'�k�5�rںe�۶b � y�H��
��<��>/&G��$��QN'9�'p������W�S�T6�=���?�=�I-��C Zw0��
G��3�{d;�P\v�j0��pG��R��@�l�ky�Ã�>����!�c5ˍ���x��sx�/���%d+��J;��
�P��n��e`M���1<��{��_��_��B��������|��j�����$\ͺ�Xg�8�l.j�����0ȉԶQ|�����x�����k���u���{PkU�jW�e")_+���{~���R
":8-�C�f
M.�_����X�p.v��,9ODC�3X��@iu/?�.�A�Yj%mJdC�!�i�0���Z�ŉ��<��z4 T��p:���Sسs+F����4��)5S�z�����(泘ޱL:4�M����4��+�9��:�%GvN]�����{x���HN�ǎ�c��ë�/��"�L�Y� �1K���(q��b�K���8�Ǵ���+X=w��EX�ڍ��T>�?ѡ�O�k�7wX��.C܊�!�x�Lk�UCJ�����)��=t�Q��އ����[W���Z�3��1�99͞�{�J�����_�4���}l���7'�6��"̞�qs�&�k�099��"�� �]��`�
i�Oz�H���V�XK�]ȞF�ӱ�#	��yH%+�~�F�h����z��f۫D_�!Y��;� �5[X̓Q0�)�X�󳓊�1�L���DCj��[(R�Ԑ�Z~5[h�rexش�5���;B,M�!�.�?�#�`��?/Ұ�$���������Xi [�
�eȕ,Y�$k6�r�Ն�괴��[b1�R�7�$��2(���ax=!�xh+,�e�}�:�d%~1�9�o�ը�ݬ!��ar��G�h�5��Z�x͖[�j�Y:q��M9Da���X[����s��]P�����Q;���r
5�n���Y�*$m����.7�6יT�:�e���Ά �a��V��1�T�6����N�>���"���珙�/��9u�6d���ƽ{����� �	�_(��c�c~n>?Ù"�B�Y��Ec��^$��_(�š��e��DZ��LqN��6|�9A�됷��!V��y�zq�T�A�������-9й��s�?��W�"�+#�i�P��v��\���55 �ǣ�=�`i���j4�.P(����K������U�/��3��*)ņ�Z����j�ۚSp;�}�����A��懄�P�":��:���%���k���i,d�n�r�W���5v���KT��y��%ҧ��&��Ҥ�SuN�����L%�X����o���ـ��0�Hi6��4ѭ��rPǜ���`��֤��`:�b�{H���(�'�+l����}*:�ϭ�r�g�9�����ý7��D��Z���/��iL���%|]f!)��E$��?��<���S��b(ML�&EZ�F��	�κ�д[�j Hg<f�,�iT���Z6�>B��&�<w��xF�y�k�?΀66���n6�.DU�^9�l�{5<K�/,�����Q��h5����=��G>����.�O��|�ߐ<��;�����ɿ�k<�oJ����S��)���>�` ������G5L�~W�+hZ�*e�x�]X�2nR� B�3�j��+%Q�9���h��5�[��� vL�a"�Bq}�|���C�RA�U�����b@a2?���Btz*�Ir�7�ܢN��L���-�\P�H�_}�(i���<l���:3�z7�.DFR������7�^����"4�C; �}��A,�w��{O=�㯟Ʃ���Zh��@���VWNFހAvi���m�iHf^C�������?����7_8�����UC0:��lt*a0����9�7�_��C�ڐ�w<a��q�ﾻq����t�
�|�$Fp���h������4�#���A���s�/�ӟWs�c��@WaE�_-�"�g+m"]mi�o���aaі�?�U�s���S���^x�;�@;RZ�lЯ��]�+	��Z@�v�jI��T:�P��!mq�#A�~����)LOOcr|�x�v�F�c�<��K��1�=�v�J�W�:7lt��Wѵ)KWM��<�Z��ssx��E�b(��87��\����	u�m�RTı�����! _�'-�(p���V^�`���s�p���6*�V=�)���'�f�jN�lm�G�' �0��@��VZ��攚��ǃ�������$����hr��ٱ�sH�.�G�?�BK�l�|���@�Y�kA���<�,i���^+��ÇɎ<pk�q��$
�(M?�czd�L�9i�磆�O{��i�	�D�wP��&� ���H�N�rS����J�Ɛ�
v�=i�Y=I�g��������!���H���ÐT8�{��m�<*�ɝ��1�J�}�sIZ�2�Ic���z��#U����S�C�HK��ɍ�g!��m�R��Zk*������,$䳭��N3h uD�����ę�v[6?���~Q�������sȠ t"��6jբ�nʵ͵��M�I<����1Fl�}���bmmM�|��=����%Z����QL���*������=�u�ϝ��\�����m���j);��u�mNa�����^]\��jmX�4��}��I�6��%TjY�A:| {voמt��
��t�L�� �~>�"+_;��r}�>�64:��� ��.��aj< �TK���
;��h���0BK~�`8�h� .��ȬgU��v0FZ!�) .^�ًW�J�^ϭ��&������ۄ���`�L���'��f�\��م�[}DÈ![�`~iU�qf|N��������T�������_,86ڛ~�>�9����w��ym�b��(�|��E�JT�?ژ8M�66LZu�.���i��7͉��$?�<mj�$�1�2�j����l4��<\�n��i7ѪT��G]��{����GMa�;wMa��	Y���&�� ��L����C�����÷w�!����.
WWHQ"GG��D����?;;��0�/����������n؋J�����5��64�Ȑ�x<�}����u��z�ͬ���u���%��:Zg��셹�=�"��E�P]��&��_y��#�NP�D�23#�d<�l&��Z�h�z]d���u�1�|14�h�_C�����A��/���Ͼ���N^���>*g"�N�Ft�=wȁ��O<��'O����&�s�=ǳ/��/��/���+rW�!C�� K?�!A�s�h�Ҭ#�c8J�Џ�4��Х�F�uN����hM*��2Q}A"�ԔQG����i��YGne�b�3DlD"յO2���3�P쮍��CP5�t�j�^�2MAzpY^�,�jZڌF	�q�{md�%�[}�b)D�	x�f�j�j�6�k
ض�����L(��@��:��}�1��-c=WG�� VXa�e&۳q�]4�o�Ԍ����<O5��O��=�~䋿���6�����!������-�����I�U�qJ�B�Dg-$�.[SD��
".�RCp�mסWf/.��+bppP~���ʷ,��������<�����R���d�9�1^�t�PC���5.j��.$?y����vTK����o��μv�䟐���M�pʊ�1�|����A������+QgW��*�r�������j�}�y�hB�� �i!`��1�r��߷S�Ҟ6�.\�>z>n
$Pз%(KJ6�/=r
o�[F��B���|���]����ot@������x��G��-ѓ�<fO����3�W�J�U����D�����3�(ͦ�( R�@��Ŭ��m6��x����N�q��[���LCpumm;Q�PH���֕s����-Z��>�γb�w��2@�4����s`���Np�������;�~�<p|�up�!���vp�sTh�9超����j����M��c/�i<�~�k�g�O!3����r�����]�E�3&>��Ιr���+:m��o��^�𾈊d�٩S :����4�g��Si����>qܔ6ayiK�-�¼W��#Wӆ�IQ���^ۮh�a���''��s6��S�}pȔp���ҫp�.�~�>�5>�@�S+Q-LpC�14f���2�ev�#��d^����$��pLa5�>��sr�Ϧ炰�M%�L��(��a�E��d6��2�ʙ�I�1�6��gC�f���Z�EoǬQQ%xo�A5_D)(��ǵ�9j`Zuԫyt{5���a�]\�<��匚�h4�)8���7���/:��R9�=�{��P�����m�(�汴�h(!���䗅$���59�޴_�ǒ(W+������&�&0�e�XTڎ��%�/-I�BZ�2������M7�M7�0i�Bz�RD�Ҡ� �Á��"2�%,�籴�A�ц7��Y��|M�x����8�2ǭD��Xn>��P���恄s�9���%��I���{�f'#���}�F�4t��Wg_s�x���GyM�;S#V5��� 3�U�T���a���d��U����J����S�cmyA�d�P�J�,���EL&���f�T�DD|��_����.��'�!��v���WHI%e�L����I�醳���m���8�;��u����Kp�u���h(�͘vB~\�]�?}����w�@��B<9�ip��������k�ݦC��0�އ��y+n��0҉�PG��y}B�1�G����q#b��ba��l���q�"�9Tkh3���&%@����C��k�����cnv	1�������f�k�~�w~�x�v��$71��^X!&����3j'�X1h6�o��c���~'N��/���B�n��x���B�`���Ǎ�?��P �mC��s���X\�}��s�B���<ڭ��YXC<�G��G:5�~��e�W�U'9} #7a�D�6ٌ�A��o3 ݠ�fXi�Y��Z�<�15�'<+��{-,�����#�Jcxh��4��0���k�B4�s7Fv�C/1�~j��'/���'�ǋ�^C��W>M��4������8~^b��    IDATc�ϳ�::j�H�%�F��n�����}�����b��?|��hC𧏼|������\����D�\L
�x�:�b�9}�t�� �e;ǒx�����[�����&��qs)ReC@�;k:��{�|�����<�1�^�`1�ž��=�Q�ȀN'�DP�h��T.��_��=I`��l�N��^����x�<@>�Bi��7�^ZŸ(��aE#r�`S�~�D!=�;6�g�m�Fd`09NS��v�Ѩ�U�#��!7؉����m�8��m�M ��S21))���_^x=��}������/O ��@$�/L4�"d/�L��H�.�X�x,�>YBa���+�"�AHn4�%5s�O�_b07%�z�&u�T*�S���̦�>��l�ٜw<�ʙ� ��)Z~5�NDq�=�n ��! ��1/b᭿��&�׏6�D�ݙ@r3 ��M���I��D��{x�8S�%S�U؉�>Ŀg5`0�s�"j��|��ۈ	?�C���M"v�F$��B���(�א<YM#Y �I�lN6Q8�g��i��i��-CVv���E�f\rM�5uDߢ���tz���g�n��|s�ߘ|k
Kʘ�۫�н67l�0n��7!���h�,)�j�fN�g���?C�Y���<�w5|��Y(̣SQM�"S����tS��1'Eͦ�M�mG��޿YC����Zu�T:<r�?���hj���ϝ�RO���b(�{����I���c�G�'�����9lN�7ܖ��6( )�>e��ى�3N��IPI���3
)�.�y�>��j�|Q�@8���
TsWl;a)���z<Ba���2� ��-"���Y�X"�����T������R;ʵ��e~NR��=�J��6@T8�z���EMȎ�#�#�vU����a!9�֧N�ѳǴ��z^�^�# @��a���@�n$���}���ZW�\��ᗹ�5�Ú-��|
o�8"X���cCp�b�������&R��.d���zQڌ8?���k;T$�z�<�����i6$�Vrﵟ�P��`:���%�%Q��DH?\[*0�Jb����8w�
�
�t�
�P��Ѩ�p��C��G~����q�S�)��ك؀�i�glz��G�٤b��[4����C�<;�?�=�h�I��@���M�����|/��=�U<^���h�FE�/�>�3?����6�xx?�4/�QN'��d��p���&�kC%�?�����h�**�a<�3wXg��h��d �>��0���|�<�«�-�Q)1p���e�p� ���;����M>�	�8�\Y5J��Z��h�<��H��-lm�@4:����Q<�w_�Z��V
ylsߕً�fY��[��!\�k'RJ+�M&�k��Ye֖q��9d�W�����߇X ��dt
dmZ�SP\D�hJ��Z&HJ"�U04�D:!��YeQ6M��m�}S��A��Q�;�d6\=d����ʨFrx�d�XWV:�����jǅ�zg�p��9�~�<��`���� ._�f����|?ls�V�\��q�SD��x�}������?�yo�����hC���|�����|�Գ��F��$�	!w.sj)Y��m��qc�� ~�����Ƅ�_ZE�TV��S�@���+���s����(C�����'�#���h�tKv}�ЍK��K�	�7����H-b� ���x�]B,�C<�Bu}�?�$.�8�Zf���[���DI~���#M�b=�G4G<�ւc'JGA�#L��G/f#��D������`*r(k��r�!<�нؿo���1Ӆ���Vn���ᱧO��L�kMdJ.�"i$��55�D���ϵ���ߚ00M�'{t� /�Ԑ���)��,������.��KJ-a��������"��7����z����Hx�X��DRrM{�hC�XG��Fܘ__Cop;g�Psl�"Ûw�h�@s��7�y��s eN�w�h5�9h��F�V�o��Й�I�����Z�qMɩ�\�!�k���j�ɟ	�Ѽ�1�[t.1��-����o��D�v{FwD��Ԑ��i4TH'|.���257.1*�mk\��P�VE���F����'즀�
�k9��UG���p�L����.5�j���b�)���6�L���kſsP����E����P+�i���0���-j�B�LPfo��ȧ�ܦ����x�w�9EU�a6���R�d&Nא�����;�J�MɰΔ֡��&��R�)��arl'9Ø���Fw�v��㇛6���f�#'�_j,l���)״g��� �i"�$�e�X9���O�<݂��e��Ws�k�� �:�:h4���Xt�"�ד�����4Xκ�wS�K�g��Q�LU8���c�;D��Ա�`A�$A^O�Z��%��ѱI�ܹ[� \���8`��zx�D�4�r������A�[���;q��.]�7޸��.���ĵh�k��c�s-c@͍��4�,W���#^c�\\[7��b	T�R�0�4���ݔ����+�cf��5���h8�����?҂�#'�������_x�\�@ >6�ժ&�a��vlZ�0k�=gl:m���q��7���p���R�F}����6�M��m�A����}S&��D�m�E��K�ى���l"�+�z���!=�l��/}�[���:2��\{>�N���}��	m!��<ʥ,��/����ߏC���̊�.��z����{��O����)\�~��^'C���W>�.���lL�-��7-��4��R�������7é7����+]��#��W~���mo�Ig:,����:�H���<��������U�����ￌ�����y�d������=t9جЭ��jԐp��}x[�i4�9�l���I%cj
.�?���3r,#e�Oξ�':P���«i �P�'�d�k��tl��yr�����e������j��:���¹�^E�>T'���bhp�X�h�tV"+�!2:
w:�\ߥ`���\��󗰚)�W����j�Z�IC=�Oȸ�1�X�D��e�`��j(h�t7_��}w�S��K��&`����6��/����ߖz�����}3Y���%�2��D�.m0���*a��m#I�����ۑ_X��S�0O�ྜྷ�E�]e�7�<`7�������/�Ņ&ڞt=t���&2S"v�|�X>u���-3���Ð�>��<�u���X�.< �y�+%��Vp�Q^�L�,��S�k[Z���WZ��P����h�RIŊ(Mz^w	��b�DtM�p�H�aNB���C�Q@,������wb���������ե&.\Y��/��ϣ܊�o%a��Ix*ΫF*���=s�ІO�;7Szޓ�ۍ%��k�~�Ds+X�0���˨/�ʩ)#�0��R)g�������3�s67z�sj �<hh���K�4Rg�poj:>7泫h�<zP��Ξ�+s��7��fm ��YC�����#T�cy�b�<M���tж����Lµnl�9�Y|sh�����ms5̤���G)���iI ͢�43��j��6	S�f�(	�	�S\pZ��:�	C�Ź� ��g��5�5Ź�*~�`hk1t�i�j>�S�N�É?�]�l�����7L����s;���r*��ڻm�Cw�N�vҚ����;M�S\���,' S0�гiT�S�fϦ|yY(����~2u���6į����_ܾ�<�L���k��L�c�nNa�8�8��:D� =\lE6e<08hq4.
3�ٶ�,1h�,q%�p4�hV�ۙ۸D��i4ύy?���bR�I�`�_6��Nb[.r!M�˺���FM�V6��>�咬�����(�^���@�/l<6:"Tz�$��B����8�LZ+,��d�ZZ¶�T�9�a�?s�e�}]����4� ؛XDR{�DQ"EQ�-�O���l�qދ^b-/�8~�q�$�K,YT�Z$�E�I��@t0 �o����������<-��Y�̝{�����>��w:�D2��K`͚u�Ӈ�ʒ�gP�6�L��/�u޿�T�ꠇ*VOM��K.��T{������Q���i��+�f�hVx�<�zO4 �����:t�L�6�s���W��Y��`s�@l{��#�L�^���p*Ӡ*y�D�GI�!傒ƹB�׮V���'Cu~��t*k(fݽ^�#��2�����eT��p�-���~��᪫.Qv�Z�NZ�)�	�2��1�e5&�8�Rɽ�R�ܿ9ߵ)*��Vș���O|`�hʬ��!	����w�����������Q�cT���>'g[V�c�,.��+^��~�}�����Bł'�:�h��,9-@�:�;�*���(7?x�!��9O�'~eI-��� ��Ro�?|�{�ع}�Dˋ�J�G��k���w�"���F�S��g���$'x&pX���##�3�SK��K���>�:,sG:�sQ�I�d����"��&R�l51�L�3�۩S����0Y���-�cu1���c�?z
I�bK�vJ��RX:vL���N��J0���s٬��t~��h�.�II~4Z��5�{�*���b^���(���L��126�3�<GeLR��8V�!51��-�a|��.��ܞ�x��,�Ul�;-����*I�֛m5犣��Tbs2���3�BZ�,���a@��5���7}��?z������~��W��?��?o�F�/�یr�E�	�����j�Ь�D*F�D��֏0�N�>7/����]���}��݆����t�5N�p`��/k^zmˍ�Nb��I���j.\�) q�]t�-�si�Y�c�9}�;$�˥%,/�����߲n��w��<��xs��[�R2���T��[)�/ 72���ˌ>m�{NXnd�pHSbS $�E��@�e��eՊ#Y�s����w�k֌�*i{�/��_ū{��|�u*�!S\$hD�E<fTWwI�C=�Wv��2F�:X�I�p,d��d:���
J��K��^���νX:2�����+��Sw��ryI%|>v��ؚ��{��O�B���agƝ�$�d���?>����
׿�6�i,2��h�j�x<04�B��Z¢bDx��z�CMf,���Ohf�Z�{#����vp�l���\>�x�����~ ��m���|�������р�KM�ZHIS0��d�E)3qS&��:� G\���C��q^����^�[�#��2�*z��sɵ�*�^�f�����+>s��A���!�McCr©�Ōs�4�GOz�oo�t�st<Np�V������:�I�avЛf�lЇC�4(~��h�+�Rx���FIX(�����܊����AU��^��4�a�`�5�Gz08Ol���޶�	��{s0�U8� c��ϟb�H*�g�Ǫ �'��h6N7�A�{I�#fr�3�+LRP1�z;.��;��k�.���e�y����5Z�Hؾ#3���,c���ۺn��P�D4Z,j��h,��k����,C�\>4|���S�6�"��̑#GP)W퉽>���''T��&Q=����*��[bÂG���K�f�{x���iY;S�� ��_���u�Iq%B�Y��b��	J�Ze�2Iyw��N`�Gu�L�h�G�)��r	I�Al��t��_RB�^�M7]�_�ŏIΙ���l`v����߰w*Ẉ'E���):������mdh�HF�+��c��W�AF�%E���~��n�~�\bro��Q|�����|Dҳ��6�8>i ���lZ�����(���,^w�9x�o��/�9�y��a���0弑f��W���x&�Y�G�c�"���P/ӛ��)d"����.&G�'���A���\���<�8>�ůa����Y	��I]�j�m\�vR	��ʲ�Xm���S�O���C�-Fֆ��◑����i��G���<I���T!`���"�*f��X��>+�&�EQ���D]^F�R¦U�p�i�o�Q^�W�p�6����=Y1lw��T�a�R���E���Zd����ϣ��z��RI�g?��"���0�U��
��#EU8ټ�錳�.�Ig��l���"91�5睅v����"v9��z{�b��<��Q�(z@�,V�y�3��j$�+����3##�.R��f�L2�c�%�z�8FR�g��;~�|���hd��ݟj��?~㉫�3��%��ݰM�7t3X��<��l��Zm"֮�[YF���vW�w>>���5���F�"7X_4,��	�����.>�����9�Zĳ�Z�#��F�{�q���q���=Yrǻ@��B�N:�n
�&���eeF�i�f3X75!��~��g�p|z���K'��S[^��'%�W|>R`x�$�Q��2����3�s�Z'.��4T��S�^A�^�E�_����7n��ޱc�8H��gFO��է33���h,oʕr�2�7�K=��$�<7�LJ�9v�+��*���mT�e4��X:8������2tk�����p��^�2�q�18r�����D��Ӕ�m�[=�+n�VA'��������eR�H��QMf#HN�NS���
b�H��xpC�Ö��4c*5G�G���ɗZ�T@(41��g��4���Nм&���\y�(������Ɍ�"rMʠ�0�3ޤ1�@E������$$z,�JQǵ�{J4(����P ���.�f9aK�����D�wݣl0`Q��d��E'eXD3�a�.F]���b �2�r�M���D�-��*c�kI���A���=��qg��R��>��e@+ȥjZX �4%�b�P��^	���xt�\
��g�nܾ��
��<K:�ty�5�Ɔ����K�\��y�yo�5���Zp� N�fLiSֲ th���aŘ���C�@s�W�3�~�tٗ�?t��3u��G��Qw�(L�>:�L	����5r*�d�W�(�y��Z�FG�����ʞa��oJƚ��{��{�����&:�S�z���@���[\���*?�+=^��*�������,{�u�6���粞�'.\�4�%�2����u�6��������@�۪qe�llԗ��Oca��49͓f��N����U
sؤ�\�^:WЪ�p�W��~���K57���-�~�o���/*+�yE�+s0���~<��>���,k��HqN0��g�=>A���)�%��5'?2����#ǰm��9xTՁ���D�0�R��D�ɛg2�F��&��F�Y\t�Y8��3�\���P���y�0��elJE�{eɟ�'���O��Z�RG�TU�y�Tv�gp����3�2�r&�R���<���s_���#!�W&4�6��*j�E%Q)��UT(u�!Hn��5����3�A`/e�R��}���E���9��Yc�]�9ߪ�8��C���F��n���#yd)�@��n�J=���C�X�R��H�u��K��]�uN.�	�/�M��bE�%d��r���b?A�Mڭ�����-r'׭Q� ��F���踒Ӊ�1��I,��8Z)�G��~;��2��FV��Kcvn�rMU�|��&�@����կ@�Ca���*;4#U:�X��W����g���7}��?q�s'm�?�~�����������?_i'�/n:=���}���w�pZY/�O��֞d��N��~���X�_v)��N\~�Z�V�4W����}�L����E|��cǁ
j�1$����Ry���X"E�R�d�JH��~�b�\`�=������Z֩�h�Zg�e�Xb��i�)]���֮�S*ce�N�?��ݻp|�>�F5ₛj	����5�X:J��W�@eJ@�t#n����v�ȌOb�gb��3��\��̔C:7�~��X	�0ӓN2m��*J�%F�l**:��L�/������ټm�q�1Kj�q��3�W�X9>�:�ҩ�2o��T1AGN�,�G��YbL���1�8����e���F�AWz����Utpp���Jj���%���t�m��7    IDATӤp�Ų{;zD2�^) =����OV�5"?���a4�MƲ��"9 ��{��$�πJ"���� �|�6f���2���v�@A�����H�;n*>�-���$c5

`L��><�L�ga�gȲ(����";�E������^|R-�l4P�&UЂS7��5Ǒ/Xf�i6����2������e��^j��?�E�4�v���v-#��e~ך��q� <�z�9�3�=(�2v����)���Ѓ E&5�M�Zs6��U��Ï�z <�$��Ж9����>��;�����.5� $@ۿ�z�ϝ0�{ʚ9����(T����k\dV�����5h��g�Ϝs�Ϝ��}�᜗�":�U������c���ps���]�Ic�~b=ދd��x��k�גyҰA� �~!T��ך?��9W�5;2��^�A�����υτc�����U���< �@x�w�5E2��x�bM�� MP�#,�h�&�4�N�M���ʶ�
�,,E��_��(���r���r~�@ݩ�K���2������	�@�lQ܀�#���=��w�?	%�������D�=�6�|�>/���&�TI�#_�����I
t��UVy�ڵ�D^X*aa�&��5p�����h�%��*0K�<�# �~�f�,VD�
՚�C����s�f����F=�(�>�3 �Z����܊)�ߪ1	G*��X��U�������{~l���w�xt�V��/|Ͽ���6&�+E���̪�H�|H�b���@���S	��1��k����Ϭ�ɢ�J����� �"��$��R�d?JW��
hXY*$c�0:"vu�&3)L�3�p��r�'b��Uj��3�2���T�SP�B*Р���qV�E���]z���� �ϩa���i[N�i��hn�9�c+%�,����Y��x����q	�<�������j�㨗[��9�>�:�khI>)�Q��F+�G��=Iբ�r榐IeP(d�j�@�S~杷_��>�sχ��'����7��������R;y�������0+cRB'�fr�S���:�XU��b���sq�o�EgN�U[F2�����q6g���G��Q���r��$z��� �&s��i��+��R�綍D>�V��z�j&\ɔI��%-j3�48����JiY��ѱ���($�X��a��:�Kx����ٷW�
sǎ�SZ6��h�Y)R$�9�X���0J��*n(�HԘ���Mظy2�Q��^�.�L�J�����E��B����}�����e=�hfe1d��$�J��	͊��jXN'g�Mz�r��4-�dmnz۞xG�����qU������Զ��DeȖz5�����%�hi�#�EUz��A�Qܸ���&\��۰�i`ϱ�heR �΍�{/��9f��ݬ,�0 ��e��xx��3m(l>��ឭ@
R�j��2��5vZ�س|�T�,x���(�?��`;�f�C�����@SP��x q�M���mt���@Nk �V#�=�;��J�ˋY**]*tp��W��V/4�9��ʹ�ENYp,ץ��W'|��5:�@�8�b,=���T43:�%Cω��"{V��!��~dc�Xʳg'���c��QT���Sdb���VC#+5�������"�5�%�	�D��3sE�Hc2��I�@Ф�B�u��l�(h�'�����)�f� ��i�e=g�Ư�
�*�<�~�M���eߊSc�|�(�=T�Bv�b&j8$���=��*�%UHsP�t=���f8ۡW�`�`�@UTCW+�>�gP��P@kn��+�x�
�,���w%�����m"�f`ߛ�*b����h"�i%��'��J���^�h�
M����耒�&zV�,�
A7�==+�gw��������2�d�P�Ut�T|91=��܂�űv�$����S��UE�S��7���K�UW^j ��ƾ��[����3/��l�fzt���0�)^'�g7�A�ߑ� ���cC��q�E��$rycxe��a�Z�۰^��r����T	�{1��cX�z��`N?��Ξҋ����ŪS\ �^cƹ!uD�i���i�8�J�~EU��UQ��GưR)�Y�Yi)�� 3�F
� �S=T�J�(�ܴ��x��L���n���>�.��O�:�L�j^iv�ǟ����ں�NRtY���*En�6�X�Ғ���W�[�,F��:m1JՊ�a��I=X!pW -��Ћ�)�<U�xN3QK�.ǫ�kJ��j�m1�Mc�1L
(�ۘȦp��5�85�$nu��X���B�j��ET��~��q,P��INJ��4ִ��{�\'�s�R��ʓV��}rM��i�3�w׮[��u�P�7��(�/a��1̔�HM�F~j����C#�Ś��R��}�d�jS���� -;��I�bB'�}�O;I˓�~��ݩ�V�G>�|�]o�����c���G�������������̟1q�Yht�J(Cڤ�S6�z���{)�G��Z=L$Ӹ��;n�y�&�o-#k#��]zZ*16�ā�>���ڋ����:�LW,!�	>l��\i(��S�J��J+���5��nM�Ծ�!C5�BZY�z��T��M�3S�����<���<\�e�$��)�о���SO���=�4�.�/�R*���j�5�p���(1���*����U�^��ι��4斀ٹ
L�����Pr�%R��L��h�pMsB�%�&�덂���r[l���C&���e8�l�^�����K��x�����]譜��͌���P���=א-7g���I��Д:��3-�&�;W~���3 ��M��ͷa�����Chgɷ�˚��1 ��Zڱ���7nj�iOW�	 �A�Ξ���(0�� �{So�-k$�	&fEl& `p-
����X�jieſ,���Y6��>�$�w'ne�)�+�����Y�2�D99�m�=:Pj�7��L2�1J����\���y��a����yp�\sn8�&�=s��&
�4/�3���4�a��[�p�,��7����蜉fs}�x *p'��Y�25$uP�
�z��V�������7&dB��� �^D��k�'��t$��u'������k�੒�5(N��*6���'�qSf��$��Mt�! �;u��ż<��t
9���H1���?��c��!���Bo�?	0�I��H:u'\u��%������C�?9��x��'�ao���uƤj= pRu#4���0�s�Nʈ�C���
MN����W0��`�-���x��X�X�J��i0g��֗A�sO�@�M��H�����bi��؈�g��F�%���gqp�n4���o���0��{/��
:͊T��r�����]x��0��>��K�7���4֬;�ݥ[���3;����q����<� >+�֯_���U���eq2Y�V˘�[�d:�G�C�R��F䍠�o�kT�bZ�ۄ5\�Y��f�I�n&0::�
m�^{����Ie����j�b�@�H���P��FM�ɞzE������z���&��
A�����t3���6m� U-k|g���7������̂X�]�R5ʨ��6*��Y�4i��\A��쑡�K�Mz�)����%m�oԱ��s��+���PO�W�������t�s�RF>C��b��Rq��}��a.��|��i�ԬJ���lUj���>��j��6f��2��b�8v*	A�4�驊EU��kg*^vo�W� ��x�t���J an�T�k3GQC
�USHQ)��Z68oX/ED�w���R	ե%�L�r|H5d_U��Ud�����N�J�Id�	l��ј����֟�?�;�{�?���ӟ����������
�7��߂*Cxq�-*Zq�6Rb�!�ٶ'a�R�R����*�w�M8k]��
���3�,�р����/e��,/l@vtR`Cґ������y��b�NҲ�A��	Ө"��j>�2�H�hqQg��h���C��fe�^�L���L�q��I�}7;`~vIe,Vfh���*ڤ�v*U �1ڭ�d��$�����S��@���J����B�T^��Z��T����d��lyp�%������Nl�"��`�)n[���<�H��uQ���h��0��n���
��GE�2�L[��(p�3L7j�r��ɔ!r����l��,�fzhƖ]�W�~+nx��(u��ulʡ�䯪H��w	:H�a�d��A}�:��v��YW��t��0x��Pu�L$�.Ff6�l�[�Z����n8h����E�����_ `@G	}=<$Y������ �v�l�����/ dȃ���E�"��iX���R`43SR��_&_�Sde�g`f8��)gN�ч��Tq�X�U^<{-��S�^���@b�K�?d���$x���g��CҬ����PAhҶ��A�A������@5;�0ʨ�<� �
թ*}�Y���T��:$@�QQ�Ɛ�&�o  ׽pG�>�Hf$-X�n�lB�+r�b)f�$�hN�J�!e�c���|o�\��v&df�>e4^��h��@E^W��jM�������1�Ɛ@{,�$p�~,���{ (qܡ�fB�?:�ˀ0f �e��6�9n�r�������_�|sJ��'��G3�>w5����/��CN����(p��s:��y�� �jT]V�8��V3��;bjbeB�����~��fm�^O�-�kaϮ��k�NL�[�[��O?��݃�KKK�?4������'���o3,K8����mw�	�x������D����[�_�q��,��QbYuaO�V�ʈ�m��2�+d~61�J�F�Z�
�揋D0\���9�K	��yy�Yg��.PUb߾�8zlN� ��"4�LJ�6�dU����s��(	��Ϟ��D�� ��Q�����H�d�;)Rs�����)9��d�0�B�
7���b�~�u��O�slܰ
4%_iv�Ҿ=�����Cx���p(P(%�&i)�;:�e�cb�����^�4 ^�S��b�}�z>��C�6�_<�H|	��Mn�L���F�L$PV�> ���?�vkFGq�y��+^/%DVV�PZX��	A�g"���q%�Yɨ�k��}���d�Z3d��T!e���lު?T;cS|�b�VAf��x���F]<Ɠ8tb���QdWM"�z5��+I�Q%~d�k����
ZՊ�S��[�(!�(��t}�����(ɝ��ۦ�UF�q�Ve�|�[�����G���O* ��?��=���_��~a��������7����@���+�+���q�v�Mt*u��Ҹ���p�m7�u#��K���R�aV��g�W;�W^;����s�5͞��
D���أh��ή&{�,(۹ɫ���O��I���"B���]��p�Z��%��c #�H�\ZU{�q���� ��P�ʕ�]��&&УT_�I�V�r��5�r4�T���F�d�M �����<M~?��R�^��:ԣMۆ�d�[Щ���-��(��N{fK����&u�A>`�dZY���B�WA�F�	��j��H$i3:��X���{��6T���o�8:�Mdyi�z�Hd��0�^����4uӖs;�إ2����V�kp�����܎r��׎B���J�����L<�S�ԕ��#¹��ȳ�C}w�Qn�oZ�(4�&�����R+�I�4����D�?�BU؜H�(4�w�P�����>�ܘ)��@���N�t�?�q��*8pl�j�6�!ޗ@����*�]KI �=*�|8F��Ź�'����fH���'���9����Y��̜���w��4T^P��=(�=�{�oe��+e���`�4�;��h �
Q�Ș�����Z�7r.,P�%���S�-ЋɝX��@{���~ŋ��J�{���k�3ն*�2��5z���ԃ2z��
�T�B��ԦT9
���r�r6(4��h�$��x(`�qt*ؓ��ҟl�7J�St��T�"�ۘsx?\�*���RA�#�"߿�+�R]ܚ�ɵ�����!�p{O�<���d �zBk,TD7���7��� yH�1řA�R��<��������ak�j�
��SQY1�R�_	��%���ʔ&��� E��
��.֏0�I`����S��x�ݷ����ѹY�x
�;�`�K�o���0q�e��*#k�-w܀O~�ø��T-f������[���cؽ� K���_�ɉq��<��:|� e2�h�Z�S���&�����v9������2���YUje�&b���Kq�e�I���Wwb��Zp\��G����P�?��D�rIs�k�Y#(�a|d�h(�ϊ׳����\�a�V���p�{h65�|!(,�i��Cy��V�4�$U�Š �^Z<�x��w�u>������H�����Ͻ�Ǿ�^~i�i�$��굲L�.��\\~��(����jvu�����#E6���1 �S}��R�o8���ryE=�!�3�k��e3��@�bS��[��VuR���T�hV��������Y���M1I��f�e�Ӡb$)I�������5]hq�YRO�����yFA Ek��+��ԃ��g�j�E�'���@���R������SXi ّUHgF��+2���9,5k��H��	^�T�V,y*�x��3 ��Eܜ̒	y H�����x���f}���S?��;?�ǿ�3��(C���/��}�ڹ����Ӥr�m�ٚ��Cߝk���܉n�X���y���뺫p��Q���d�Čx��c%�n<�m���ٯ=�=3�����2�I�q(�S��c�j��o��:&�YiW���>#.L�_�d��a$?��}E�}ZY�F��(YfĻM��2���
*�%�c���KeU�[U�Ԫ�(/�P��vd|Cn@��'矍/lRZ*��\����`�@,��(���h�z��3��<;XLI�So�q��t���,��Ӏ�{�ֺl���8���/�#�Q��[A�5�0��?���c���|��؃riY��~(G(U����� I-��$5��VV��@z����V\��;��m㵙Chf���� ��D��$HN�1�L�󬇧�0��2����hCe �Q:	y�:p���ԒBs�5T��{��r>Z���Ã��^ga�5�q�1����B@�𣴟�A�,���5�Z�0_��mW+؉f�# ۲ ��B�����4o�Q�f��D����TDf?%S��@%�4������^ �r������%��U�N�B�'����r:���<,�Ȑ/�/}N��ړ��0T7B�i���Ԯ���QjR��d -<�5�ea�y�1C��`JN f�U��4}���Af���
:��uoTfb�E�t�ZH�ވ(h��`�i�(��RT�H[���z��){P���q��&C�ă8Ѭ�Lʿ��S�l�ƨD�W�5�h_��� Ga]*0�Z'a����C���}ݞ��D׌�s0�S9�>&Wl4k`�g�}-��PE�Vx���JV�b��s)�|���t��s8��	X��>���P����ҺjO��#�E�2ҰT%�*�1\%Jbw��:��D:��{�c�ӏ��ξ�
\w�ͨu:8|h�^��������\�Q<{����/�ͷ��F|���(�
	�_�{ �z'���o�����s����~N߼A��+�VM�t�pM�zbaǏ׿��9���&X_�~=n��Mz�t�޳g��0��)j�?~s�X�n�;�<я���ѣ�5^#�Q����2��ǉ��V��m��b_��t6m޼�s>�F
�s�>p�O�Zq��i�><3h"�WS���LNMa���Ԥ��3���wan��^,-9L��G��7q��oǧ~��X35&�J��������}O��K8t𸜿������F	�O[�_��w��[�E��6U    IDAT��L�V�H�rH0��f���^�KU��I�eOf� V8J�e��y��łƏ��?LR�4�
�s��qh���8���9tU1.�E�gS�>���n�Z��O�-���"�ϝ�H����I�Z=��.�*�G�W����7J�=*1,,�(�d`�^E4gm��f��S��u�Z�&�lD23�D��n:�x>���
b�rtU.��\Z�̡CA 64�7�.J��7!,³�B��	���:�y�S�g�}�M��_y�K'������S�!��������_��Nzb�����"A��ߏS����V�%P�vlJ)�NS�
'Y���W㎫��M�]���$FRT�hjsϏ�����K��4^�q���8VΡ�Z�J7i\0ʍ2��p�������e�ʁf&�Z��fMU������/���4�|F��r\v�K1�C<:f-�U�	�sQ0���@v����F���$�,Sqs�aT��X�0&���R�NJ�ȬSɀRY4�4��i���߾޷PȡQ�����
�ʫ�bQ	K�c�TBcv��YZ\�k۶����@m��E�1��{�.q�������N�>�̪M�D(Ys�O����[n�MoV��;�A1G���0 d�����CV�dL�Yvp�ˀn2u�8�����C}����Lф�g2�h�^L�=���`Y��u�<�sr����!�(���(�@h�� {��m΃�<��g0��/�+~��'WB��8T?
jHݞ+~b���L�gn���o���9�U$J�� ��LAA�!<�ISճ��4����fe��,lA{-��t@�Rnh��\�Nwwe�<Hl>�}��
NӧT��ЏQZI4������A?�0�0�>u�y�KT�@�a����JG��#�dR��g%�=r噅�P��/p��W����Rҿ�7)�h��,�C��@u�п%H5��Ȼ+x JΡ�ިJC�zL<!Wa0���{X�<�gә\ўK��BA��T�h*���Lz`bh��n��Y,��g��`���$Z=�k՘G��55��%�ϡ��]���B��Ẉ���Y�n�0&����n��1�����}N@��Ku:E���v�*����"�ڇ��y�n�]�z\{��(u�ؽ{/f�cn�4�/�_�#Ɋ4��4�c��7\q~��?�7^u	����2���G����G����o�[�z��ޟ�����ȋ�@��m��]XX�=�����Y>|XA��_�w��.l\�����#�<����,��@�0}�����,yfR=���r�|.l,^�n����P,..+���sߩW+J"���kar��k�ŭ7߂��ש�w���x��`���}�Y���˥,#υVO���W���8+!�Jm��
X�vJ{��Wv�k?��{����*�
D+���7�7��'�z5q)CM��_�����xjJ+ud���(��~�t7�r~����9g��e��� =���=9ڇĈ;,k.�������~#f�j�E.���Ϗ,�<��٬��M��p~�j�ш*K$��e1"ڕ:��2�k5�g��5Vl�Y,U˪n1�*ݶ;]��u4q�wT*W�J��`�?g�^�5(��g���s�����Mn@ft-:ǓÊ ��:m͟����f���_|�Z	ٴ)N1�#�#��	��zп�(��&�XB���&���릏���y�$0�����_}���W����8:~z��J_̀z@`<~f�J��7�j$,���])��vn��R\��8��H��T��IǸz7�.UyR1<������Ɖj��z�W;ʞ�3��!%��T\�g=V��G&��o�ۨ1⬛l�K��\���L��:��&�uX�a-
E�2&G�ef��L�'%�=5ɟ�r]Y��Q��Q �}3&�51��(.�S�e3�:f��C˃�\/���M�U��>#WՐ�v~.�:(���3M�6ҩ�&m*�C���2Yѓ��c�<���;w`f�.���Z
��L������*�l�:�0g��R-�}�64KIc������7߈����6��8����֠$�fn�y3��T\�(��E'1�?nCn�9ݲ���5@�kA�yW}�^�H<<��w�C�i�j:�ud�4��l��_��U��;0�<��k��u��!bWAN���E_b�8gP  ��J���C���Q�8N*'+h��E_�q��tMAJ2
���>�;Q ��
�=��8Y�ҁ� ܠR`��A�0*�载�c�He7>��Z�.r�N����$�����������F����������T��q��/��F]:P��!��]��J3��0 ����Av;PTLrZ���0�g.`x󪼅�`؃b|d�읪�*N��p��`Z�C�|��)�p��a�>)c�b��� ���������@A@O� y7kc2�ǭ�(�N�� �r�N���a��������6
��r����2��D�<���N�ճe%1��q'���2����a��s�oE�S�U�\��/{fV�L���q��?��|�z�f�϶�������������rӎ���w�],�T�w�~�3��{7x�;�<hj_�4.��L����t�������?�kټy���ࢋ.�SO?�/}�Kؽw���Y�\�����u��a��*
�Acw&���LI��Z���ܦ� ��L*e������:����pƖ-2�z��g�����jy_|1ι�\d�#jNN�����x���%�m�d{�$�_(�;�~
_y�;X�t��Qo���8�T��{����	#y�ڨ�;x�����*^ض[ƥRUH�i��iW�zUx�x��ލ�B����@��������L �n���_�%<}|/�\����Z_f��t�)�c� �Jۖ ��Н�x��n�j����+KR��ZmVZ���Ǳ�E��}ӇgQ_�l�By�ːݶ� �N���hdKV��rh�J*�E���- %p���Dt��1Lm8]t�J�#��>'T�ׯ]���?_�˯���C���`��؉̠K�;�X� ���;%T�pS�.��%��=��;������{^�	b��~��_}�-���_��F���0~:�1���X@ЍO�A��F���\<ifV���Jj )��8�&��sq��c�d��.
��8��,4�i ������>��s=�G7a�ƇM|\��#�F�]���u�ͬ���r�nD���:�8L.��a˗��:�Y�����X��u0Q6����e�&�uFÌz�WP�6U�'g�J�$�aMM�)k���6e��6V���������(�U5MMLh�Z���L�e���b-XF�t��J>���2C��N�/S���6: �Fž��c����ۿ�1Y�dL��Ǎ�Fn��{�~��3I3�����~4s�te�t��N���[oƭ�|�ʎvH��
%'C31�@R�@��#4���qP�2p�\P�-�4�3�T�(@��z|?PN,�f��APYz�̻te����=�y�)���� �d�ʸ钼b.��\���0 ������u�쵫 y���hU ��x�݁�߫!o4����t@��1v@��yRfT7\I#��?�(0>����v���g4�#�ۯϫH���:�!ȟs���ʯ/�J}��D�}�Q�&4����S�a ��(0P�8'Dz��K�N�S������7�ac�kr2U���M��B�!\OtD+�'�(���92��xuNk�A�@��di^��Y@1��G�*�&��e�5d�S%,��D���s4�����J��܇�D��y���M�����Eш�`,�d��ϑ�[ Y�y�9;$�Plߧd���0s�{�'P�z��"V��15���׶���>���W^�X1���Ә>t��%TfN Qj"٢�F[8ڍ*�e��ʋ�O}��|�~��������O��f�D��wގ_��wcl�<�����#>����XZ^m��O<��{�o��?�	\y�U��#�೟�,^پ+��5�j���?��n9n���ĥ'��}߰a�z�(O>:��$n��v�灟�کժ$=��G��7��NW_uν�\іFWM����L<���	�Y�J�lͧ��yf'��K�����4�1,,̡ߨ�]������IRڷ!Zѓ��ğ�ŗ��+��ɏK�V�"�c�C	S�
��O~��&�%�"-v�e�\�,�0^��r^p|Ȭ��V̄v[�ȕ��l��g�K������m�&�Zuʠ�M� 14���g�Cme�҂��v�$���%������m{��cOb�΃(��Dvl�U�왒.��g��h�!Ms�P�	G�����zp��>���Od�%ݻ0�����4� k��g�*��p�ƍ�2�����=J��8/4�Km�8��W4���R����T����Ҕ�O���ۯ��g>�3;�g�O��j@��/|����_��j'�9�j�(���^��^�l�챔�3�~������ll8W�s6Κ��Y��0��c�h
�\Z��&K���m`�t_��K���z�uh��$�:-��iЮ��0�|��L���6YPE���fO�C�Rs��߹�v���9V������2ҁ��" �9:V������R��0o�.���Ln��	<lr�c1��Rf(mS�P���byyI��f�9��U^^�ѣGU����f�ɚ�,�qm�;��S���>R�"6�s��0�RQ��l3sG�c׎�8qh?:���ǆM�AF�u� �����Pc9�e'	ތ���6И2нfɉQ\s���]�`!��ieJH��¡n8է"�˦3 ��:_9H,�(l��r����I�<�;�6����XB�CR�K��Zm�2��fU���?�A�Iy������V)Se󂊗�zB���G�P�C��ep�s�3IP����8�{@�����t�8m�k�E� v���e޼7@�$
�"����aC�1�5�Gʹ ������(EI���+
�e2(&↯�V1���O4C�A������B��&��ow�>5X:5p�Q���j�1��(���q��kX+[�4@�3��W�zj@��j�(�VU�����H��kũr�@%��8e��q`@`s�+�ޫcS#�L�����A`'*6�Cp�Lh�k5:7< �ߙ��9�<��l�!f��}���0���f�mmY`�ʳ���c� Fe����@M��p�y�KRD�����V�fѪ� ��a��8���Î�{U=�.���u�`��,i,٤�U��[n������+/F>C��£�{��7�=�����$�o܀�o�o���ذnV��ٗFi��cǎ)�$3�LJ&[�#X\���̌��;v�3��/��:�̳���_�2~����}&ɲ��4g[��<cyF���� �c�&Y��HqPae␉@j�s���"<R(���~7���2�����=�o|��׾�*\��K0�j�\^��Ջ��J!G`�N��jb�VA��D7��+;��G~�c�5 E���Q[:�{����D.M����N���g��M<��6��ZV:8?�.��8�x�����x�[n�!)�ʲ�TA)�1R,�ݭ�a��kC��������s��~�H�%=�� I�0���2�i,��JJB�j_}%9S���O�+䙡߫#�ĪH2��**�j���W���^܁t��$�0X�̤�S Z�F��KaJn�-�,2Y��K,d���"��i�q$ؐ�/������*�E��4/�	|O
6��W��L����g#�Jj���?�D1U�̿KL�^�~�'3�����>�[�ۮ������O5 ��_��m��Ͼ�߫�������Et�P�!�2 ��8�+�*E-[�/v�j
I$q֚���s��3N���ǑC#��X;��n"�F,�Cs����
����d� �U��vYv�/��� ��� ���уd3��i�F�)�q:�$bH�A30�1�W��!�[镁��5��R��Y�u繰:���k��o��r���D�Y	���H���P�::��s_�r�t�t$cciJ��_�W�13�߳R$f����N߂����<��΢��e~Dz�ˋK8�w?�Duz���k��C[�h��t �2C��@M��c����p4�Jŷ�N��x��A9$�
"��6���8<� $jhl��>_5������V��������FHPU��5��?��#i��.���U|�6�5Yʠ�������!��{�4�FA�'@����x�L�R���6nZ�oQv��sY��@�q
���A��5���Y?�ڽ�� (Z5��d0���K�Q�@�w��C��l�2d s��������W
N��H�p��-9}j�^��F�o4p����>5@8���!j�ʪ��#.���::_df�(��E�y?�E�	�i�)�a�f����������SA�n�}�g��e��2��������3�ȩ���3H�^�jw�<�ml#	�NV�@Pk�~����^���x���l�9�q���P��6�l��l6{�Ê%N�i�;� �ԜhuAUK�JUR">���o$&�d���6�ƥ�;��MbiyϽ�"���/���J���*��>R��f�H��@i�J#�$��v|����9�&n8���Wv����⩧_�=�4즛n�u�^���	�v�Ԩ�9�V73���14�5,/̣R)	̳y���4�;�|�=���>[�����������ܟ{�y{#~+'���)��s�&V.���l٢����Ǳ#3�t{z���~��~��{�������'�͇���٣���p�%a5��2��!�}�aO�,�f���[��M��m��`�+�Qa��0&@�����#�p㕯�o��b���{:�_�q_�ƣx~�~L�߂M�O7�g����,����߀���Ez��Ѩ��s�N�ܵ[~���}�}�/����D�A ߗ�f�F�\S�Ne������?L^��������Yk��i��D�K+JQ���hk֌�-��%�b�V	�^xa����aǮr�m1�O���W��=DK�cC�O_�$:!1L���/'TBZ�>���j�@�/Ic��9ؘL|H*�Щ����Y%E�>�{M��z*�Z�%H5�A8�ҴlIc�R���elX����o��c����v����5?Հ���������x��k�����-�p�xqvM��S��^t�we�F��FS�\v�x�-w଍�@��L���C����d�^{f���ן��?���$�����]�ͥ�Z<�m[��c���"� D�%�f_Bْ���Є��o@�2~��!�H); �0�c _.��;���3C�AzƸ��`��V"d9���.ҬC-��O�]sP��շ�Х�k����!���@@�2T�2E�t^�i쌳����s�����ѥ,�$�h�Z��w@��ʡ=��,H�Q��9[u%��+�
�"�H�Ǒn�$�7��w݁�'�u��.�j�sީ�{���c�C]+�Ԩ��+Þ
f"d�R7ڇ2�p빆��3�
�(7�  ��;�!
�¢��0MRM�����@�����4ό(xd@�>�< pz��U�+'N)jQ���6��s�nr���Q0����K̖m5�|n>���xM:=��(�M��Yց��7|��/�JD��6^��u�o�ωr�}O
���澃]+��~O��;h�&��(��o��`�5�c�:"��@��U�h0��g�i�T=-rW&:����`�1�r|?�fW]������Զ��zF��دك�`�5x��0�����O}>����ܪs�U"(��``�r�.��M��R1:�+`��f0H� �`?T'}.�\�3����{�|�_��<��~���  ��+���雯Y���g�7M�ȍ�ڦ�����i	�,p�y[�n�(N�ž}{D� (�Ek��kH�Sȧr3��Z�t    IDAT� �W�vr���{��<�͛֠Q[�<{��}������S��x�&�q�m����5����@i�a�RT2%������L2!v��4f�u��� �?�B�#����{��ź�p뭷J�����ضm�*�sn���q�
��ä���C(���7��Գp� }�Q��}� �Haw�}7��]8�s�4���g���������w7nZ���:��1t	4��1)�P���X =zz���v�s�B'WDfbR�k��,�O�������p��	5p�Zm<���x�k���
�cSX�q������+�X�=��.9z�;0UL!'� )@ֿ��3�<�/~�a<���ba\q�e�*󋀟ϙ��O��I.k=��{��߾�Y"ǒR���u���F�䛰ē�<�V�����j8���x�}w��ֳ.-�E����K���<�;��!�#�x"-�F�&cY]dRMUaJʃ)i�(���Ͷ�_���L
�d6�'e<�,165E�3�juT�a%3�U�|"ڣ'D?�$��3�>2�d�Z��:�]3ɪ>q��b�T�{��y�����b�����������?�dV�]�MFZT�P@@�8�G�H�bH�M;t�%el�"�,U���D��y6�{�}�`˨�&��&�9;HX����(�c�9]�C_}Om;&���Ȅ@�D.�3�F�_>�g��U���P?��<F�A�;P',�o ��ތ��{�TB�fǔ 0�Ճ�5'4f�c��.��	`�z|��\��('�2������N�XS�M,������� ���T1��A�Ar��1��͸���q��߈݇���)��l�f�1�� �oͣ�U��i6s|��7ʋ}ȸ�L2Aڇ^EP:P�1�:���T�bt�Z9_���<qL	�ȫ-A�;�3�����A�]Sh>#���L�� R����,��@M�Cv 2X�sH�zP0��ٚ�]�}��8�Ual����$y]!S�xs|4�6u�-dQ}����>�� U�@$B�1'�a��d-$�Dk�fzO��CE�(�q�س�|��=�qp����D�c�C*հ������q�P��"��r9�A3�Шˁ�_�v��<�*#���f����=(����Ų�C�S����� �:�'��̫a�8�X0�C��l�R��v~]���x����P�T��*��k�g{�'<�����R݆{�p^�ar��3>X�S�!��̽χ@�q�Qh����2�2�҇�������>��5����)(N�C�P�փj�N��q"PH����)z���(�\�9����>zᔀni���%���,�K}���Z���rh�*�B!C�_*G5Р�L������߆�gp�����Xc�ϼ���~[�D"�ӷl��o�7�|��b���۷++K��z�tZ�f�#9�����;3s���R��C����zTjU|��_����.�M�6�n��wީg�}�>��>���s�߇N��1�x�����O�Qk��nP��Aݭ���#��DPx��W����4Z����x��#�
I�@8�Mg���5���Q��$R�2��肜F;�Fi�Y�������}�gދ��Q]^Be7\r~��������(5[��_���=�^B'Y@:�S���Rr�{�E�v��/>�^�M �i!�ëx���?ܪ���uk%��*��,-
�z���F�$r�5�ù���������sa�@�b�#V��F'0�&�5�3Pe@������b�������y����\�blt�y�%|����g�َv�=�Eyh0@pO��{3��>AsGa�OA{��w��GTF� Y�CI6 �G'�Gn�&7nD'������5���Ń^�G��b��UM��k�*����=�k�	u��HJ�l�T��Z��������k����������Z!��?�ʻ���_�#�W�[�uNN��Rn���<zq��1��I$�%�֑��q��V��L?�D���#cxÅ��;���7�6u��@&c�G��N,�Z?��;��W���W����Bnb�ZW���i$�X�8�~�˘��,ОE<a����h02 ?�[w�@��3���X2���٬�P~�9 ��+Yv�XDS���#Enz�ܒ�c���5� �@f��>�N�Z@�_V�7#_��$�5�l�D$��T2�"��32���|&n���;�B�6}L:��zWҩ#�"f�ƞ�_@{��1�RU]8�e e�  ( ��x&ۮ��:J~���DM6��ȯ���܀7��V,�ۘY��l��?Z����+�^��$�7 Y���V��X� �@���h`ͫC?�( s�t*����!�j��s, P�},�d� ��B��%|�(4,�FmJ*2CB�fꐣ(�3�N4hg�������A��ݰ�ҞϏ�`B���*<�ςF��z<��`G��eC=H���{*�gN|z&I��H� ��v���O���p��P˟E�~���:\�3:tQP��G�<�9����ީ�= �A}'��>�B����D�B��d��5��|9�3��r��,�;Ѡ����cjOC#?�N��z��v���U3�D�<�(ষKt�G�D� �7'm�<�T��u}R�	}8�Ӈl^���S�����y��(��&L���Y3�)v	�g��7Wp�IR����oŀ�j���eu:z�C����i�
	��d�d��*�������s�����2���Ld�oT����8s}I�6ԗס1����ӋI�������2����|�C?�׽�l�����O��O��o��Kg���M7݄t.+jΎ�v�q�X�cRY�"Z�:F�yL�E����٣ؾ������>���{1�<��~���Cj<f� �D��G��׿�������ʆ?��������C�j��׽�BI�~经((au`|b��{/.��lݺ���K�teig�}>��K\��+1�Mb�3OcǓO"Ѩ#�
�X�y2cy$ٷ��{.)2�4'�JS�&�^��r/����S��ӻ�a���Ǚ��N�^w]s9>���cj$�t,��fS����l}~R�	ĲY�Z�u)��c-��|+>���ጩ�<Z;<x�������C�I�݄hT��F�����U_��J����TVA ��q:����)|�Fq�6>�j�� X����ZKKh4˸�����1\x�vf%Rx�����|�4�1d�􇠐��2��M%�e2'���Q݉XM��K��\��1����8�6��������g3X�k4{xz�)ٞB1�U@@�$bVU��+��� ���įg0A)}:=s�m��~"�����c��*��W��������ȯZ#6N��B,͛1��d7�d;����5��]�Ѩ.����N���#���+��{ގ�]�3�Iv��s.Ymm�1R9�����ކǞ;�fb��I�i���҈�g�����kO�@��d�"=r��Z�V:2��J����C��G�c�gSoD��E(�{m�J>޻�	����%(eH�P��>�t;�NV��I����Б�d@a�;�&���nh��� ������p���̎�.��o~;�S���14{��N�Yk#�Ob����
�l@j3jg�BG��F�(��}Eb58i�ׁ�������U�^�����+n���|�YgQ�,�vW`�,��}�T7 �Ҏ�6�5{,Ȱ��x��2�N* e��P.�S�V� ���#Vg�	��ß���U$(w�ʎ�T�O��D���cm���H�|�~iJʒv�5�7��f\j<��|�!�Mm<f� e 6O�]t}�9<>|xP=|���@l Lp����3`95X��d@�2��#���F�՝\�����:Z0O��]!�<8P\[h��VB���i4x�=G?o0�O1�6�?j�\�d���Y��Pɇ�K@ƿ�L�����ѨL�`lN�/E+7�����{�0��+K|=f(V��33�Qےc�Y��qp&�L��Lx�3��t�����q�̒�d1c�J*��ӽ�[����U���t:��O�
�w�^{-��������]#�Ҩ"�3H�̪~jj�>��zUЮ�4X8j'�25.�JVX@�	>O7:��)n��� ]A����[�;R'8^r��T�Uh-ZȀ���W��|�`�N�ҟG��P,Wq���\�z���u��)Ṣ���d�9��_U2����EN�.Q�U��\S��Z�޻��W1z�Gd!�WEl���}Uj��-����a�d�������	�t�|TJy��܀���	'�{ל�s���9�H��k�nt��#A$��T�l �N��%�h8  �(��?Ћ�;�������k�b<=.�G{===�D�׾�5,^�X�¯~�+����_�"�;�8��������_$��+V�����[���Ѓ�n݊Gz��vJ�d�����?a������FT�i���(9aVx�x�MR%�x��â��^2��p�qo�]�;�a����^�K����u�����.����`֤���+7�A �
O8��"�{�Tp�-Kq�mK��T+d����bՆH�3�`�<b����� �=W"��r�פ�ڥ�ւ��|���L&EU�!���"?���k�����l��@�r��	Dc!,^r)l�P�x�o޺|�q���*�������Kv����d �s� �hT�^��]���Lܫdo��H�xc��
��*���h�<��68=Ke��'ஹ�Y��6zZxi�V��А�Q��C���[j��y������NJ�k��V�娿����\����s�~��}�W����n��3/��+�����i��\)'%�/�2�Q�F!/0�4�u�ȍ����D�\x��Xv��8��)Bw:9�������ۋ��*i+�X} yW3�Q6���wU�����+@` Uh�R%�GF���V���SM@j�-I9�l/�&��d��c��v�QYm�UL��d\ܔ��r3��]Ӻ�: ��`�������A��,IP�4)�QPj4��!3�J�RY�k��
�5o�f/�9��@���:2���ɷ+Q,<x=�w�<6���=���P@��S��K��-�𡀠�I�M�T��8����8g�G1R)�o|�^r�`��κ��__���m���ޘ�Ӂ/��)`U���j��'P�CY�͋v:H%ʪpX�E� L�O]c�+U�(\(5(�3�))熋�Z|r-��R=J�}}I��W�%��AޤZ�n�|�Fŀ���N��+��t���fإ��5Vp�*Qz�KY�J������P���<�:x���d��b��|X�h+ A��E���{t0Ը6 ��{p��[�Ff�O�� :��k�)c|�M��'�@&�{�;1�n]��c/@��l��<4�k�wx��
��@_o]������i�_��J���� X���."=�d�mFc��?���'��_'��z�B˞ښ��c-9_+��xu�������ӨR��(J��5�H7^�5�����\v@ '��3�iY%:N�ǩqm �v5�կ���l�u}��n9������y�<$�U*�P>A�w��Ê'����]�������\��+�-�;R�aҧ�jW,�������.����8�ϟ!��|�5�7�'?�� �b����sp��c�W�unڴ[�o@��@�P�����p$���(�(16���^�4�qߧ����\�t>�g�}<���k ��o|Cz	,<� �����z*~�_`�Ν��cWJ���^��M��6�1"p��Ǯ��o���}N�H��L�6�����K.z�xzw��009A>��X&���Pe'�o�y�ۭ�G�~S�>[`ˁ^��Ѕ������ħ�#�A�Z���NÏ�~/BL`:�(V��[����=�������U��������.�Zb�3I�Y��?�4v���{7�i��T�������z=�I�ȿ�
���TH��d���ߺ����W�8�:�����p	��N,��r�t�M�:m� ���y�������|�U���R���%�g|}6���Y��Ĭ�QOȩ`E12h�V�(�!��j\����55���"�/�wL  ���O�F��U�Y��V	����"�XƤ\��ZH�3eP�jI�҅�0s	c����nX���|避؞�W���'ox��Q��)�U��Q,唙�u�~	:�.?���,�.��ƙ�,��o�����Ͼ��z��fܴ�:�y�	E����6f"D����@?���> �߁`�$x|�*��LTG���1е0��j
^3@t�k����Yge�1��h�i��q��R��8���	�l�l���t(�-�|���RK�D���
��Ck�.9�+e�d����b�%�*�j�%����"�d3�� Ȭ���{/jUf�0��'M��-��S�E��(��2�57<Uj�
�{п��p?PʢZai������}@ͷFFU�<�B`s��f�PY8nf��&�}٥bL6\�c_o�,`v��cQ�dY�2��iJ����jʑ��j-�a��4�lxSp�r+5�b(S�x8,Q�(��"b���]�|��;8͍BaQ�S6�{��E�M�C0���(Lѱ�(1F7MQȨ2��+Y��)��x�񘌍Ȳr<,�7�f���
f%��Z��J�˪ZsG^��1+��փ�������4��h�����B ��j�Q�xk�}퍀ٚ?�JX�9z�����U��D����������=�����q(5��9�Ϩ?���֞��_O�c�ԃ�z���~]-��'ip��Ms��[�Z8'8���l5��e�Ys����كi;�Ҵ<i@�9>�"V����6`��]�ܒ�U�~��9$�y��A+��ԥ��`X�[{@>�����?D']W��ϊ��%GZ�~��2&�S��� E��,�:���fz���ԥRQ����R>g'3fb�}��v!��'��i�$���?��
E��Ѓ���QB4���g?��fu�E�
8�z��: `r��s2���j\t�G�Eq��A᷏���μ2�T�C�nʚ�rH%ƑI'1�Ak<��}������eĘ���;<xPѿ�n|��O�ꫯ�[��!�a��?�y�~�i��~����ᮻ���)���/HǊ4����J���.|��JɀS1��	���q�E���`|�z��@��)��e�N���w�z������_��C(:C�NcKW/��;�!�����#���(�#g�����/��>Nd��f~��3�`c�Tl|�y�A|l��Rˮ�_��.�3�ٹ��>���%�񩠟 ����cLDi0�ְ�����/ �� g�%.�J��I�]Ȓ~�X�\yv�K���4*Il�Fc`tlC���5Eq�����n�/���_X��>:N�vQ)��U�7��䭗�¦)�A#�DJ��D�uR�]K¨vT�v�ܤ��u������� i?<�)s��Q3�(�0R��}2&��uIs��,��, Q2c��A�!�RY��Ҝ�-+n����|w�G��>���?�� A�Vs�����7V��g'y|�CQ�����Xn_�P\$/K���*:[��?��]��ډ�^�=���E^�s�>nO�	�jSE�7ǃ\�����6�5�@t�m�u��7\+�[H�k�k�۵0��d�vS�F����[<v+X��͍�j��MqCU�j0��Bu�ˡ#\�n�$�޿��ZN�܀ٻ,w��O����>,�e^*�=>�k&}�45^���X}��ұd�9�ep�PU�
U63��Pv"�6�^�ϸ =c)�$�֜����?��{Q� A� �, i���I�����{4�Ҋ;XEa�������«c��a�Cp[Mu,9K���"�@��	7$]W�؍C��oVah�N Ţ@0��~U5{K#�ڨ�Z�`M�(Z���a%�h�F� ��}�V9UKd�t9��P(�I�Df    IDAT�����z�Nd3���!�~�wO�� �5R�y�(�k�7�W:�E"�B�U�	ʫRM��V1kX���X��=8�gz�j��[�q�s�r����1�;���W|�H ���{@�N��uP��5���A�$�@U��s#���^{�� ��@�׫	{ n_�����?ĩX���'�����/���0�wZo���+-|U�8X���qB���fl+)R�UUm�	�|2�Vf����*�!���@�}��sU�_�q�ԁ�'�C�-j�l綀_z���P��*����x��ړ�E�.K.���]>'=a�>d(�&��#� �ڣ��5��@ɾ���\�CQ
u5�TF���h��*A�Z�@4�G��,��0�������2p�3}.="J4'̞��p�x����"
J&�F	꺻ੰ��D���γ�|��7]>}�-؟��٪6�{��6o�-�Y4ބ��='�r2::'I¤����I�����8.�!`��b>�B.���~�~|�_�m�nA&��O<����[��*���=��ƫ������{���`������?��N<E ��W����ҥK�5^ye�z�-�����M�$���?�1.8�\8k�ݍm���,a��$S�H����� )"f�N��"��/ol�%'�ŪM]�O�P�z����fQ�&�����ӿ�Z�!E�\���l�o|�v@ �5NRZ=H�F�p�W�s��/�8�s֬|�w�s�*��ʦ4�O��9�󌒡�՛f-�^�Y%�a�����)�����x<���ף̹�$IfQ�t���( ̴S��R-a��.��������;k�n��o�޾ax�ax=a��&�$J�ʭ�C�ٌT���|m&Ԍ2���E��JY�+��ǂ"[����O(��ˇb�	�/'�_�PLOG��(R�#��M4�(��L���h��y�,*m��/J��Q����ӘN͉���������+�]�7^ٷ���G޼��U�E:N<nfN�@G<��#G�f�&���C0ގ`s̪R_�|���h��pڱs���+����ޝ�E�w��yp{x�J�qp3��4sD�:0^p��]xm�TB�j� >��(Ù����qd�@qHz�Ϊ��۠��;����!�(M�ϭ,�ެE\h
00BR�R�ꐘPn�9�*	o�����i%��fXI��5�������O�TFu���C,��\d�6�*�#t�-W�(�0�"��+Nۦ��EK0���e��I�_�B��1����^���
=*��eH�ҢB|8 �@�?f�(C�6s�������A�� j��fa��Z�@��2հ�SYt�=X��x����Q�KƝz�4na���q)�9q���HT�g�^5�|�f�Q���9:��k�ӓ�X.#�ɠd$����)�*7BQ�`��ʬNΨ�����21�d����L���`t,�\� 1��73 ��'�,k�'˔���@'�����������u�&A��a�����gR��T��%��ց��\�k�_
,��2���	���; п�kک$�5[7�kd�u���uMg����RY6@Ŀ�4�~�r��P���������_g����@L�^��4�H:8�����o�@�xJ��
���\�ʺ�Z�F�%f
?����B�]7�|nT*��eF�� k�6�,t
H����jݙ2���S�M��phpD�#~�:�1�kTӃ���ާ�X����O���3K9A+���j씲����J�ݿ��fS�\��;�{��y6�UʤY�~.'{�hԙK!�sbfG3zvm�;/��R:���	�)�i�����V� ��f ��H�\ɦ{p��%H����^�f� 6�kio�9瞋�O;U�ž�~��Cɴd���cB��B>�Z��������� B~7���/��;nE�P@��?>(�|f�ٰJE!��Ħb��g>��s�Y��O�m[�J/�H�='0����q���Ϗ>���$DBQ���1Q���~�s�:S��=;v�������~�%ǐȤ���2�]vB!�97ʦ4��H/Gk�O���,}��8C�NGP,��2Xr�����,���L�xk=����iW�M�t�Da���иo��j�{��?���~ ���QI�Q��lio�`�
JvY�I�&	0H&SG�x�5%=/����Z���I��V%��%+��t�kX<Xݲ(�����SV�Y�Y��s�4$SY�B2����W*=J�z�+fQf�i"��6�������rtKvx���Au�LN������<�n7|��V���n?��fF���F�v���$�N��l��"�&�r�Y�
�8]�`�Y�I��@`%�+%T�bg���;�^���q�A�������*o���ɧ�}o���O�:e�ҫ.�9�����#��x��W��K�a$k"��	_�N���t��ᦏ]��O>A���n�X��υH$$��	����i�T��(^z��W�E��O�^�M��P��al{o9l~W��U3�Q��^�ֿ���dL,@�!J<�T�]p�C����`�����2C�HE%C��{��'�������$�l�ڈ�"���鑅��H,�q��ʬ52y�uZ�D�-�e^��U�N&\0��iL�r��s�iM�+��	w�g,Z��g���\	�C	Y1�v�U���ې:r ������O�)�����k?`��Ԇ&R�8���@���RC��ٸ��+p�%��pz�^�ʎi� �iK6��u��i� ��l�ͤq��"҂X�Q41f�yؕ�m]���u"���Sc@�I��r82�GWSf%x����"�OQzJ�7*������P��@�IFܡ�M[Ϋ9�U�J�T����8� @�	��	I�t##cU�bYmX�>0б4�	
���%Z7�����_C�@rBSl=Pѽ2��A�~}�l:(�5��ve|� K��`\*D��^Y|إV�"��NS+��E=X�SI{f]��6@�_S�7);���ؒ�����v�Q}p��������0����-�Dm�:;��]�� {Q�^ �F��Q�T�t2�}S��
�
x�I��9 {�~���[��AA}|m=/���ڡXUt�c��V�'�Ru�c��T��Y}V^�)IP��$`j�����؛�uŉAw}��rҶ�����7���+@ ���\˸[�
\'�[��&]!_,�k�����
���R9�������s��6D��صqV��U�@K[��f��,+e@�b>�a��� G16����8|�7c�����y97n؎��a��D�b�ٸ�+p'bd|Lh>�Cê����O�+��hXV��J�A:���� �c�s�(�=��3Bb�����Y�믿^�~��Ș}�K_��\( a��}���K����}� ��;＃-[�Icm&��ף��	'�����I'/g��[��Ï`����Lb\��Ц�f��O�4Ebf�墘��q4w�Ĕi��:�ؓ/��U��|g$*��ύ��_��v��J���������G�����ʣ�L)O#�֖ ��Z,Y|���`ӆ�8rp?��	�Vz��?�뢚�CZ��129�Ƿ�G�=�	IVx�-� ������r�հ���auB*%5�L�[�:>�R��|IL�(��~��Q�Q�	%�Ru��c�
��Y��ǃc������>�T���Wr�"�C��~&}�(���]1ӈD�h��.�d�be����H<Uf`ON���IB:��=�t^�,F�*=�T���fe��.6���誰�{h&Y�����m�_����rɡ�������翽�`��ϼ��u��|f����Z�g/섗m�`��#x���x��5�𶰑�}���_�#���S��ߝ>N�7c#9$F�Q!�M@���d��)�%"��mƋo��+�u��i�/��ׅ�p�t�-�c��+p`�{�����*c25�U�r+N+7V�|��v�ߑ)^w�e������o�f4�N(�����UF�jF4+2ai�!lf 5��jb�����L��+��L�>5��C@�� �ڞA��:$xh�,]~�x8I}p{"˚���p�Gc�	�b�TA�H�q��cGz�g�z����:�Q���/��L�9ĭ�hq�~>^�ਚ��sJ%�3�oX�c/8�G1�O�Iy��H2u6@ wͪ��hP��M��ۉB>�1N�ba��Q���ϋ&�4�QA����:puÔ� lim�8M����L+J�HX��,�$�A�BU`��h��l�"1�п�eNQ{����/�	|.��.:C��=����a<��Y
7U�3�l��:`T�dQ)�/��Fy�e��IO�ζ���ؿ�2��^C*�Q҇�����C���xu0�0�A���u��R�d�G+��}M�D�T��mu���C]�=��t[����?�y���~,����d?|�ﭯ��]�1���"�kBe^Z@Z��x�J7dn��^�p�5�y��Yb�C`4 ���r̭_UŬy��cC=o��n͟��C} ��n.�Y�w��w���Pn�j���-I�?�e─�k��P�!���%趚�� �~�4���bq�sR��b�I�QsX�U:A��b¡PR���r���U>�T�t�@�a�>��T�h���`צ�X����pҸ�aɘ���V /+�Lʹ�jʹ�����7.��_��s�
e�{�ͻ����ﾷZ�=�Y�P��d��Kf<�h��J�⪋n��~J��Q*d�}���тo~�����[�
��/��_�R����s?s�g����_��ג����{�t�� F�G0}�4�ٻWn�L��o�Q��h�@���;�m�����:?��O�p�B�6oX��<� vlۂh8�`$��i _*� 	��i�%�TvT���BЍpS+:&�@g�10�n<��r���:�er�����޻o§��Șe������g�޺]p�C2ߙ�b���]ÔIq�p��wL'܉m�ס��!�p������$1F0���<aҋ�#�y�*괽z,�y<�ċՁ���Jn�sK�N�1�C'�����v��B9G��ߏl�pxι�aQ�48�I]*�P)1{��q��8����IY������Y�Q�{���#�(�N����p�[Q���c7���/�k�?�r�t/�kR.���s���cf �ǻo������R#�"�I2I(�"=���T�#���L'�g�?}�͋��ͫ.8��9?>��
���G��?~}���?餓&}�֥8n�4��GJ���=C������]B-��QǸZF�WFGS �[#8���p�E�%BϐڨPE �c����P���A��E^<�����TB���uH��z����k��{��8��} ӯ�Ni�W%��,��Z�Q�����+����,lцt����X\up2�X��1�:_NX6�����a]l&�ld��\�L2�&Q<�j��4��c
��4�t#}EQx��"�E��a+�]�d ��uP�߇@�	Y�	_Kλ�*�Ι�d���q.�b��pa�o��|�ܡ����D�ʋ���?+A#0PJHbe�Z�?�@��y��0/�<{6���F�p�Y�=x�R�sK���&Hj�x��r�HM������(_+��
�
\�T�v�L���>tv�#�Ju �UyQ����O�����ٜ4R�Q*�����8F��DLwLVg����H&�+d�lnmJ�E�.(�l*��`PʋMC���� Z�!�7�X�����*/ Q����ټ��M�p�/�\�2���|e�@WQ��ݟ6�B��VO��u&��_F�̬����������ZʖA�q���� �*�%�81h�5J���j�r� ����:e�[��4`�r~s�Y���v0���b\(n�<dT��末D��۳=P�`V(� 3�{�Ħ��:3��ف�=p�vB�+��"����5�~�a�,�}ph5�r���F�7UD��}:�mץ �RR��zgl��-M閷�����P��	r�j26�*���%_k��=�A�
���ʒ6#�f/�Mq�I7\�L��w��2�5/���#U���h�Q=�u�w" ��%Vy�{<��u�=e����5,>���r��T�.c;�+Wv����3�a鱂Y@{S�7��lĚ��B!�<n��@R!��v�^6�^ǆ��p��W��eWa�V	�X9ٺe7��?��W����9s�aѢE8��p��A���!��	��X2��e��l�cE�	&�JH'�̩�����m�n`������glݾ]UYP����.�{v��K/�$Ypҁ��n���U��ob�ʕx�wd��OA$��0:<�U�Vᙧ�@��z�g�'?�	N:�$��|�������P7���e<H��2�pϘ:M�T.rF���D[:Q��1:X��o�ƁC}�DH�,#�M`ʤ|�s���[���m��pa<_��o����}�v+sS�M!�W賊��(.��"����o�6l۴���ړ�M�4V�MQL�2Y��6�2��h�ƵL@ �SK�G�ΐ��j�[�J(���b��E�X�*��$˔��H{�z���*�s�J"��{P��T,��Dt�dT���+���罠x}jd��L�7��5,��b�"4~�l"\��xg�&<��cش��
��5�ri�
c�����/��>'�\��=���Y�5��|�K� �ES؋�o���l2y<���b�F��J@��x�%�I)j��H#9����~�*j�Lv������oc��D����" �����-������={f�e矅k/�Ӣ^���\e�7m�����AlܸcT�-��!q#�ᄉc���������Y��1�0�����Ǡ��B�@���ӯ��K�m��k�?�*��s �
ý8�s=ƺw �>��WL�(r�<Y\'*���S&���T�|d���/:�	Dn���I	�F ��!?���E.9LQ�	�AO36	2�N-z6��#��	���h�A�2/|tC��&�����G���������Ç�#T "G�A&V@(��׃`�+�,G�H��xq4O��ؔiwLA��Gɬ��v�Q͗л��{� �{ ����@@�t9l:���kT�le���SYMa��1�cٔ)�J��L��Spŝ7��Aw�$i�}*�^�I�l�)<�Z���G������!&�0�py�k&���!����"�<u
�Ѩ�:�BI� _��R�P�dJ>B㠜�2+  Hԥ^��2��\R%b�����}��i�����rFYއ �j{s��C�M�(p��cQi����S��G%>7_�K�����>�"\�LT.a�@�@�G**8�B�E	�SΖ�:խ� X+0IK�=���FQ�ӲiVvH{R�]%+N�t��������dS'���
+ ew��)�T/J�Y�ESat����t6!�{��=��a�r��-�L��$�N�:3S�����u�1����| ��)�O����y�d�P���A������� �hjV�e|�A���s�LY�?Ng�c��ov�%����:�ASU&��y	֩OoZ�գd���
٠�	-����x*K���̲��c�iM��2��OUV��RU��c�� 5���DSo�s�@�+��d�**�Ȋ�{�
�)���4�s�a���h��� �G�r>��-4 � J��TG/�*5�O��i@���h�[�M�����T���~�̬��g��XUD[u[^ס��u�SVBK?>���O h	���b��Uز~��4�T���Gw]1y����uLz{���%G�Ĩ�wވ�^�Y3;P6iz	t�9�o����2�ך�`>ο�"�I�Sғ��g�x*��є4}R�M� ��YܫG�N�a��)��׾�믻J����xC*]���՗��gs.���� FGǥ�{��c�,��?R8    IDAT�d
��Gp��>I ����Ta*T�IIա��e��y���_�+wܱr�����~���A	�3�������mm�2��p�\Z�^sG'�&�B2]���7bժ-�+���;2:���Zq�7�s��>WY��C�4{j|�%t���A���`�, ��i�/Fq�֮Dz|D�P�$���,	�|6#�8h��0� �i�h�J+ܬ>ə/g�j\f�KW�<T�s*+=�8��t"-��b|�
�����˓j�
!�X�I�!Ǚd�"Y.x��*�kJ�`V\F�d��5��x]�I'���K.���^�����d2a�7���݇���/b�Ɲu��B>����� #@ܿK��?�1|A�{h/��6^[�c9� J�fjUMA��e��ꏜG���{ϯxEx���\0.ʗ�DR���c^��C�q�1�>7��3��2���|���>�_��ܾ���J��W�Ҷ���z��n��鎶����8�/�;̛�	#�G�d ��a�}��]��7lŶ��H�5x�A��B(�y�B~�}�	�����`�L	��팄|�9g�Y1��b8��M��ċ��Φ��6M�7�*�-l�:�{7�F���H�'��|6�r�D9� g�/A$߁D*�Zh!kM\f;t6(�ǂ�HX�`\x�Y6�
��?J���M�Ur�<homF8LC ����B��D*�#��K���A�+(kNx��ʀQ�`�������S����`�����l��e�O�7�D���^��5�c�bF��; ��1�̠���C�D%�q�C����� �\<�7���X��hu�s�<��_�J�I���Í�I��W�%�0�C��ȍ��U�Ŕ��A�	� 
yVR ���U,�H͔9@���0i��l���5��hT�.�,�@G�I����
E�ۨ`����Ȱ4�
@c����}<\yH0���t�=�0�wQ7�5��S]e�U"�9�l`��HY�AVJ8GZ��:��-͒�Q���Q�"���àU�r&<�vdK����oh��|n8�
璃@WU�$ش���Kc��-Ҍ�z&��8:*z(�[6D˚fh� f��M�0�̡�*��	5�O�>�&7� �@2A*h�3�" �T {�V�:�b���%;�T��h�V�v�&LD�6@��'J�U�
��<�̸ζs>�y��&ݖt�r��(~l�&{�(T���Fs��q&�8'��M����С��G�_�~��[�g�嵺�l 4�Wu!Z���_a�M"Г�](��K��WX�6�"�W���`g@ =>N��֐���r.�G�,��~Z*%s(FGl�'��`��E���G��@ $f��Z.�ټ2c0�c%��t��N�)n����э�Z*Hϖ�5�f�Жs��O�y���>얊�	h�9�[�(2}�X�����M#�sP5K*o,��^�ω��^����G���^��hP�t�����L��Z�׍��Fiz&��E�YC�߅�[�c��u($Bq������T��)���2EU)��ZEzlM!�g�І�Om�(����[���[wx��y��q�1�e��9�-�� �I����bT&��l�d?�����6�����ŗ�Bѳ�?��_|c��r�/��Ĺ�Ԙ�BU���7��*s�!

�<16�b6�ϏX�>����grg���c�ꚫ0k�ll۶���a={�A���{JR��`9bʤQ��Z�v�x3��Y�@�o���>��\Q A�QC��Cs$�O|�&|峷��)�{ ��CO��|��FU��k�J�ժ���8�Dg׎-B���#?��ah�&�sR�L4�JonRB&^U�֪WL���d�%�H���R{���(煇I&H&�]Nr)IeE�����@���^�}E�n7L�zz�HU$�y�၃��e�M��f儙Ϣ���������߰��"[�b݆-X�v���H�
Ҕ�$A.�@����k�����O%��f��}x��7����0�Ax|MR���;�ُ�o�7/:բ��V��'_zc����6w�� 92"qלAIx�r�ʥ�k��@�D13�_0���;���;�Xz��N��=������]��s�����ⶥW��y�н6mێ�6�z��h�x�+�����k��s/bϑÈNj�ɯ���%Kp�i���)W�D,PZ�LDs�xQr��Փ�CϬņ=ÈN] w�YJ<:;\H��o�6TJ	̝Վ��?F��=G��uHʌ�XӦMA{{����z180,��֖v�����U�RGGN8q>�%�ɗ������=`��Nʓ��/����Tu.�f���-tV�RyZ�S�V�u�
�"kGQ���L�ç��8Q���g�w�\�_d.+
�x�U_�C�bf#
���Ș�dS�?��7<���Ad��s2;�Gs�A�#���g�6���i�CP�|( ���
��m֔��|JXV�u��-�pf��_�@hRθ�b\r�Ȗr��h�mwW���Яh�]u�Y��k�#@��`�R-	��ZGK�ڛ��-B$�Rp&W���|�9<(U*��@>�� �ĝ�� <�@��2��8f�ع���M�����l�w��b�TJ���A9 ����V�^UWl��V �9���Y*
�i����$������)�V�` �M���s��7B �MH����GG�L�EQ���( ��@����H�_]*W�Ge�"jR)�&���T���(eR8v�\̝9>���y������s�A�^��M���Q!)�K*�B���:��j޶g.e��������!Ki����Q���с���3h �Fϑ!�z����������U�;B����I���/��9�`ZsK=�1��R%�5���Ё~��c�Y��h��r�x��6��upi��`?'�VYq��ȰA���2xƩ�aHRE�)ܒ=�������g�ܩ������2��I��G���h8�p���U	u�_�����{R�����qH��Ũ�_��P-���U�dg1L�*?�
2�ŵ���(�|I}֪���a��*	��A>�JB(�.V���^����c�e���cI���������ڿׁ�}=�^�S�)�т������+ȭ�|�Y��UA��ܸ��mB��G�RQ��)��Y��\N��>x����YC:1�X��O�{��r&O���H�)����?b���ȗJ�T|�e8��D��k�.tuu�Jl�t�z{�eO���j�lp�`<1,����׾�E\z�Eb<��_�۶퐽�|}q����J�󜷸쬈*�,�����228$��'���C�&FG�Q�����ԩ�q�u���%�1::�z/��\^���E�(9^�`D�\.� m(��1�N�ǝz&Zۧṧ_���(̊Mmm�SծT@<��=w݌��w'���3�L�Ǘ������Ҥ픀�r�wV��ڄ�J�P�^��]5$�b�%U�{L�X�l�N�v-�����Y�0�6��B:Q>]�}��)�E㴢���^��!�HL��:ax*9�֦8T���9��+�e�9X�0�1���1�) ���0�� ��I�
"� ���;��1/~��o���?���0�<���8xh7I��}{�l��^�p�b����� �S��������/aWW?��XK�a��8��*ܾ�BT�V���,#�
z�Sp�È4����e?#�Ҁ�����>��5T�<������-O�v��������~�@�_^~�;k7|���t��`.�Yv#N�?�֮��>-h�K��.D{P1N��X�n=Vnڊ-{�c[ݗ�D��f�,��%X0}
��,�!?*EEGa�U� <��y���Uشo�����!���qM7�����&?,���s���ְy���׋H�E�,��0�шL��	�(�G�/1����|.#�Ķ�	�X���o�;�~����0C��**I�0|��8��X�����'�[��y�jE�јEc&�	&\x�%/d�L�������f�l�I7G^/�3o�Xp�OJI�����\�}^W �p�`X�p3%Yf�ܼ��7�� |l(����{0�{��0@�Q+؞X!�� ��:�WŪ��Nv�Hy����W�D��'_z�Tr��\X�!`ҁ��QVL�f	����P���L]�!j
�XΚ>3:ڥI�%���C=6yU04<���Q�,�pL��l���k����	U��Ě�̱J���J9@e�j�LOdL�JTV�(	(��dd,�< �$����sf;�
�3A):�Z1s�T�#aQ8��3g]�4���������T�"���Ho?zz��&h�Qq˫lӅE�#��R�� 5��
x��dl*��id�%G�������!t1�,��pρ�\���#�;_(*
؊��/�2�/��ɸY��:���k�q��	 �/�jR�L�jq�R%I(��)z�|�V�Ipf��
��z�ϪQ]e{EfN���s�L�dS��Twx�%�縋���~yH:+j?Pcbʚ�w�ĥ�g�4#�':��A�4���@I�@pV	E�cfV<]H#b���!�s�O5����'N�4w"�H���MSb��ժHp ��h�3� �R�j�[�4��ɓd���S F��|��4o@�H����jU]9�\�"��yU��,\{U�w|�rGz��X�._%Ry@[$�~�����l=��١ֵ�׊e�%������:]�2k�Y�lpBe�� ��:����go^��i�bd���a�Q�)���ǉimM9+x����k�z�{���
FU:GůGK�z&Ŏ��
�M%����Vܾ�JLj�k-�Ux��5���	��t#�70u�t,��b\{��Rڷw?���Fbd\�����'p�p�q�Џ�I���0�RsgM�7��5|l�b<��c�?p��[�k5ŭs�\7��l2Y��GV��d��6%��9���R6�G�4M&��r.2�L��ٳg�䓎�g�.�C���_{o��򹢼?�������� �bq�SH�Yxʩ�x"x���x\�XK+2���/ѐ�����L���+��C�bϞ>�L\�p�2�r�����$�xt�_\�k<ê��t��KPLO�m(�Erlx��|jr�k��U��``xhɱ�|~��T����I4EG[�P#y~3��4�c�è�I><����@*�5��Ba ��x#�d���Qz.U/��@q�Ma7��|�]��l
/��{�E�I�H�&�O�A[fSèXz�"���	p�Q���#��d�ު�x���S�2z��0sJ>y�Rܺ�"��«o��"S���HZd�]���(Վ� ��07<�(#�@�U1���p~Zg��;�_�?\vEO�\�˾���<��`���^����|��t�/�1��v+�8~.6m܄��ߢxg�s>�,Y����C,�_���C})���<�Գ���-���#�y�5X8w:�霔��V	^��>/����<�v!�1�7��LJ��!)Mze���`ΜɈ7��ylڲ#E,\x�l\�0��xXp���Bd���E�pѥ�	X(��G}زl��ln�67N4�����Z�c��n��-��p�P�-_ï��IGI��#����/��*&�QH����T��L˹�����,�H���
t�5	�yˠ>��(t��Ȧ$:�9D_e!=F�
R�#�� ��>T�Cҋ�` � �g�P�2d�Q�����/ p�T������s�"�u�E˲)6!�i��ȟE�C2�U��2��"��(�q�bzg&w4!B�B&-MI����!�A��U���p��_2��`�Q|Gr5�q��ԼH���
O<�8W����^�p�l�۫6?>_���ҙ�
0���Z#�K��)���K�K���R0�&VJ�y��Jp�JJ6�D$L��rK���R�`7��
��� ��J�is��Rf֜Ҩ%@���Ѻ�gX���4iG�Q-��q�98㤅�����B���̙�:؇M��Io���'V�fR-μP�t������:��gHu��ϩ]�>;�BT��>�9&r�	��"�;f�����˫,(ב
j-��h�3���-�xMǐ�p��Z��j VA��YT��R�:.S�G5�k�Ή�H�`#�9�T������5E0��M�); Pn2��]g��it��gd�s�0sJ;:�Z��ڄ�x��?&P�KB�=f\1`�@�,}��J�ť�#[(H�� L�6��Ύ6�����0)��@"�C"�C�H��$9
Eu?T�s�̸�HfϚ�yӧ ̽�,J?�({P<.$	�"�Z���+���{M�3���2d�
�� �,-�
ع�z���_+.i@�糞����>W5�G�/=�������#I�����E2G�>o#jc�D	�qׯ]0����h�E�`�dj&^y�Ily�=ᤇ�*;.���g.V�B4J0ƾ�\	��(�A�Tn��*�����g՚u�l�u@=�;'�y�p�g��)���Q �upP�ٯ�}HX�e�-�&�BZ������>�%�_��_<� z����^~n:���D��&�䇵�V(]��9V.	L��D"�L��S��7�GKKN=�DLg�&5!҆���#g�І|�6DV@�I�XX��fϞ��'�i�f�opO>�^|�UdrExA9S�VB>7>��[����+F��蓯�?��{��L�9�����*')�~Ҫه���@�f�y�g0�SC��Yp�yĹ+��:ø�]��>�c\�t1��>�������<�~���f����>�LS %��x��@4~SU�� �q6�N�N�3E�Je&�h��q�^#J�g���A[g���o��k����K/����_���,rE�_V%6s�L�� ����k/ǯ~�O��0��?��E�H�����Wb�� ��a��N�w筸��O=��<�

� 2e��D*"��֫Sh�NwU�L�I�e�Z١�ܔ��3�a���M����羸n����nw���ܵ�&�w�|lٴ���o�ko���g�y&�:�t?.��x���lH�
X�n#V�]���a�O���ŋ1w���
�����;dfn�n�xz�N��5g|*
�`$����Y����{C��
�{�4L�9#�$�n�B2YƩ��%�.��H#��@P酊܈�0��%�T����j�%}QaRV�~���C�&0Ţ����"k�[~�"y���S��Y?�Tr�� �<�Z˶����C�
7n�tƭ�J�f�Hg�0���j��Dx�S���Q,����]��~	�8�I��%�Z!���%��,K����h��z�@�6~UM)�HO��*k*���i@@!-��oE�ڳB@���B�"w���b�93�w�^��/<=��1�J���>(�lf6�7)EJ�&��˼U�6����ތ�������������d���b4�s6n ��ll*��R�,N�:�ESf�3�C�t���d9��Ё�q�~�1<�u����=c�a�u{<+;Z&}ǥL)�3P5U�@��J
�Ae!��,'ηP0����������}н�ZA6�G�d`,���h�DE��9�r�E���X���FD� �|��9T�)�]8n�4\xƉh	{ġ��w�-�#9��b��J o:�B�I�ZK[���u�u�!��ah�%�������M�} h�9�k* ��;lj���<]ACϚ�E���
�l��� ˣ��[ �`p��@�|\E�Q�/@��D-_L�@��(K㹮赠�G��h� 
R����YU�T*5*�j ���?�	|�
Dk�̯2��w�����Pɉ��i'�Ǽ���' b�/q���x�^/{~�B��� O���bQ-�Of\I�b�2+�����i)<TK��{�74��D�-�=�C2�.��q�8v�T����������)��I�r{ѵ��mގ��$�� <~�q�-����Q�C*P�+�i�X�ש��������O%y'����v@,�DK�@?F?G*Τ�J gɂZ�|�ƽV�9��j��$F*I��Ô��5�x�׭b�A�<�(��'�� �]�>������گ"    IDAT�G{K���2,[v%ZZ"���Z�v~����}�}������M�&Q�����T*�l�flH%2˪"G�䟣Vƥ��SO9	���êU+�u�r�$b`J�)gK����A�n���NU�cr��M.�}}����
�Զ�dM7_���H�J24�֩7��RFkk+�3���Ǵ3��q����ؾm�$���&�'+� �}w�����1<��
<��gp�w\xd�p(��9�JpddhH*�D������&̙5>�;�m�>/�E�`��P�N&�X1)[�&e|���G�1�L����E��RI<�^Rn��F8H��Z�L��	7��@.�D*���1��D�&���؅ޑ�&`P.����j�J��zǤ���#72�i�:�o|K��T���g��#O<�#}8ܤ��~��\�$n�a	����"_H�o�n���S �#����g�����{�3gM��?q��}�e���_�o��r� LwH�A�]�G�LV� ��4�)t@�F0S1���Mo�p۵��S���{Z��s�c�������xG,�;n��>[�t�x �wlCk�$��̚�������1ӧ�=�b�������9ԍ#���6�'OE����.T�q���J �Å���k��a� j�N�kn$Kx~DB!il�E�R������ǡ#�ضu7����@&3';UDڊ4�i%Eቒ��I6��`6$�-{=��g��Z��)j.6�����br;�Ò�'݈Y�!"F}�'�oa���1k��K����tbf�T�&��WndS����8MV.
RN��fP���:�J#4%�Z�j`tԀ&Ϗ�#u��b����2F�/{��l�.אG���H����àS1ui& �Vv��]��T�� ��Y4]! ���7]��?G{�B�����t	�+x��#@�'��PE$p��9�)�[����(����>�	t���t"�fi9�����2�adՀo	2�xhaZR)��(���,w(WP��<9�yr0���EM�A�
,=s�`Hh:�����5��5��\��eeKIߊPI��p���c!D54�C�%{P�eC��ՉD����dF3E���x�x��d�T���[9.�VG��8j�$�O��E矁���E���d��P�y~����Z}�Y�f08���T|O+*MX}���u]�
t5MHg��R�{A�l���r,J]4uE@�*0�@�G;)?��ld�2�:��*�4�IӨv�m���w�A� �j:���ܱ٘Mw|S�)]�ݠ����/Ҡ��|��̼W��+Ry�YM�"�jֳ�eU���$#Q^b�@jc7���0�s���لsN9���DɃ���ZIhM�B�*��"���(���
Z�Έ!���z��J�{2�L��|�Hq{�'е�G�FD�}�L�ufϘ��N���-��悋"g%��Q9�UY~>u��!7X���k6as�A$�8�Q�%����z�N��8�J����A�� �>5�Kg������h�״ =��\��!z��1�b��GQ:�uso�&i|.e����ă�ۥ�C!���U1�UMl\�>���"����D�ң�z���֖	���?2ЇΎ8��f�r��hmJe�������O~���!D�;
F�3�(���˜3|Mm�D�nV��p��=REktj.�X*�����5�d���_�ʒ.q.
����Ī/Ar&��,��=�t�� �.+��Y%3��aYdk���ğ�y�|�wM��!/$8�1�]��jFL�x��"_��402�m�wa�.����r.�b���޻o�W�Sz������X.������s	H���,�7ED��`�>���s/{�����,U9�U]����n�o	-��a�����Ѝ�����+�3f̔
_� ����	%���2�F>��x�N|�S�JZ-���ρa
�Vڝ^��ֱg�_����r-RF�@�����/s�eYy��>'�X9vW�[MNJX�B���Ì5c�,-{<W�������m��e � %�D4Bdh:wWN�N����<���%���K�?Tk�j��:g���������i4��i���:ʮɛ⏾�{��C���<���y���p��p�}Bg��U�!Ы������b�N��B���-�2�S����w��{x�����$>x�T|Ƿ����ͻ�k�5!h�<R0��'�yX2Ă��!^��k��k^��'����/�ÿ���~y8�=xr�o���?;:��D"9�p�G~W^�o��?����_BrdD!�Hid��q��x��12�~��X̬!�/!�7�h �N���P"_M�sk�Ï2��(*=7����*m����U�$��	�M>~+�iFї�? �!o2<t��"�ѐ4�Irb��/�^ (l*�۔�j��"I�{=��J�,6��/Gv-�S'�#��B.�VW��#n"���ك��A]o(�P$�T��@��E�Næ*ȖZ�$�;�4gBl�D$^;O�<u��u���tx�l�X�/䰃�Ӕ�� MK��=t���*���@a~hV�d�D=��ڐ��ҟ���l����9����@�]D'Fq���ù��j�
�;�o��ӡCw@z=42�	<زi�c�
,� n�d%�`�@O%�vׁl����euR�H����g���r�����P�ǌ�z
b~�1\b'S�gK��p�ף�c�m:���Zz9v/�-v��Pz�4��ՉV"K���JZ�0.ȼVI�����up���$�S��]����&Ć�bQP�R�|_Pf)�����h;|���̌����$?s�rsv��p��p��طm�^y�����-�Ud2�㎪�iP�B��]��S�ȕ�px86�C��σ�8S��y�,�&dژ{[��$�fraag�3�3�����=x�|�	[��3\��B(i]N��t{�>Ν�-��i״���.x-̛ރ�OA6�Jd���-r���*��!���[_O�y ���		?�}����[�G�c&6G�N�I�9�;�ض�� ��<Lg��\]�]==l��E瞅��0�lp�Ȭ��c�������溒b�H�g&26���H������>�GD�%-=A)�5��e+x��i��^����|�LN��9�v���&1u"t��¤]�D�K�^�ˤ����
y��^z�V�d�F���S��Aȟ�0�
ef��3��ƀ-�>�ٲ�}��0g��.7� ��?�$����~~���9��A�~�/�ؙ���A1
=s�K�G���HO�Y�^1v������T���a�	:?��%�>�d�Z�bq����^]��P�}�#��ǯ��H��U�<������L�,��e�٧�=�${��M#H��8AF/Hb�}�+�߃J��	�G�RB��F��|&i��2g3�V�.�Nce��s�Y���J�9���N�n�h���8%��X�~������<{�Ss�_������%j�� �ϛ	���zU�ձ��"����ib�܁�KU�>s�-����� C\�K�i|��G��;Bz��{�؈ 4�\��ଳv`n�4y.���	��E��Ԛ�,p��kbA�u�i)�\�z6֔4�NEx�{���^�{J셢�4s#W�4�v��XZ�G:��_�'\|���x���*p�1�ς<+w��l_����ڷ��Z�|�*M���T�ԁg�K�C�V1���O�����M�H�C?|�>�C,, wP�[��u:U��5|�#����Hg��������~c�q�����`?�3e|�oᙗ�C0���?�!|�}�"������ _���kN��<O��cJ�B��ĉ�'�'V�J��ժ�U�����߿�����_}��� x��顿��]��C�?���L�����} �]�Ǐ/�|�+x��P��x4�ljY��{�l�G�~?���r�DCN���BjE�{��p����h�����pa)ς��~�z�!����k�k�����p�� V�y,.���\�!0pR��~v6��#iT�*^8%ɉ� hkT���$٘M���ϡ]�� �P���B%�A����U�bi~�l^H��ba��m*p��A�`Ӗ����1��Q��E����**��z-;�#̅��Ö������Bj,��뫃e8"�::"fRzKp7/c��z���ώe�!S�x ���7�Day�ZI�v����2��k�Iov��vVG]�-����Uq���
�"e�Z��#� ��8�+qޕ�"[) [�[�W^��g�pڵj]�^��	l��pB�H��ˉd<��H��n?2�=��t�PX��u��Iu�Y 8tp��&o8�h��0����kD�4	O�YS�Оp�Ç	���������#$I*4gbgX�.[��(��@�
��3�Tʘ��C|c�@�Ϊ�N��J���2�� �brj�$q��)���d�U,7���b~��;��L���3S���̉5%������ٵ��>���0|h��h�����"�R���	V��]��j+�
��Z�֤3&'`=��y׍�4��L˔hX�LM)�d�LL��݆Y��	�*Hmؖd-��-I�v�%�UBH�d���mqL�ɭd��da��y<�h1Av�8���m̵��F´�SVW��S�KSr�"��x+q��ۿ�b��ې�����$^pҏ,�����X�����j�eMAl��o6ǈ�Nh���D��D��ÎM8��pK:�#2%DJ����3!���*%�J�~��!����,�DRe�҃L�(����p�I��_�S3�8rds+�Z�J�����8g� F�{D���Nq�@ilWa�o�^d���o�᥷�c��A���h�D�
$��p�z�p�Kj
�R���e\-?	��,ޏ�зwj��{�������01����6�݂}Nk�����]$0��{I9ɜU�Zwxa�t�o����c���x�����sϡV,��gM>� i�S2u�]NĢ%Ҕ����>��?y�JHY�'�|����
o�}J�P�zoP�B^7��_�abc���j�<�4�����Z9�v%�6	�jN8�����L
\0�X��<p��)F��:��gC�8�c�Гi��-8�5���`O���%l�gby�Q���gǜ�$�/đ[f��En nO���@4�X�� C�y�-����W,m�YX]��<����8�h���n~�gϣ�[����`~nO?�GgR�cA`�m?:⹆BgxF,^x�RA9�4)���yR�4�~�i��=1�;v��p2�fM�X�.��B��zC{��vbuy	�\��u'�굢��ս��@(�;��L_���y�C�[Ρ������l9_�QU,%���Y��� ��}7|����� �Ɲ�aa)�?*~����.R������ߺ����K�#O�P&u��W]s.��2�0�?�{�?VV��n�MW\�Ë�~�$����x��i�D��ϒ{��"z�t\^�u���('��n�b�21z�k/���}��<��_8=�߾s�_�yb�W{.Ox(���I\|�.���a|��;0���p�O�"2�(�h�0����ql��瞍�.9M'%��Z˨x�&/�t�/�<�����౧V���_EÝ@d`M��e��&����|h�+R�`'��W�<�L��f�j�Lg&��s^Ȥ�>�P��*e�t�j��*V�x��@�C&A��
fO���l�xx]/�A�p'Ǝ�`تc�x�K�!�7C�o�#شe�d�.��At�n�,汔ZC�
� �#Z�����Tpb�m@J��Qv>�H�	��7���Ǯ
9�Y�=����6������h��ͪ��88�h[����0N�2XxX�R5I��Y�7:N��LA�
�u�b�a��"8>�׾��})��,�4���	&���0.�$V�%+	�ߛ苅ߢ�*���a �l�4�ɕ�(D�%@{n�F݆$ȸHgʺ���l����7.���V0hm L���d�g�l\k�w�s`�Z��;|6L4����gI#;u���&;�:m8����k��;�F�x�ֵ�y�f�B%ݨ�Nx��ؐ84�t;�Ƒ��B���r:�t��t��1�"�u,�q��i��i�Ь��f��َ����~�=�0)lIC�X(H��K�6V38:���l	�BM��&!>����䎞T�����P;�5S�3Z�Vyg���7�p0�v�08v�ׂ�P�|�Z��r�+k&x��ҟ��yLWP*e���0�]��	1d�/���fvA �}��F����?c��F�R	�E8�{n����mw����8Xo�7.�y�R��u����<˚��i�2��Wm��k�q��ٻ&���-��o�	 #�` Q�PZ�햁wt��~��J�:���e>3�Z���o:�'OM	8=At]n�/q��N��G�TU�Iu������;5���}/�!��ŧ�<5��Y�K�C�u�7�.�_?��
Z4���k�Ju��99�#d�Rb6ɫ��%|s��?��LA`?�w�gְI�b�^��>�����ޯvqH�q�l�#�1�qR!
Z���޲бU��: �ĉ�ߋm��@��g���"�xnZ��d�<7��'�[��ݠ�L���[���?��n|/"a�|��ƳϾ�����ĉ�rq�:�q�a�[{}�Iҥ_)�9��(�Ѧ���X��f��H�Ϡ�&��>U](�'_��pN����&>)�5YD.D�W?�5E��2c9��4�,U�yk�l�A�ꬓ��=͸OYp��*l,�A�CDe�<!M��yv�M���H*n�X�iB��߾���?�����S�����?��9{�ܛ5`�����S�%��
��0/��$�ڮ��_������к( ���Q!�^�:ŧ#���_���"FFF044b�7>�r�%��ʆc��Ć$c_f-���n����o�&&&FP�t<#�U*Մ�hv8x�8�y�x�Q�/��.�ڒ�!�<s�\$�g��4:�/���q�u�A���܏;�u/�VJG��Dj�"r��
z�on�4��������O?�?�f�Sߌ[n�$�;�k��x�Q,,������]���㟽�{Ͻr�Z�P���1�/�|�)(t`x�r�(�ΗvL�?��.�q�M�v\�E��S��CC_���<���8\�`��ƍ�]��/� G�Ʒ����ȈL���$Kk�hS~�O�'v�ރ��?O��R!���l���ق�g:�r[��w{���x��+x�g�Qw&�@&H~C�dG ����l!�7� �hL��T#��

��xR��xr:3�q\X�T	�Df	�;hԊH��P/籶��J1�f�"+i�g����O���`����U�-��)-_3�m[Zӄ�h�́'�G}Ɩ���"C����ض�l�oى\���4f�WP%��f&r���w)�H�Ŀ��A�/u���a��MW�0��+�=nL4K�@�����N:�Vf	�S����*�d`F��c�9�&*a%`|~�9�}�Q��E酼H�b�%41��{�
�T>�T����g���>l���c�F���!�eV�З�iĤ��
�rzfG���H.10(��O�Y�䪺��Oԁ�r)�!�F� ��K5�[&�-�P�@/�F]�������;�C��*��@0h��� �������M7���D�Ru0�=�E#z�B����%�d���F+���HHd�Xȇ-婒�r!�/`�P9���j�H�Uu,��钿�,��Ψ��]Ă^�߽��َ���r�6�)�>7����x(��tczq��W��v�����.�Pm����5�%A!l쵓�d�ڴ��vw�.�dx#��H;Q�����Y��Q���m�s6�Cr�L��-M�䙰ҵ��n\w����^k���I��!���<�τ�k�����"y!��n���H]~~u�:̙��\���;�����B���p
,���򕁨(�� q)qbRƉ���U�̾�    IDAT����..9w��=���)���	~@�)�
*g��ȱ�Ν q^�}�2>�y�)�\vى7ŵ=�3���.��y0��cf>������BJ�?B"��[�ؿ{�}aM��$[�o��X�	&T�"������Lϼ�6ϤQ���J�*���-ʞ�zq���G C�ؾ�v#�N�m�����i������Wٯ�� ���b�1Ʋ�KC���"��ÔjmY~��Uw��m�G
NZ��6��6< ��:�6�vb�`?���}�Q�8tA�W]]q<��,���E7�.��V��l�>���w��믻� l#�;sz�<�J��j��r�n�?���=gM�%���y�1��F> %3%� &@ٿ�yEU�����j�
傰�:5�M1H/�F�#��B�((�'��������2/G�z�;u5�(�۪��RLn�4�����7�qϕ��h1��^��Orp/�H�Ӵ��`C�����4��ND��6�O�3�~
���C"���^ZƗ�~z�	�.���D�mx����`�WV�q��!���l�:�H�`�k�]@"G02�^��8�eH�l��l� �.�?�������'t�C\��!>c)5$���ra~V<������>��<�˭!�+"����GÝ�y'�����Po3V�D�Eu?����E$X�Z���@��Ͽ��o���<�G�{������p{�t�P̢V�` ������/܊R��ǟy?y����q��=|���-��QD#N�}+3J�a���]A<�ӟᡟ<��`1W�+< o *R8��fA�f�A^M��:t��\�����6z�'n��?}�#����� ��o|�^;>�����P"���m[��^��x ���P �y���@"�g�zG�~��QRJ<2`�c�G#��uW㼳v�C3'���Zp<:n/�nB�z���gq�xm� *]rt��008��4�"J�JV��pD���d++)Ʉ�{!���x�>-T��� GK�r�j�Z��%T�)8:e8�uuz=N���p�X-���hx�!���8���F>��ԤȒ1��a	�ȍ
���Ф-YrL��~��0�}7������=H�"],ci-�B��eYizeA��d��(�,!4�pJ�P�	�C��Ȑ�H�ɗ8���ZH8��Z�sKX]N��M�]͡�_3��m�auԕ K�rN�"vJ��8s:�:;2d���Mc8z�s�����	A���R�_NX4���F�ZU�||x ��`,�쵔�0�g�a�լ;����������>����h��ĵCD��{�="��I�L�y�� aN-\�-C�d�^$�Rr�ZRҾm��_S+�
~vg�A�����R�$)�´\'[2�T?)"��ČIy �pHE߇� ����V$�� ��@c�Z���љ������h Na��èXk!W�`.��4(] }~��:�譗e@6`��6�`�P?F#�Q+�R���g��S����/�e�-TIʖ�8:����"��¨T�14I;���evW�N������.6< ��X�^�M���0%� 0	H[WB�$)��aA���Y^!Llm��P�:Mn(ԤraI0*��ޱ��l!&�Xk)�j�r�d'{v�hC��@5���*�,z��-2�]iT�N�����ɀ]d�Z���}���Aŵ���p6q�{q��qD���e �u�ϥ�bȳ<��[s2��h&��L=�CC���X�Vh�%�E�������Xmcy5�7���󨷺���Lؽm �vm���8�m}���K��P)FM)�>l��fO�^<x��=��l=��PDv�	RAE����ݬ=Q���`v����(y�`c�����bcA Ȋ5��߆�B�t�ӭ��5��qz,6K��([X��k)lY�ʢ�G�Q�2A�Z���¦�$�����8}�-��4�s��Z]y�� ���Ʃ*�e��9l�:��}�pݵ�"f���B�56���x#*D	�Y�WX�T.��'�]���,��P'*�4�5�I�ku�,�
"��,�TȻ�x��W�G�P%��9�⟌/�m�<~B6i:M\y�����kd
Y�f�p�8�:����."~���Xa�Gg�����$2���H�Ơ�g>ak���Z�O�Ƈ����.�yg� �sL��Rk����-<������3�r��:q�?>1��<��,���g��U@��i4�u):�y�d����A\���h��5M$�A@Wi��ɱq�B�Ԏ�ŵz��CȤ��j��_�"���#��Q��Xt0^C1	�|���Y����P,���{�i���=G[���E�W�%����a9��w��{�G(ל(V�*FixجW�&n|��?�/��o �m���œ/��#3�(V����c�����閐YY���Ŗ�	��=<��Oq�#?ơS�H�:h:�p���Fc�-A���q�0İ�gAPM-���2z�-7_�?�����`��ǿ؄�����O���?{�O�ON�c��(���=���y�x��!lپ]t	.������o�W":8�@8�\��b.��x瞵�r��p�]R%�X]gG�p8Ps9��{�����h{��`yv��|Oj�8�B�Ie ����� ��e���X�C���vb�o�n̜�`n�8V�Qέ��*��VA/'F�ֹ���3��[�J�_�_X�t�Z����"k�����8TOq�`Cl\ ՠ�.�M���	��®��Ǿ�.���$�?�sE,����
�Ocl&)|O[q��L�չ$Q�ݸ|A� �7C���G常���7^;��Z��:�E��Цe.�<���N��=/�u�7m�!h����lɊyt ��r���ͪL�$�ʎ���tȗh712Џ��6���Y-"H�;���O�B���R*� �͗��O���E,3<���-��]�Mbl�YbG��+zC 6Deʭ2p���QTL��t���U�M����T(b =z�N��\(�Y� ̳��*
dCI��dX"Y�"Ѱ������`�.''A*��ٵ���:�I�\�k�JC>�?�����B��L̺Xʗ1���J��J���:�*�嬦E;��p遽�<<��x� ����Xw���u�N��x	�p:Eচ���Z��cs�8|r�J�Gp&|v���Vo��������V�ygQ�	��l*)�8J���6	���a�����.)~�;��.޷�#a_U�좀���~��[-#*��Eh��t�x�Ů�QAJ����~r�_ϗ	N�2!��s��_z-r^,9��QB���p+�܁�4�`��}B��:<�6�v�˄�N"ɻ"���^�G��};7���0���U)� �"z-6h��Y���N�rE�=�<�nD,J턗�ȏ��4%l �+>G�_<�Q?|9]�[Ǧ���iT]��QP���i��=[p`�6$��:��l�)8�߽�ї��� r5���*���M/j����"��N�o2[�eZ-�܍S۾�����=��Ov矟�N��Z6�;�������}��a���t��R��zd�KSkZH8�&�l�����Ss���E2���n�_��̓}�V�x���q��C�<*ȯ �F��L���H����2v�،������ ɘ_g���m�L�8���x����T�6� M�&�O�_�ki�S��.��Nr����s�D�Yv�x�7p���O=+�;_ ��'yks���B��ɪ-�~�-���Ʀ�a�Ir�CاဘB�R����4���?���4u�8U�����l��H�fU�=M09���1�L"��������W�����1JE>Ө�s!A��8<<�͛&P���0��������t �"�XS����|�<˸֦��0>>�I4�G�>ƿӧO#�Ja��͘��4��l�p��ƫ�-�R���P,�qť�`j�b��
N��uB�&d�|��q�7��J�$�E��B�NQ6�<�$��=ૅ6��K��p�u�A����|_�z��UN��x���iD��뿊���Z��{�C����1���J��l�� ��󿉑h��*��=��Z:����'�փ�G��F���j���ۇ` j�UPf�������g�;�li�d�ݷ~����߳����/V<��|��q��p�����xb�?��;��+.��� ����/��R��1I�4��{��?B��$���mINE���g��MW]�}۷	�I�Q�1��`Pq Mg/�����?�R;O�u����x�Q/��l"v��0�v\dnb���s�/�D2C��Z�x� �KY�8���N�i�RSh���:����_F��yM�X�QU��R��chu\� � %b˝�Z���m�p�8�da�'�XꆒQ��[�Ax�Il޾{Ͽ�ѭ��d+-d�U���c;!��9�f���lN�<ة�؍�M�+u�}�j����"� �cm5��_|E�d���`��wk�H�]0�4_f��Ȳ �����}� ���ykB�s�������2�}��(7*(7j*ԡiw�&o�x|�016��Sqժ!@�!�򳅔��/�`v~E8�>�PXxv<BA/��1)L��T��āh4.}z&[<@	=��	sL����W���5G�L�F�����$���}&�$�^���K�d��/R�h)�Ù'\+����4�2�r2�X�9S�C�/����&D�ZC�PB6W��jF�5	j��Ӕ/�sc���H�}�{D���Z3+,�_���B�YG�����.:{.=��?�>����C�F4z*W��4��;�^&n4�|�lI��KY>5��\�	�4�1�̊:�͚��x;�ߘ�ڂ�v�n��	�~�Zv�,l��ڶ<�=	�b�:y�V~��6t6쉀:���[r��&���^�K%t�daG�I�=��Bv�8��y�(X�G�!;��eK5�h����,F��$x&1�t_����e%Gv������!�򺙘�[Cx^��G����p��;6�&\ݦn96s�f96K-��c���4;L@{��K�`��F|!�Ԓ�@JB�Dne��B��M�a��$Ws5��[��sH+��'a�J9���7��K.��PϜ��]��K*ȑ��)+�� �`9��s����çe�F5��Ã��A	�� �^��ɒеȕ�ɯ�$���~h;Y��V�iI��	>�/6d���^���.�8D��>�߆o�
6����F��2�EzB:M1`��Q�!Qb���KDQY[ų���ǎ"�P�ʪ�	l�e�˟R�:ȦB����v�݆/|����k��/&�nrY(.B��&
nN;������D�@��>�a�N B��O	c����p��	W1vBF
Y�@$N��#�.�{����;��������.�E]K	ʚ2RƲ�k��h���]���O`d�DW�Eio�<.!��0��$������E���#J�q5���'m�&�)�y���+V>/�v��S����}=*'z��,2*�1oI$�06>�\��Ϩ�wt[h6*��Ţ�Kϗ�V+F��
���
�s��c�A�����̌�G7mڄ�۷[�3��ţ����QA�{ahpP1/�͊��N� �a���*h��&���	A�y�I<�G%���Q�u�l"�}f&f�c,��%�R��=��_�#��}�"�K���>�;�q��.ܾ�ԉؐk5���GB��-�_���#�o�;�<��_|�up#��������oo�{/؃�׉&���T����퇾gdŶGfVQo��'�׺T�#���G�pHk�0v� �U�m�}w�r�_��߿���~���+�z;��C���?��p�?�srvo�u���GP"NDB
����	|�;╓+��IHO�!�/W���Ӊ���ƫ���Јa[3������s:m4�)�F��i<��)�U�pc���pQ��x�-�sH������c0��@�8�A�&��k�V�rN��x�簶� 8D�A]gKw_̋ZfK�'Q\Y~�h�R.y���f����C�6����JΙҼ���$L �׭�q�JB�ny%C�;p�ڼ����۲K���J�fӘ���V��t?Y��c\��3�{r��^���$o��XZX��'P��st�Z�G�������I�� j�V�f�ϟ�P��c8:'7Ȏ�B��zl�$��q�5�ƻ.��R�@�x-�V��v�&'é�aL�Hn��4�5���9N��[���
��>���Q7r�~���	�$	2Y�^���	ǌ�!���5�ă�C)�,,.c���N[��M��زy�T��)��!Y�$�T=`�Rl28;@�`�Akj5�T:�r�&a����aL�� �:��H^���e'�����A8[b�i|���\��T&�͏�'N�¢���*UM����6#��DGdf��R��i�^\U��%���V�������dOa�� b~���R[Q'�J	]��s����ۥ���,����V׉\���tY�Ǆ.[�[��.C �,�������̬Cg,����K��V�hC8d�g%r\��S�z7�"!���1Q�ђ~t9�p�{���V2\�.S�>���2�ki�([+�Ɇ��J�-)[�GΨ1�\��B������wE	��`"���i��2dlө6ɨe<�5)��mQ� �q46��V1&�^��y$��#g����@{��a�Y����ER=U�����S5�t��d	y7�����r�:f��d�-�Xׁd�}	$�~��E	y�m��K��|Nĳ�j���)<>����*��$��+�#`A05֧��G�I��Є�G1�2�U�+=<��WWQM�2y��ĵ^d���nْf!�� �z� �ɾ�^�g����!��	���ɑb�b��^������x8L�YXҘ��j]ym�z��QK�Hs�Рr��t��"A�3kx�'?���|*EP&����_��̧"[�q�����O7��^D࣬ ��e�Ra�F	��l�0[�!䇞9��`&��flI�z��8�!ω��0�&�T��}OV�J��r������/�/��-��5��T�Qj�$\Wl5����������P\���o4���ę������P�e��S���Ԥ�"/s�1G�)�Mq&$f�1p,5 �$ľK�9����pziw��}�y��H�e��yo
F­�R��K�P��Tp���'e�rAf���I�[u!��UB|H 6S6�Q�����#��kl����YN��F�a�DaieU1���[N���L����)�<u\ӌ��1�#K����8:>�`$���XYˢPi�����p��-�~��nL|�!�=��/ܿ���_v �v���x���cf.�B���I�(W2��������o����u����������r�!��� ;7\��~�ո�}��^�������~�����n�Z��׏�"_j �������`*RɲQLwO}��^��T����]?���{��O���tջq����6:ddń0�M��7��_��}�t�#pGcp�����w�1�a��8���.�ܼ]��¢�F�G�=���n�����'�;����� 1r2d�_����V0>֏=gM!A-t�� �&yTJ�zp��	,LϚ]�������DP9#� �ת�S/bm�8��54����U��!U�TB�x�($.V=d�9`'�r_��5
f'�����\n�p��Í�b�O!���|�&�6n4��[w��w_���Jm O�F�!�>%�L	8�cd���m%~@i��8t'���`&aT�;r�tNZ�RBm��!�@wR����c���0��ˆ	�!?+eGd�(�(�[7��T���o��E�g_z!��)��פ=-R%�9�61�L`����c���c��`#ф8#o>�16�B���:���GG��irL�b�)���4���W�A
L���g�|�KKH�
r�dL��XT�"!8��y]�&��Hp��I����`�b�}���[X���'%e:9�	S�&ї��p�$~Fve簖��    IDATN�ް��nM��+˩X�4JV���'N
�ȃ����տ���C,2]m��\8������I9èy:�	pٹga�н�t��à�TW�z���ujϭ�V{�+f,��P�
1�i0�r8QhtdV6��aa%�b�aГ2��!Ɓ����"%^
�����n�U��� 8�x�硱��$UNd����mR3sg��_l��q���:P+R��"�[G����֖TP�4�� �% :SZŃ����T'��?$�?^wWe���3W��:��<$H�0��a��D���:�5�P'�·[\��\{�ᤫ�D�A�����^�P��lՐ�15ڇ�ݍ�c�����$a׍?J��"L�h�������������YzRT4��U)��E"�TA�}�(6Oc�?J�\8:�D���)ȇ�B��A��������C&_�\4��#}1\y�~��mɦ��MaF1N=�99=��χr��L��S�%�|�(N���A�Ѱ�,��$��Lf����n[�'�3*Y�����҄�eȾ�3^vqa�+a|uk�d�3S�s3��޵aEvajs(騉c���)kY~5���0M9�~�HI�F�f��\�
^~�i�>x�n[>�;�5���Mڷ�L�wu�m���o�l�u�\������Z�&,9;��;6Z��<q�L�L�C�5�N����C�H�g��s��H���Hؤ�V#�1جw���M���c�q�������Ln_N�W>@�����X@6�ZV���7	2491�zW���D�%�/�y�˰�n��H��b�qL���	�Y)����R���+��� ���{�h�,g
����qǝ�bzvE(	[�����-yѐ�luv�{-q�&ƇQ';������`2o��L��sB��~�TY�Ĳ��ӧgԼbG��!+�]��H������U����W^yy}�&���V�T1#O �!��ˏ����L�2'܋9��\Z-L�����p��{p٥099�`Љ�t/��&^|�~��A,.��X��6�%8�e|��_�_��籜i��'��#/qBЃX��:VgN P���\�����8o�4�@6���ދ�|�[��r���Gg�&�rDrj]���T�3�VuHƹ�Y-��:��_�������4���_lB�L�������|�>��_v�>��� ���=��)��?|/��&���yѮ�Ь�0����_�����"�'|��N.�������4��ޣgA�YÓ/�ZэH��Tb�6ҹ��y��$!���+�aח�YbT�}�ſ�ӗ1?=O��dЯ侜YA���`2����ԅ�O��I�Yʓy���m�C��׋-[�h"@M��`2�]� R��-�T"�!�\��IXl�e6e��M d��BȪ�hE	ǆF��[0�u&��w,��BQ�L �<���C�b+�5�R8��@� QrO�IV�ȡc�k�x#��(-�D��L��a.Vv����V�eT,25�"U�����r��d����X�;�J��o�.��l��.����y��{���j�U�`jr��٩�4�j�]0��Ǐ�B�م��Sp�{��FU���Q,��c�!!دB�Tj��#1��i'M�� g�wi�477���j��rrdE��PJ�+�.�+h2���r��U௔� ��Ѝ��E�r����!L�����֌y4v�]X��Ҋ����pTk�I�@��"%�J�2V��p��G�z���`C#I��T�6=�DU��^�St�[E��A���E���������A������L5:dwGD>vlVBv�F��q��]Ҁ�&���i9,���8$y��SR�i�XL�U��E�v�u�[��3��R��zւ�
U78�z������#l�1�z�N��Q�&��yx��>Ƅ�P�B�(O	��[/O�����fv�+USk� �0ԁȢ��"V�2�i$�BW]�7�0	��j(�}� ���!��c��c{�F%��[?�a��@,�m�a�&��M����n�bQ��VA"Bdf6���5���<�4ڏ-�Cr-�!�g"Ԃ�����vWI�׸\%�(���xGO���4]�ˈD�	�Ѭ5$�@���[6	81����U9���I(%�]���XhJ0=�مU�,�B>�n��vMat8�(9L�(�H�{��"øD�P�6Pn'�s8��šC'�Q��� �_q^�/!����NXR&6� wҮT�ΞxY��S/GWE�q:>�b�n��;�51�gT�X4
��uH�Q��J2M���ф��)[V�� �PY�.��O]ɱ[&|ƣ��lN6�ig�ˉP�ɜ��O?��o��^��F�Q$�۪Sp@u�9�04��b���}|�un$�)�p�X���0vi�����9���%e)�pX�"����.�,OM�|4�
c|xHg+aH�v.S��	_G����b'O����
�
�tz���E�L��f#�͙6�.Ɵar�(�}�e��s�&	7��$4��dV��i�̵L�)7\/N�wZýJ[8�1��?2~F<��;$��aH/�GI/�h\~�hp9p��|�λ��%j�x�p3VX���3'��*��H���c2�� �K#���^��I��8�|}�3�+P*Y�$[+d(�R9dÌ��?�gP3Sw�c>g���pD���"��ge2�'�T;M�q�d�*b56�V،u ��JX�L�6�yghrid��څ�������aDj(���{����w,��P�wQ�2U~g7�W���y���}O>��^{'�id��\^tȟ[]�z����>v�� �Nd�{��R:x������J�FK��=N�|~x}!�!�k�wM�;T3K�s����}ꆿ���H�������o��/:�O���&v��H�����Rx���ջ��g_~=o������p5�v���ބ��=���_N���(c�}9^o����q �p���^z{�J�"��ڬ�֪��k��� cx$��d�	.��%�"���2����'�x괔�:�,�H9e(������N�:��Z
n�kF��z��I�R�:Kč��t4��*T����ꓚ�z�׼.:ҩ�V�ݪ(����\�ǰv�γ4&i7{�V�����o��QL�}�cSh�|"i�[�!þ֖̪�rґ��-3�w�[���7�M��t��:6�J���ë� 7{�|�Lhr@_�2j� S�`��1�m���L�k0�H���8�a����п}3��е�z�^���pX���f:��Y[�ԡ�~r_�Қ�����3;��F¡Qr�m�l� ���~���h�@�C!].k�Lc�"�A8�� �j���N��j �Z�u<_k��ID�w��y5	��J/���ԍx(1���$�y1�i�H�@��v�mp��Z.�X�x�A~Ƕ�j�sH�s�f�p��ך8
L��x�E��\W� B������B���a�Ƥ�Āۤf�/���<fWH�Π�ȣ�_�x?�s����V���Sc��$D,�8P麂He*x��I�8���l��8p��ضiD�0&����^�VSң��q��<r9�.ٸw�F��`�i����Q�zgA`:���>5���-2�!c�DɆ�,�*	�<��A/7d#WHI;xz]Bk5�\����0�i@��]���\���gL��1C8U�$��4��xKՊ���<+S��Ũ�{���y}9�#Q��(���PT�Hb�0�69x�m�!�=��ZJM*�7p�c�"C��j7���;X���h
��+��x�:=��������\>�^ZƉ�e�Y��J^�@\1�\vc��崽ur�� ��)�S������*c-�1���ť4*5I`����sv�=[�~�l^�:��,�Y'�sR��n�NŦo�Ǔϼ���B�axLb���B�K�'��2�({�<��O���!�����DɾR��Z�lb�u��!�T�� �"	�R@��Ʒ�6֡���Ǳ
�@.�@�&�>�	�^NBioEWtv��J�8!h7JH�<�Є韟����|V ڄ�PA�r�T�!_�q�"�iٖ�P��&Z��<�������$�%����Ntju� �5�-�F�һ�̿�b\�CA��5���J��k��<ë�|��#�i�C����Q�	J S�lP��(���_O�G�S�Uh�����D.�yD(*8��K����|��{����d�d\�]{Z�#6\�z���|LuyV8��Y��g�Uʈ�?|�0N�,"F���j�h�"�ÿ�6%P���pt��\�|�w�`מ\�7�/���4�YE'�,�lNxx�

6u�ߚgmO���@_��)�mPy�t�/�H,�uO�(��4+�E�g����������h˫��f�BQƢ�� >x�5��Gn��][��p{<��!����+(V��7q��C[6��7܈^Џ�U�ʤ����Ϯ>�K�;�Rgm݌�}�j\�k/N�:����<�9pz��khtz�R�>��E��]�d�b���-�P8{��?����������/MA�������������n�W��������G��˯�C�=��<���$���-/��CH�:�59�߻�V����XY&63,<58g�R���A��E�L�Zxk:���*ܡ�T h@VmT�����8�H`|b��R���.��?��'�dfmq����o�IY'�C�#p�,�8w44)�XɐcI�$����I��L�HX���^7;��b)�h8~ukY�͎%-mp��VS�h��cϘ<��׭�����&���'�r�Z�M8���/�Y�_�Zϧ�n�C,85�=�r�2��خ���h�����t_ؽ���pa��<
�<����(/�@��6ŀ�����Ј�$cg&g
#�0j�[���]����l��4�{|�L�٩���j"�HhĘM��7�`bx�F�=��%�J��r�D�
f�5�&��]ܠј�qDc!��9�g�Ǣ�^oK�he9����7v_�NEGN)���j����o���P�'ל��ouսx���h��b� $��atxcc#�Y#mv\�0�!q��YKM(1�)K3�Ti`zf�LQ�>A�=N�LA`�x��Q�����A�W0)�K�İk�݆�=\�,�aa����j�4B^��,\�/&�C@��%���O��f�P'O���^�r��l���ؽe
��wF��.������r��8���8rt�3�|t\n�E���{��di���b=ѷ�+��A���3X;��cc�y9M,�>8	��B�����k3��VJȮ�Q��Q.�(�.��*�RR�A��B�� ��C�ZG6���Ґ��2�ǎa.W��gA�1 ��>\�0|����(��	��h����u\5_�ŨMb�I�6�JŎ�d�sf����̖��'/AMv�Y�6j(���훰oפ
��g�&(��KU"k*�����l��(��XX+���"N�,˃��R	�׆�K��h��6�ɑ>��m��qjK�|���.3Ki�
M�d���O!�/!"$����={���+�G�׆��iu��-�'��׭���6�D�Bx��i<���XZ-"ѷ	�@��1v�t���h�E�Dx�(�*e�(�Qc�/Y�X�"��4'�$^�C��b�!���۱ԙ�l�W2֞0Dz�����Қ�D�]��'�<$��}�iZ�8��N���p G�?�N��:����
^G�P��U0�l1N������������5�?\n5H3)�Y��d�m�Yn!*t9�ܨ���F�G��m��~�S�X�~f"�6	�\�[RDb�E$!�)6M�����l��E�YM�`�c�bm�&�v�v�����0Me<#�)��lT�e	R�S~aA��Ӯ��W3 #��n�.�u�$::t^(�y���4��
��4�:$��q�ё��56�b�0\>69��O�|9�I����Ԭ&���S��5i��W3S��iҙi%L�9a7^|��'\8�agf!���x���@����9!qE��R��8��d�'�)�j%L��⒋`��ޅ��>��_'O��G�?��՜x�$-�Li�j��H4��@?\�It"!)�l˷�SF
)��4
9����;%�==?g��.7��
�
�2k�+/�ӿ;�:�H��^�D���jf!ζѯ�����_����Ǟ�����Ϳ�;�W_v�徫�{%�nǫ/��~�
^x�f�3�b&����8��W_��wmC���+�}�(��66o�"3&��2��ܖ��r��bׇTՋC'���U�PΓ��b9���*)nD�b�C�������wF�CO �Z�F�T
���2���{����6h�2(�R(�����N��t�h_X�p�Lz��Z�j�x^�/��Y$ͱ~Ќ���k)�r!��H�)�yq3���kb�S�-�	_*��G�\�I� ��v`�������\�5v�}�_�����j�4�����8j/��AX��+Ȯf��Z��<EB�(��r�%�[CD�@���,�)n�L��?7!�
/;i�&�<���]�n�$�,�9!�Y	ݤ�68���@	v1(�֪�UA�=,�d�x�a'�HĂ��!"�$:<:]��e��%��lA�";f��:\���ԫe�4	�bj�8�<����X��g���0��f>�2��4t���>�k�#4J<$�0�m-s���{Ȯ;�|	��(W
�.�'��	#�i�ۂ�3�3X|����v411�ĶM��y����jˉ��˘]Jcyu�V{wnŕ��-cIx�jW�#'�K#nJW���B8t�4�� J�ʀM7�Zu�&���}rL{��&���W�K*���t�|��#H�*pQ���n�!ȓ(�1q:#�h�Nl��ܚ��Rܱd?�} ���v6�{�"0�L�,�0X�`�&��"2˫H--�Ʊ�mt%D��6�y}��'F�'^��T�i�K� �R��Z'��k&�*��7"���Abx�xL�a,�@83dw�n�\!�R����Wb~&���g�l�Iv����'��,�	�T�j�QΧ��l���{�aj,7����Q��nBi�E�K��Pd�����E>v
K�Yt�4SJm�	�Xp��:���>Mp��
���	�<�˂�Eh��F�XÉ�,.�
B�W.�1<ŵW]&ߌa��|l��!7�C��6���͞GO.�g_�j��x�$-�t��脝o���M�XU�G�3��MI� kơؘ�� ���5�Ƃ�E}�>!�bP�M��F0B0#)Y���M5�#��m���c��[L���p�p�:��zx�D
Ut�g]�k�H2�P����~3�D�\Q�(���2��zfB`e�s[��ru��U&��
M����7n��C��H0��QecM�4���4)ƅB����w&�$��9���xI�\�g�&72S3��	��$N4Fq! �<���s�󔿊ϧ�.��œ=�/�F�o�i'���r��4΢[��-���T���6�=G:����9ْbԵ�}��̻<.xk�D^�i-@S@^�8{����}��BQ6Ձ���^�s���Y�^_ιs���%�$$H2�L*��s�����Vmm��Z�\��1�	#�H"�(����FI�C�t�_9ǭ�z�wf|��?�*��L���y�羯�
U�*ZkTAb��4L��k ��꺷&SdM�X[[�ԑ�ݤ�͋h]^�>�믿�R���c�qEg�P����oWt�V]�_lڸ{U+NW��[4�V��?��]ݸ[z.N�i���^F��9L�oqy�jU2e�	g�ZMt$���"<<�2)��~��#��)X����&�����=���b�TjuTic&��O@�>��P�����'�j�:u�2K�}SC}�����~�(C�������/_Ng�w:t �D�{����x
5�p���͠Y��S�P"��o�����"E��j��t��t#C�8������>�    IDAT����]<�����^lT�ߝ�ᵳ�h:�Fc�W��oJ��#K8y=Z�~�;б��1�]����zn��4�;w��E8�e�rk���Ѩl�^�K�ʃ����lv�SP�U��b�X��9�y�R�1�����l��i��Η�Xp^�pďd"��(&��~�;�M�կ��?��ǸtnF�`�MD�r�����Y��+܃���p���@09�����hs|�����M�%^n�1�����ʗW��tc-���]i�Ө��9/�IZ�Y�7D���KCS0���� 3�	۔!�ؔ!~�o;�7~�^�G�����a=5G��Jtujjؘ�%����
.�.!���Gd��wW��=� $@ۿ(z������g��U@ԽRmaiuS>��Ey9ei	�b�j�L�E<B*��0�M��L�Pgspya��G�l7��Q ���'��}�.(Њ�w:vԉ�x%ТO�ym~U����Ng�j;��0�AE�5 �Tt �~���*�H���R$�]� �q�M������VWcS6Dk� n<���N�'L�W�f��m�AuQx#q�gN��A�Յ?A�� �bA?�ڎ��>�3��H}���*�jM'~���pn�kt��8����+{C(�Ud�6�#��C�ᙃ�jCp���>��^�.^GN��!lm�Dg����u[aq3�Z��F��R.�J��=�3�A��}�᥆���;��u��h�K�%�d�&xݸ�(8�B>�E��ޯaп2=�r��xɁ>5,���;���U|*�Xz�ȩ��j�M�����+����S��e�j9����i�d=;:ǡ=۰k�a?�jV�%�Kt�4�e�H���MN�����u����YB�z��П�u(�}+���_ "'�\����Bg/��r� 
�����b�����cj}� ��6�L|f#���$�I�h�L]�7�ұSXZe RJ@��*�,:S���'�UJ�����j�:R`�����֘����Ÿ�v��.�nil�6�=���@��t��]mTXs��cY#[{�fO��0:eQȅ���M
�\\��B�8Q*P*��su0ڗ��QǱ���ʹ��Q{e�Bl�Rd�ز৻���,Xy�-Tj�H�a��}�M��wtQ��s���>�;�׶��}H�_k���dcP�z��Ϣ����<Õ��!�K�_O*�5�t
�9ɣ��5��p�V�$Æ��3�㤛�5r�Rq٢H�b������f�|���"[�!k�a�gM�]�^���Hi��~Z3�.�E��;�?Y�iF��E$	�o1��L*,p*�	T���*�.�8�ڳk'R=	�8�&2�M+;���Ȅg�9��e4���[��rEZ ���צaW̱�a����ѣ8z�z�^xAzi�D34�:
~1���X�ҝ(%a.�{B��W[{�hVdܑ�E��m�N�D5�R�H�K�q����Ґ��n@�"A�?�TBÃ��Ƚ�f��*��i8^Ts�(.���0�;���z�4,�(0̜��ܥ��Ia��s��QC����75���?��߯�����0�_���W�,o�I� �J!_�I�é[8�'�R���q�iIX/�!������߉�}a,/����<�S��ƽ��G�\we���P(V�!��:��=.\^~{bW����$�ڸ:�B�5��kr���[H$��S@F�z6���"6�f�]^��]C�ZP3Pή�QɢU͛�1�N�cn\n4�3�>L)�P�J�;�.РC���Ƀ�� iBSSS��������/�V-�С}�G.��fzG���C���,..ṧ��3O?�'ϠP�H�9?������&��1�>|�ߌR݅�l	]
�N�%��!�)*o��(4�NW��:Dr;�e�H��Q͗��a�[A���� �#z��7W���7����lVr�Prn�S�GW�����~?���tyV�.�&z��U��ѡt�Et9��F�I Xq��63e��Efؘ�X^��"j`;�
�Q�{������D��RNo.E�D��d�fMv�"G��@o����)�4�@�99�ha-�G����5~�mZP����+�Elȹv��!��ȾV��nDJ��q�f�*��(�=�����U�e�Ce��lF�-�ɥ�7D<�4�6�J����u�q�
Ͻ;�px�L�� ���(t}Jĩ���.r�Ƭ��9�I2#�އ���qL�bd��	�ܘ����/#�;����8{aǏ��Z��\�8����1A[�.���e�fTg���u%�kü�	�*Ux�Y�领vš �
��Nt�R�aaf����U�E4+����v2���Q���A���O-���٧ج�U��@�0�Fԝv�>�D��O�S�6�̃3��"[��q(8��:����#��n�ݠ��!��Z���j�X[���������T�EKaC���8�`���l��W!W~W^r�8�>�j^�sǩ	P�̮lH��)�銍�]`�ȡ 5����q<4i񵊬���]J��5�źl�)P�T��)#�[EOO7�x {wmE��D��@��}����%a�֤�_��mV3%�8y��Q��	�����yV�&��J��I�'���\�`7!�xXz+̬Z��C��x���8�b�g;m�g-��@C����`�����;ż�k�Y6f*��³	`6���,��i���ZF������P*�N!�W�y
���<^�j5�����q-��$8��Qa�@p�*S
C��ǣ��R�
xS¶��f����	���bE�/ݟ-s/K��#��K�G�"R�9! ~#�o�iB�:�"��nD�,�Z��:��@��Ԩj���Z�_g�ҍ	k4��3�m�a�`�4�E� �R��&h��t[��������v��k������kh�v3@�� ��i|�|<5V,�%8�|��m��vuj�M���NA/��.���A�>�m�&q��	\�|����μIƓz�l
�6ۺ�y�רյg����v�v"ƿ#����Oׁ>���א�~�\Ƥq�LR���4Dv�18�E�@&_�C�m���|�c�G����d"�:m1�\s�֕M<S_��AFϕz��@?�##p�"����t�IʲO�ג���QC#�C�XhAJ����N� >��.��g�3�E)ߤV�%���?=��O����������/�����.�o��/��%�zŹ�w���rЖψ���"z�^Loŭ������9|�_Av#��~�<��l�Ws?0h3ܪ.֫m�rz��Y@�F05 8$n|M�|F�U��;6򭅶���PM��ӈ8����S'�p�Z��!��Q�o�VJ+���,�>�����-�21���6�*�Խ׵����P�,��A5���H�l`����am�.������s��?E>����_'����	�Umc��"����'���o��d��oL��/�4<�Y]G�e����{=6�U��w���I�eC�'�D��V.c��0A1_���6�@�wq����A�! ����9�M����8	���әD"l��`tvC@Q���n'&������a���ЊPms�*?l
�Iu�(/��\ʙQ���;�W_=#��X|@(+�uD�>�lڍ�>[:)�\����eC7htJ�	y`����%�����N�)Gν�$�R�krQ)f���ΐ&ڋ�AY�T$�嘵V+#�M�T������^9a�q���BX��IP����$���A����"r����?r���U85:�����,�I��VA�Ot�n����%F*B"��hE�\���e�y��F�7�߅��荻�B[�Ѣ����D�]�'Ϯ���0��A�EA&��{��̍�#�J1�n��m�.������CB����\�[B���Ój��\�,�b��}@�IsS	����BJm$�
s���]���v�%�6���Ni5�K3R����B.�x�6WV�~٪�6,=}���>�-�S��g3�RD�qC��f��¦	��2�BemZ�b=���4�<T5]�b����sB�\?z��k:$�I��kj��Ĥ�a����S+A�v��t@E&-��� ��kD����t���r�ڳ}�����ߢ���4�]�?�7dф�>�BE���P��ߥ�b���mB�B~�l��8���c��0M�b�r������,�\E��k�&����M7�C��E��@�`�ǱD�b�H`(Wץ)u���KK8{q�kET[N9���DMe�Ll~���D�8�
K=��M	�%����uަ1���7D٬/�V�17V�! [xC+7�׸�slD屨:L���M��<L3��U��df�h)���4�c,v��{P�X��g�Am}1�_A�\��f���� -��@Bb+<��N��"�7���vC���ǩ�����+-�.r�	���ִ�ʴb�ĽOV������UI�q3A���U����{�Ӵ��O%E�U*9��8���Z�� �� \�y�����Qj�E��笽Hoa�P#��Zt�i�!���f�
/tW��f�d>'M���
��c��1�����0��Ts��~�P��j���B�D�Z��e�ģ�퍊�Ө�D��f����vE����.xf�2ן� �1��`)���P����#���@�
�S�h`fjFǾ�����¼��I�N��F�HCC[�-VQ(���4T�{����YS'f���n��[�A����>�}�4�&x�k՗J!::�V�TV:M�5! H���Y]:PU+�M ̄�6P,�~�@@S���}�p{ec����I�n��[��1�?���?���vg�l
��?��,9�E��zv�_}���]X+�#�;l<��� 6�=��%`:;�1(�eCbڤǉ��w����'�ۿS���>�}�����)�5-vk\M�F���@�z�4^���p�©!r�My󹹹�f�R�/���,70�׃j.�מ{
3'� �E$H�Y]@�\@���L|�Jd�q�zq�-o�G��6�߼�N�8��"�D��=�����-�܂�{�kDix���	�<��ڒJQ�l�7��J9�����?$י���=�wv��`{v��Ėm��x��q|�[��w��O@ǋdr ng͎]g�B��	���w#��ٹe��Ia�+	Q�0�7���A��Z��8�r���kX_�@n5g�d��,PT�qd��e����!�e�)�ݲU���!`iǆ�7c�G�����0�&�0���b�*�6d6n�*z"A�F��0�+e�����d}{�Č<����.��Rq:F�0ЗB������dJ���*
Ŋ���,+Y&�k�Ǣ
t3aHSQ��6��X4��T�X}=18X�UK�0��{�
Z�,�5������6Q
����"a+t���C���z��Q�Ě�Xo��c3���Z�F�T��^��zUkqaK��6�LzS�ni���=;�0:�+�7G&0�g2������e9tvn�`*�¯Uˣ^������>ml/�����o�-�d[�t�F��-�!ҵ�t	ý1���[�/�t����Zi������bu#��t�fqiam�v&�qB1�!��n��Z��Km�
��?��dA���TtV!�f��Q�Z���s2 ��h��:B<�s9��ϡ����hd�lߵ�8��F�J "[, W�&��av�
�T�ψ��D�
Qb�.-���y���u�����-//ayn�h��!	ȩ%�IA�$��6��~�Oi��s�T����K �����\��(R�?��VJ� U�j�}1�?�]��q|R/"@2b�,�~��'��iG�D�dY�p��� _�)Ř�:��F�,/v��!XD���l��5$3��`��X�PQa��pҴ�^B�XE�Q�����@�{��O��8c��m&'-:���)��
Q�403��S��q~n���p���uU�Fp���돨���
��P|N�,�H��
]יG�h���ۥ�iN<׬u6��7�,a�VC����ոџ�%}�M#g�}�8��/Z��և5�j���	q�x�� ŏ�N��9���g�XO#D\�a
Z7S٣�vdp��i����cf�<{�v��Z;l��r�sO�>����S�Cֺ�F�ƞ2Jי���:��˽��=3��u%A�t~�ea��W�K��ψ��'ɞ>x!��Z�
m��c�xf��DA.�e}V�� �J&�s���55�HM�)��V�܋�1Eo��ub�}5�l����g�z�Y{?o�c�N��׎|y�{|}�t8�B��$��a����o�4�7�q��qM�wLOJ&�I���?#c�z�nY.�� P�DE)�s1�����ҙ��5@��iӖv��	h�f{�b5|����@�iP�� b��~~s3#m�����~���ȕj��r�6;:e�aٝ]��o��o��6�Qo�F�~��ؚ0�af�G7A�ق�f�^�>�H4��)�V*q�無�i�{�Q���Q���WE���'j�p�h�!8�{�o?�����nٗ����ҿYC���<?�_��Wg7�$�e�M���9��<�ޕ��@��>^�j�V,���0=���X[����;��c#��*���_V�7�HK����;7Wd_�H���nur�حʞ�+w/9�.���2�!/j�4N��6f/"�i��h"����ʂ
?(l�c.�J�زu����y��������`}3�W����`pp�M��G��F��.,b��� �Ã�MB5�ř�x��_�_�LBݽ�v�mo}��x:�K5�|1�ص['���Ep��,��7_�?<�u������!lsFp���1�� �%���0�3^Ӥ&���!���sM�#�U���p��������@�hS��xR��1�P�k����X]��n%G�߭�@�Y2�ĵmb`�6����`xzs��(��"���c��02k���&b@K�vۅՍ�&�f�^B0�F��!�(>��;ɛxyuU	��rM�4�J.z���Co�nC=Z��M�8�mq�����0Z��P(��:i�ϘNy⺮Ԫ*��YP�AR��A
	7W"�����ur�̃�p�$��T��R�S[B6�r#�������D�V�'O ��F4����3	a�����B�(n�0���gN#O���sl ��6Z5�n�
�İ��ca��_>��T;nxBa�*�;�v��b1Ԯ�Ь������c��-�5��m��2m3���fh�z~v��VQf���-j�,xixe�u
�.�7_��UHQ�%��Q{Re�ė&���Ht7��|D�q8t]s�^�*�*Q�Lce~^闉�al۹��Q�A��植��B[IS��5boŕ�$E��t�S�Yi'm"�U<h�����M�H\��&f3��l������G��m�B؇�A��<r$��f�,��TO�69��d�hc͘��C���k���q�Q5��}�0n8�G� K=�+p�j�+���n�(w�� ũ�edK��x���gS�Ϙ{h��G�T���Դ�v���J5���v�	�`e=�7N�`m�4�Vng^_7�x�I����)��g���}���[@�����5�~j��8}&̨ط���!�l7:J�DjG4�3��+o�F�9h��0�l�,Ꜩ-����u̐G>�lJ͔��i��c9qI�f5�f�ZX3Q�T�1x���x��O�٪ʚ���}c�_�*˫��15Dn�h�lp���v���FD�!��Ǝ�lo7�{wO��'�B�͔]Y�Z��Vn��᜛b�ȯ�~:0�5�s��T�gis����ip�7�Cم6���ܛg�p��E,��kB��x�6���E�-#j���&����&zRq��J�:2:�ϖf!n�[I����5,�����@{P66�^�`�%���^ �i����<`m���bE�
[S6K�p��p��S�y��{���=�܁������a��عc�&q��./.��s    IDAT*_)i������&��>�C�`t|܇lʐ��]3!�����B�eu�i�E���j�l+R��8��{���V�x�mL_�O������!P�~��pS�o&��KN`�,��V��5�f{�,�9�� N��a�Z	bp�a��˥�. 5'պ�Yj6����:���2)J�R2!��7��K��Ԕ0���F9��yp���~�����O<���i���^���׾�������q�ӛB�xS�M��{��`^�oUt�&ǔ�{��yq㾰���v�Mx��a�֭��R�N��[��!����;�҉E�>��P�4�^�TJ;@�8���S�p�T7��nM	ѝ]^����+��3��Kh��(�� �^E�l
�V�HWYB��{��]w݁����Tr����������LLLj�)�M  �3.h!�^��)v�V�@{�D���i|��c/J�C��[n�A��ܴHF����a���Xo�q_�[x�;?D��F49�HlՎ�����;�6n���C�'-��F�����Qt����F$��{��,\�E'����F��)tG�U��]��)�Z����y4)�kg��{��v�!����<J�n눂Æ���ɱ!Ye2,�bF�Q�<�kD\�B�%���M�x��QP�`o
I&n*q��l!+�[&����U��3�6�p'��BE�c���:�ZV�@�I�hժ*��m�5��
C6f�i��Dr�h��hamm�/����bێI��2��4<9.71��A�n��5��AJċ��@'f. W�	�VfC$���>�(ڪ��5��k]�\ǩ�g�}��}8z�D�Hۮ����@.,�w<XM����y�yv�R�`\���DM���LK;Y��K��3����w���i��>	���h#�/ W�b%]��f	���L��RG@Έ��v�JW �뫙��5�j{�7��H�M��_��W� &ǁ�fIt�-xju46��-,aci�f�&�섏:�`Rt
ч�S�0@�!kjF����p�%#$�x�^�^K��k��I�Ԥ<��z	esK�QD��ss�e�2�����|�
��5������Ƴ�5֪OacJa�N�j��3�bSXq"�'�%&�zj�vnCiY�!� 0?���ƶ�|&�4�_�Æ�VG�|���q�yJ[�v6BјV�)�U��:�w�No���\���V�NӞ��,�\ؿ��	�%�
;Em%�R�H�G�*��Z��F������x��e��f�w�%qa����p7��2	 �b���P�Q�If�H���~��p"���ڲ��Z�����,��1���7)0A�gZ�J�`>ZF�k�n�8[h�:ZKR���l&��Bg�[�i�uw�(�.��/���7�ݑ��%�N���� ��\��j[A�۷M����m�"�I�Άў�j��^-��}���h��aq�&����G��j���-��%w%���w=����~�}���܋/ɨ!OJ3�sT����k��W�D�!��3���a�i�9��f��2�Ӧ��qP�����yf�
C~<�R�3K"]��g�TT�Ub>�����I��Ҕ��NKK+8u�����p�i�Apå��S�#��G>���!����!��@*��� �(r�fff��e�<|/��)���>�Mg͉'U��K �E�����l*$W�?Z�R�`�r��х��4�S���	Q�����p�����v;^x�U|�?Ź�9t�L�%_�dvH�+����&
��A���n��&��V��R���q�q���F�6���k=%m��&�ȻR��%k@�oK`���ʪ2�t�Оפ}s�s_Pc��"�rys���~�����+��_=�Ķ/<���E���v��[\������*������	yä�4k5����[�
����ҥE�]>5#�	�t� �q�͘�܂Q|�tnn�u�kz���x����Ө��g+G���P,B�D(~�Iђ�	E���rǞ�g���T[z(�Wp��c�XY�&խ�vn�[�q�߃O}�c���� o��t9��Dbp	�X4���H����4<�)�Z\\�ɤ144��;�%X���}gϞ����=8r�\n�&�1l�gUhLLLa��n���ěg�<���<�:�:�V7+�Dzq�{>�m����F	�ٲ����,��5���aO≔�T.�>���%t��(�a�*C�,��6�Y�57Z^�!�i�p��\�jq�C@��E'�C#���?��lф�\��F���&kT06؋=�[%Xq&�n	� �~=���@�N�@s�������!�Mđ��_Z����e�y�
�-W�H��&g��
N	 v����dum�k�j����ăe��F�./�Yt�8�Ř�BX0RLZ
�b�3U�H�-4inqK�+HD��1�D2�һ�F��Qn�^&Rp��Q��HՕk�=�R��
��D�@�c�z=Ȧ7���,�RG����,��89��ޠ����^�}�Tj]\Z���i�)�?�8�D�s�W9�ff�n]Q���4{�ػ}��BO<,�D´b�Ց˗Plg��87�����C �1��wo�iEK!�lβ��AdL
$
����D��� ��!���ɩE�R�\��u��y��qD�/���!�e�NU��P�~'�N}F�~�4 �>Q��U��;���&�}ΙK��V�yO1�����xuXszIԱY�"�al��z��s�
e$�]�SL���0_�E���hL'����V׈�y����z�]%u�fr�i]ؗL��091
?�:�ذv5ᠠQE"�Q0|j��l7�i�"V`���J�p�v�р���S�Fڊ,<i��\kc#W��r�έcy%��n�K��&'�u4�m�H����	x �����#�Q.glj=^\\������jN&�ӊ�a��Ԙ�Db�I:u\�D�=�i�R-�3$ji�?�
�^����r�+U�Lс[�o>]SX*A�U�vڴ3�56�5�vT�˚Z��=!��d�)Qظ�:j�������7�nр��9���/�x��"u�!#Q�Ȑb1C�*��1��լi���[o�g>�1\d�\�:n^��x�rЙ�5�-$5(�)0���eѬ��**���۲E�"��{��WWã��$6��[`a�������wq��Y��a��������msj��9	fݧ?�q��waj[���%m�ױ�&����^��ѴFv��!���.�H69��=�)&�yZ`����f�Xǽ��CXYY�SO�
?���87��?��'��BF��7=�O~�\�a����ӿ���g����䍔���u�+:8���Ԁ���Ȩ��k��f�_�f�I�_�Sԛ�����럛�\�\i"h��a��m��;w�_����al�v��ǿ�7��]�8=���x�u�1nY�<1�B�<Bw�?k��ɱ�O��k��B�E�J8d5A�4���v�&��׎g?�èTѥ-��	r�$i6�ҟRW�=՘Y$U惡J3�s��6�޻m������|�37����!��?=�7_��&�y��>���Z?���̙3R�c	4:]	&4��0>>����h�z�1�9y�uu�ƃ8|p�~����Y���Rn'���|�"�z�4'������P��r�D|[�=���0h�\E�퇣V������&����PZ_����a��)�|N�v�@�'���t�����u;Jłľ�Xuh��\T)r	+�.���'���о������+#�B�����f��d��ʱ���^��؈��;�ՙ�#W<�c�
p��%,�n`xh���~����x����X\�`3߀˗�F����8t{��8�
U�J%�n�3G��m,��t�xc���6��r:�z&���"����\2Hj[Aj��S})�ǲi�p]�[?b��pV�`2��X��#A����O��k��F9��߃����2�Mnm������7�g�%�b����^Ƶ��H%��I�~��+G�&<��$��I�h������$��g	ʛM�o��g�E���1�
���J���Z��͸Y����fDhĞ֡V�����%5��q��|J�dc!����&s-�  �Uɝrn2����76����l��$jN��z{1<�/�5���U��ƌE�����.��ݎ��~����U�=�YW����'����*^;uAH~�w��d�,bR�8)`�%�r�Q�|nD��">$��łHF��E�ㆩ4�r-��gW��+o`v~�hbѤ	��d�4+L늓������(�7n���9(`4S���>�q�wk�M3Y�����js���D�^E�VF� i�N�a����=�9��O���x��8��#��鹵^H��ƁM���	x��Ѵ�:�E���)�犈����ST+�ʠ�f]v�L�`qށ��O6}�xq
U��ӂ�O��O�a��nK댯��C.��ɟ;|� vl��h��Td�ָf8�,�dY邋���L�)[RWD1d����C� Î�eQM �gf�`�}&-����ׄ��aK+y,/�0���isk8La|4�];Fџp#�n�k3����G���S\��a9]���q��2*-'�
��o���V,?w
�IC�$�'��\.-�8�,�y?T�u4��Ɩ��;g8}}=��������a�{����-PG��W��u��X���g�gR�Lcl7��L�ŏ��Y�["O6�j8]��2ԇ��<~���7x6^�RN���i��,ǵvCNc�r��_ӁO}�#�O��J�!,Y<���I���Q@�y�6?�v^34R���@T7c�ˉݨ����CQ]���]�Xɔ��E���O>���m���px��F8�w�0D)�z5�T��Z5�ٟ}���'0<���6ܤ���TrD��T���hjI������h��W�f5�W��)�7�>��18�Q�Xp���4�x���Շ���^<(�ƹѨ"_؄��҄����(����P����Ə~����+Zσ���I��+6�g(.fC�ό�'O�縦m�֝eMl�O����u�t�c�5���!H&E����O�Ї�����?�(N�����2!�Z�k�ə�S�purl�>$��F�^u�\&>5�8�Cj���0g�j/�.���1��c�t���T��`l����H[�=Lj2� '����;���O>v��&_���ۿ��oyh����g�p����Gy+k�${����������u�͢�|�����3sJ�3A������s�{b(fr:��Q5����	��p�翹�_��M�mك@j@´]oܠ9��[�����<�0�)S�����y��D0rc��i,]8����X]���#�д���wݎ?��}�E�Y��	��0���:�x�˝���+���/|�o���g�	�yX�g���|�@��C��ff]��SS��>=�(o�V4�&U�Q�%[33����Ho�q�[n�mo'��<��o��kobu�����CxZ�'��}�Q��V�:��3dB,=��:`!-m"_�T��V��V����,*�3@5+$�A>��$z�n�ܚm�
=���l��1�5>dC d��P�������0�c��+��
&ɏ��nj�<��"�Ƒ�;�*��ː�^<��,.�c3W���>��'zRI��+I�
S���\�$��	�q�ˆ��UO@�r:��z:����4p���1���yV��5�'�>Ģ��5���^����~RFܘ�<�K�.k���9 �����1>ù�/�7�|DN�6�Y���2^��b�nSEe��ǖ�Q��/p"7�.r�99`��.+cx8�Z�QԘ���
��+	7��&�7������s˘�[B������{%���#��pz�px���T.#	ax�WB�N������>��J����~��1�:sQ_0����u�L5�'���썝h�ȓ�SWh���l�\:���7�k\�հ��@�"��4s%�Mس7�t�.`��C�!�<�y��!W����]
g�.���hW��uoX։:ܩy�M���`ь:&)�_<5ffWo��9!���\��D^�pQ I���xT�A�VʩtJ�4E�lG[,���s�Po[�c+�!l��>C�I57.iVҙ,VWױ��"�����n��@Q��ӌ��ȭ��J!�f���/� �-�l
���)��>R8Nd�֎�����X���3;�%r,�����F�C;�6��XZ,ay%��L+�u]�d*���8��a�xJS� ���.4��>#\�	n��Tj`n5�3������E�X̦�֜�*��N$��̨V�(������	m%x�����eM�9]$�-�V �����#~��'q��,B�B�Q��<Y�G��,
�튣"�Z�vC`'�H�
/5D�M#&��B9Y4�rl�wNmAms?��c�.���}�Vw���ӓ9�#EU�c^	q��:r�5�����?� �{�(��������aSGʅ�K8�Ϲ�َ4j��M�3J��P���}5�-��sM��D5��Ťpx�TikF��U#��c?��}�|ESy�?$!3^
�	�l�/�\,��m���ޅ�>p��F8DK���i��\�;M��U� }.V�ߗ����3N=�Z=�ߍ���e�x�wR��@;݆��ϯ���/����<���sp]������}����S��[E^]^���S<��w$ 6�X Cãz�ex������^���ӧO������\4[��1�#)Df�q�>d7:Ϯ�����8�J%�[�y8<2����߰��a5�<�#��7��7G�M���BGG*�,i�v������|]�\��W&�&�����K�/��8;�2��r�ʖ�R��JU.C���j}�ω�!�$�q���irIH��Ԋ������V.�������{��ɷ�i����۾��w������������;��PƗ��E�򩧕�5��;t�ؽ{
��6�~������u�Q�%S��w������AO�\U�assО�o0��ۋ|ˇ���=~��ić���D
��h���Q'T��.D8R\+(�������(m��+�a��I2����${�����ě޵{&���}" ��R5>��ݡ���(�,$/]��������zFH+Ӂy���
�����'�\�gЮc~�D'��q���	���7j-,�/aeq�3󘻼�#Gn�;�y�F�?�y{�2��h�
7>�� F�����w��V�BQ�:6��9���i�S*�Q��ht��ב�����y���!6��S�i& �xYH&т�͞��}��aű˹���A��pS��9�o'n���cd��W��_l���ҦޭV�(d0�e��|N�4VL��8z��wxQ(\W��/��iCn�
���߫086e� �<���B�:3%x�T��u��٘��������z�u�U�%9��G"�M��g�� O��p��Ff$lW��!&�	A�L�]O�4y{t�*KCȢe9����AT<HX��ц�5z�s�a�Ɛ�����NqzS��^�˃"�K�l�7�Mo`p0�����T�M~�~��-P�����{�/�"[,����E]�B�s��uHcAp�L�����I�����N���BC��5��PؚˋLۉ���������iX@��+�%�/��nt�[���6vp�w���`&"SVc�5ˍ��{Rq2�k(�3@��X0����;v�@��C����&D����֘~��T��Q�k�����j<�\gt�����-�[h��f�ڬG5˾�?O��E���".�=�b��f�z�p�4[���n]�P�X�ɭ��B�%t�����&�bl���t]�h����@�ƉT���L�5pmNnG*dޯ��h,�H؇r!�j���?�T8��\<s]&OFZ2�#�w���F��B��3N2�c��m�Cyz�S[Ӣ���`T���j�/g�d2e�ll��O���Ė�´*j    IDAT�CS�Y�VM�@��
ٰ�.�|V6�u�y�2��
ES�Ky�e����F�06:�h$ �h��<Ξ9'�����1>��
�l��x�hz����gj��v�";�;v
�?�4�e��/Ӵ�kV��v29�(������^�6G��mL�uOX�i��'�Z)(�rj|�r���g�!p�ڨ��Ɖ�M��DUm*��{���׉z%�����s>�G���>���3.�駞E�\7)�.f�0��%��lԩ�26��6z�dҸ������X|U*%Q_���4����T�#m��p�D�Z��\�o_~/�|'Ϟ���G<٣���V[�X7j��>�[�z��Lo�@�^���E4LS��NH�&�,����m�X 4@˿�nR�Ʒ44����7���[�2��h�36��)�ǡ��_�jU�'���c�͋'P.S�@J�5���ކ�����=��S4"���Ǐ����_|M
��a��m:o�_�y
�BS;@���/�ƌ���8�K�}FH߲,g:+cS��׶W�]����Gv8ġ���}���!���ׄ���e�}%Ӛ�ź��i�! ���\A�,ꐱA��ٲ�}ޛ�7]�ܩ:� ������Є�����k�d6uЪ�	�Me�+�qш�w����M�S�gW��zx��������~��`�����\���w1���~�Aw0r�7����;1<��˿{���#x����ˇ��x|A��[������@������%�����F��V|����`*�r�lP�C�(�i�Ɏ���b���<{��mG��6�,v�)�'O�Ⱥx��|n� ��)XL�yk3��_:���E�6� :א��mbh�(��ȇp�}���H�:�b>�qΣ���Y&}�i�Y�^���g���D<�j	�G����(G]!x-$��(��h%.lf�P(䥅�U��>��|��_^\�����W��,b��V|�bpx���w�������
�&J�6j%
���">���)8Ca�u�����V��?��=���\/VP�WP���e4�.�Æ�虜8�M�#����v@�E62�M!g�r11���!���t��S����C{q���E�Ը��|N�����FI�Sv^���uJ.mɑ��h?��D����Zg簑�=sP(�f��W���`ЇP�$r2ԅ7k8A(�����|1���F��9n�q�<l(����@�,y�}��޹�h�������)_�#_丙�1�Չ�� ��Y�u����6��� RL;�dqנ��*���0���ۀ�Z�o4��~�ʴ����fVt=���]�&0���f	�V~ҏ��6e��L���2~���`u3�p*��v��W>�qs�!�#���A8�П����L�bOκ��X<7��C�t7�����v�t��.�p��y�={	�2�7N�YD^3! }Ğ���kt,�ݚ��)S�`B\G<�E[_G~3� �F�����~�ޡ�ט�!;��R�(rl�LH�i�,J����Z>9������R6J��h:���lz-�x�uz|�}pO��I�G��/]B�I��0�&�"�H޲�5�󛇼��n:m��k�e�I-��@ۦ��pJD�\''
,�,��/��M\Y������F�$���hPS6�DX7)(C�p/j���2s|N��ˡ�BJG��E��A� 	A�o6�6�T⡫��-ݻ��8��書<���r�Ed
%�|'�c^���q`�{��j�Q��7�������tQk�Qi���)㵓piqNwP^��3���὘�:(n<��g�����3���?��^��t哟�gqi�2fg/�Y߳k���tO���q��@������8���5��B���׊�	LPO  �5����D�bu�1t}Y	�l�iM	J��ڏ��>SQ?:�,N��C"]��7M �n�ۦ�`�ǩ� "��Ѹ#r�޻o��>rF���>��&���s����/�x~�s>fėlT9b�CWCy�L��I)!�QӢh���U�A4^<{�,����ajj}��W&�L�޲e������B���x���;���h�b*4Z&00T3BMM�T���"���+F���`�GڅD$,
�Xvфö���i��~���+���g4S�I�Sށ��&0�ͤް�<��A�О���_~�a<��+�U;Ңx<N��WJ��2���?��w�P.uv�����W����Z,�����+e�K����5s�
���>����VG$�B�A{`7v�+��%��sp�-��ߧ�ZOOGo����g�e�ʵ&������3��p����%.�������mj�U��� �v0_\QWnY�k
�|�d޾$:�0�td�[E�V
�ǥ{7N�&k�Z5��Z��Z�e�9A����<��W:朤���
h�ӫo9<�~�����o�]�WuWb;�����/��W�<7NOo���p��7����co��?}?}�I4�.����?��n9��ῧ#N�p/J�'�w���m7a0G1�3?�V$)���Á�ۉ�+95K�.������[N���`�S����F���7B5��u̝~��_�UJ#φ�K;1��X�`��m�̧���~'≰B�<ݖ�N�&=��_L^$�j ^��+�Σ���`7m�8�Q'���G~g#@Ȃ߹X������ؓ�:��n�r�lk�k(fJ�Ɲw܍���aaq�~�wx��XI簞+�Tn�\$�����r��FvDbh-��yC�s��f������Ppoہ�F��KH_��6�rF��p��J4�E�Eϰ|�U���ӡB�@� �Z�b�i�1jB`	�<��.�ȳ���p��"9>�| ��ڐ���Dg^��2�؃�-J�&�M�k2�#�s�P�|_���W*�]�)�d�D�P�h�I�!�Rt3���JQ0�S����K�Ɖ-���BUN'D�kB�>>"��P硞���t)D��62��Y�����R.�����_�	���[Z�+\SK�"n���#J�J��47_6\S�[F�X��F/�VKt6�y��{رm� P/��*�C�V�HӁz�%���8��^|n�;w���#��LF�d"��.�Ue���j�;H�jiã=��<J%�<��)x&�J�3��a�ٔsp��<^~��lI���X�JZ��\_�gs�D��6ȿ����"������ΐӌ��U��1���F��سCCC(�Ş�x��rö)@�im�ψ�}ͦ
��6~D�E�*j�N�DꢬyMP��'Ytq��nh�bk#x+Ź����<���bx|�����Y6�M;Aנ�lޘ`N$�^+ �a׎ql���P~�~D>I˴�N�lҰ��q![�b��".��au-�k�i]ۺ�6���W�iU0x���'�a�����pRi�]�h�؆B/kҪ5Q�c��p!	I������π��K�̮aee�R�+���E"�'�g�IVvtʨWr�F�m3p��r�ZF�>� :��(C�N����e���䙳!l�06:(����,!�x���XZ^�p� <�x��Z@&[�������6�];�!c��[H&ӏ�.:��Q� 'N/��Nca9�;�h"%Q�ֲ�M0ދ\ZsnKx���ʂ�nC�����ٍN�kM�(�MN�C^x�uחp�cj8���� R�8�!����p5���ݬ�I���^������?��{�n�E{��c�?����N3ׅH$�R��b�����r:�]��j_Y�	�i��n��&$B"ޫƈ������#��w�n�|��֭��ڶc(����O~�=��\��y��=|����^��g�	�����v�܆��=�DBx���X�����3�BBʭ�$)A�A��I���Ɣ�]�P�pP�H"�&�i�nx}&�altw�~;�^D�G��	�!���SO�N�+���&���NMm����O��w�.G�b>��_�-z�!K(\A�����-���[u�WVW����N뺳��ԚS�f�	�=��ƍ�[�h 3�����GNh�b�%�y�8w84}  �YK��#��#�`��]����9xֲ|���Մ���:<���Ǵ�u{h����چ�j����x�ɳWu�Q�k�ѱ&�T��^ty���L�/�:!��>7��1��hh4�/䮸g�1�%64a�����j~����]Cuen������?x��rǑ�����7����>���_|����}���{��Q|�wcߎmp�O��?<�~����R�1�k'��N����%TJ]��FP����������;�%�앃����7Kx��2������J�I�	�ހ-84�*��s�M�Сgw:��f��E\~�V/#�:��U�7��ti ,�	D�M��=���}عm�v�|N<�H,����6�/�����XKo`׮]�6�]y���A�I8dUXd��4N��~�������4����PC��b����'уÇ�`���**.�.b����6D��0��յ<f���5l�pG���������-W�A�;0�٬Pk���Ku��������l��2��&3!�bT�-.'z	h��5T�*]�6�M��9)����4%N��mzW���<��=�Ć�1;�($�1Q&w�"1���-C����.T���W��b�4;�7��Q�ѥ�E��/�`7�z�h�wj�����I��z����/��j�ShM��Q�6:K� "�Dxɣ�m ���PX�]�4Ʒ�xwr]���L�̰/#�fKʏmG�Ɂ�\����!kH,����>C�D�h�ki����4����B!+��'�������7�(�b�n0�`�r�h0�����щ�����C�B�.�&D���r��uN�7Qz^;:��J��p:,���I�5�S]i����
�܈=~�{���+���_��J�^8�~tQR�09��t�����1��>���n�bn�������Bv3�	A>�����x�Ԕ
�^�\0u��Z����/�-�٢ؓ!E҈���,q!_�Xjj�I�J!��(��e�&���2�g���y�gϞF�RP�50����5q�b�B�]\䴒�Т+V�S����q"@>4Qb�vZ�6'4LE�a����{�(���L�99�:U�rΝsR�Z�-��,�adƀ=���3��26\�}=�Mh	� D�D0`�BK�j��9VWUW�u��Ͻ��������j�^�N��g��{�7<��D2��s��\A,Z�(��
�� ��d&�R9�ρ����c� Z�.X�E�(�)S#MɊ��j@�ZC�f@�\��R8�d:�׃��f��@_-
GF��$;�Bn�W��ci5���%���J�Z��e�u�a��]�A89i�&`�P��"�wrd��nv���j,�KcS�1��T�"���2���}�.�ڶn��ZI� �/����;��u�F4��ڊ������x�R�����^Q��t���TfgN<Mpz̘Y(�g/Ǎ�8=X�4B"�Y���US�I�ͦ5b��ȡ�����i&A�G�/s�G_U9�j&�Z��XF�ۊ|,���_CnuI����{�b��nSb�K\�5QX��x�46L��z�]x�����/�B���#S����O�6%Ґ�DF��%���/S�:�a�c̤K�˭�v�~�p6���~����ʪ�IBO8�^�G4m}N
�+D��R8��%����w�y�Le�]�.�Z�#�ohmE ��}���|��`��U���1LNL �H�5Ѹ�g�N�K���A��^��T�F�<ig�T���`�Y`gV�w��"e��ho	����'{���Vp��y|��?į���y�8���2�����������A�P9#��'��ѣ8{��.����$��bfn�PH����p��!x�~Q�!o�ω��aQ�}�?<�x��}l2�5<'�z�E���L�4���ꁄ�q�#���?��?c���X�$�����;��b	�]�DB�"FnQ�IAԌ��ٕ�k�۽>!P��@:�e�6X(|l���A�lF^��jBM����N���U3 ���P�x����M���d�	;$���&���r��J��жM��ч�|�O���!�o�~u�_��3U�eock���Ň����ك���N͸z�"~��_�ĩ��=ٱ{x���ꗿ�ɉX�sU1�yǑCؽc#���Ԟ��%|�zdy�y=XJ�q~$��7VQ�4��G&�C��.`!�>�͌��V4x�(�R"�R"���f.����%TSk(e��xPE�lV��T2h�@ؼm��O>��턭\���	P]Zi�D�q|��Poz{�d�`�<>>!�OKs+�u��g�ٔ�G���2�#�d�ɚ`��qD�1�#	I����㮻މ�@��r&��p}tB��%�f�pcrc�XY��8�J&?Z��c���p�7�d�!��KB�`Í(��X��`���B-[���I�^�Ģ0VӨ�b0�R0閚Sc42�pM�#��#�v�9����1�"w�\�`d�"];M5�ڊ;y?���R�A�ٛ$~r�iv�~?6��nC.IY�<Hk dD]x�~eVb�`)���4�<u�X,(\��s�G�$[�BD�����}�16q�UjJ����v�	���{�0R�U�@��,r:�p�<����Ȫ�+�4MyB�Z�a�o�s�4�p�*��Ƥ�'�J�Gb�9��3�����L(���
��Q�k,B��h"@�{�,�=����V2 ���ի��󶭛�y�:I�j��\�1�k�C�9�h�V�u�#0�~����w�	1qb@.vŽ��;;�V�Z�ɖ0>1�h<#/��&�#��(��ɎX]Qϝ||<�覭+Nkk��T/�,t®~@�$�T2!X�x4"ϟdY�b���M���Q�E����#G�|�|����t^K���wbu�*���B�M�\o!���q�kſAS��b�b���s9�</<���^q1���..�&�V���S��.ކ"�l�؃��&��Z�(��R	��&&&�����ٍu���W���d	�K�vu�}:v�s�$�"m(�`�^l��P��n�,fجYF&�F�jFd�U�k@�X��"I���nooC���x�6i�3���;��-���gs$�W2NxD�TZ���b��~��\c=B�7W�.�~۝>�54 ����[p�ڄ��c�Id>�®�p��n4���RHg�|}��>��� �ػC�m���_+c|f�G�I�u��]�oC)�AduED%��������q`v��c�����,`"\) �FLxU�B}�
���BA�$�&�%Wܒٛ1+26�jTTc�|LdT��Z�����M���W�Z���.�ղ8��)�͟�)$'V�q	/�RN�j.���߉G?��V�
1m�ri_��?���Q����T%豃^%6��f�d0���Q��v����g��"�sr1�5e����������$��&�+�T6N�z�!���q�����@SS�4Z8��¼XU�"���t�l^��{w˔��������_L���l�-.gxx����>}�s��/Hל�����BH�OOmQu5
<1_�I3������ȇ�k�X5"�,��ً���?�����G��)� (���߉���'�@�D7�*^y�e|��'1::*
�F�E��,hҩ��_��PX���E�H9mX�S�ދ�=4�D����d�aA�����M0���G)���9�^�ի��q��w�/��/008�\����~�x�X�dEL �ɔ��Z�c���HT���H;����)�{�g��ʹ��ȃ����r򍍀�+2�i�|UU%{���T�+�a/U��y�����M!�K����]��we�K�=�*��E�B;6v}���w� ������W�~�4�4��2b�p�ߏmף;`D�\�|ǎÅ6��އ��N�?7&瀚M�}��[ZZ�l����t�պ��Bt-Q�l��L
'�O`9Z�3����ˊ�����ϔ��n���U-�Z]Etqˣ�⌴    IDATW���th�\L�kL̄j4��u��L�ރ�>� ���{���$�i��+M=�D&�+׮�[�='�d�m��H>�NI�����=}�4"���:�-���G7C��%�V�R�D'�Ue�>��BXYɄ����Cp����.�(�u-Ǎ�)$�Y�L6��6:���U)��K��o��w�`� Q� S� ��
�Y�/Nv���m���!_��`nd�XV�`��Q��	��y)OgDv�X.�A��|��$9a4�nC(���U5��B�cqRU�G> o[#f�9!�� `BBK�RQ�:�,u6��Xj�8I4$��r��wd
���n���f���g�3���3���������D��v� @��^+���jMLFUa��@�N	!5�� 7o��l$!#��)m��jH:)VOY�K�B��_���=�
���������N.ﴸ"�`H����zq~F�7���p�L���7����!(t^�R[��ǋd��ɩE�$��Ĩo��=����Z�)�&­��Q�r�t?5����+�i��_e5e��MyP4�Y����$(3�n;�n�L��<
�Pŉ�M֬�PQ�Q�wV=5�RJX�K'��8j�_�w�CNG>/{���Ʉ ���chh���'D��r��S�Ј�Ⓨ��uID5�VI&ד�F��I�-J"\���B���s�H#��ߕ�Z����N�*���n��R�J�J��)�H�!�,Zy،e�t7HA���F���tZ��V191�kWG�ɕD1g`�]=Dp��`s3�8a��D�($p�@U1�;9���ٱ~��z��@	sn3���#Y�X1� �@�J�''q���ilܸ^��8����T
2���9ȖL���;�U>0kQ�7T�D�����ᒂ�X+�鰈0��;�V����Hf�S���XKea�:D]*^���^��]w����|*�l����'q��9t5p��;�n(�t�Y�`rn�^���}�0��C9���Y���`5��m�oCs[ 7�
x��U�N, �����(���"JB�dLyI���&�7j�vs��)��Ĩ֓A�^��v��rv+���rq�X$�x��_!9?���)����2�P(��>6*��S�È<�� >��`��A��,Μ������KW�e�0f1Y�椓됰9~�X�d��mҽ6�H2�)w,Acɼ"ܳ p����	>�7�8�s��I�^�jiD��W�D����N��%5��u`�!P���K�
i��yr
�
��p:��>���ؽ{�\��Ąp)2��?(Ϳ����+W���D$���(��ɳ]�+�9�K�+�����>���`�d@*S�o��w~�#��W�$�3���|�s)���O���x����PTR�/��|�K_�	p�\6��a���^��SA!Js��J<l�h�9��I�&����gB�cc����}�u+l��zA�{��0Ꮿ��Qd���������He�x�?y��դ4��U2	饱 v��A����ӏLN� �R��hD�X/�yC���]� gs3�~�ٚ�uQ�
�T���	79'��r�����g�K1KIx60(�B�'�{���k+;7�|�C���?�]R��s�X��_~�aW{o7`*��`]O��؂#{w �UNo�p��|[��o;�ͭ-B
���0l��-��]�PRf-�2SϘ�e&�*��Ud�L,��ʩ��D��5����z?jƒ@�,��K�w��d$���
⫋�O����Jr��yT�Q�~ld.�����pz���3Ё���8�k
�4�>�t]��B�+�Ï~�c��`۶m�Ŧ��;.p���q$�j\��Gss#��:0�nP�諡�B+R��ˢ�_�-.,`iq�h\
 v'��v;�l����x:�Y���E{{~)�s�KA0zc�T��Uk =�a��È��X�AU�Jg�ҭL���nĝ��6_�����Q^[�ݐ���D�F�C��B�����<��VA�;��4����%$?J���
;:N2�n��iLƅӳk�Ȏ�;�%�,7����''�*�[,h����As��Ax�UuM�E�Y��%*Qհ���̼���H���I��.�H�q�j��@R�XD%Z�i@~�t�D6�A9f
$��vv<	�bW_�
�K��?�κ�4"�t�dڢƋ��J�S����I%��ت("��$iF1*qtwt
ƛ�NvIJ��h��`�X.D��S�9�5}^<n�n����G��m�0��&�#���s`gkݺa�_�M� �8Q���L�x��ͤ>��J�?�� j�ӌ������_3_���Ѯ�&�2��YK�G���y�V����C���Vo������`�@(�����0�Z�a�F�\[T��^�8'�U"!�J�W/�Y(e�5�XI�$LM�O�ߧ_���)n��i��>n����SI�z��`|�Բ���M-���K
�{��\1�VΊw��PZ�vb��t� Sޙ�eq�����{���%P���.]��b�S"�&J�*el�x\f��m�pw<�
|��V�xe�A=�eFg�Fق� �M��7N�f�c��h
`,g��q(o?��*��p�J�J��$�'��Y�b�����&x=N���8!�P6SI����$�&���Kk	\�ō���3�>�v���މ�N�L���N����W�����}X7�֒�Y�O���So�����0��	���T,,I���8�<6nہ��^���^����&�IP��k�p�v�zJ,=��t%����Hɶv��c�4�#�W�6�8��@Uȧ��
��|��ȭ���CO� �ȓ�$�'�͂��Dĕ���(�b,�{`��a��r%�|���FF'��v8���l�������eZKN�����Ę�T�w�܉��6i�,��bt�:f�e@�WG/�Z��s����"��e]5��U� %Mʘ+�P�bg32���o(a��
ZjFC0 �^8�"�B����4�ŷ��<��;v��@߀ȉf2Y)���payyY�t��I9��%��<�U�BnWr�"b�8������᱇އrA�x� ;~G��N�<+Sv�f���N��/c�uR���C�Lǂ����?��P)���DrZ��$��ϋ+;;���ݒ�K}Z�����[�L�'æ����8m�՟t�4�'����06�;��@�>�臥 �3���x����ɧ�������bZN?M�1��7B`}�:����]��o6��	�;��ǇlbSO -��}�75����d3�D(_N�)�%�\�Db(�R2Q�Ϧ&'��A��/pY����&�q$���7�8u#7*����}}��}ב���{�7���?��q����Ó�}#Z6���.x��8]��ہC{�c��A4)SFqAePeuOMiJ�1b�vUL�XHE�J�у�%{��V�[�`�9�LW�0����
�V��p��z��A�-Mhlv�q)�afl#�#������ER\&�Lx�|R�ұ���mN'��*�zP��}{w�=��[֯�j���0��'ß��ghk����%x����&geˇ^�H@�flij������bm�.����fO��
��La~~��>�%�\�~�!��$sy��c��Εqmt'ߺ��˘�ZD�l��ŇΡ��}�;/T��!�) �)�=�b��Ǫ\�Xe)��^�!���E>��ra(&��M�|��Z��*���C5�\��A�H��pz`�AD�5���b2�o�1&�7IA�MC�&��+�?v\�ɤX�����؀vŭfص��j���S��L�H���ǿ�X
˫a�I�H�&e�h�c��ÂO��2ac�\3�b׋�����	�WϏ��$���h�$ҥ��S�ȓ�;�u�4�l�k�"D���/Ө���hp7��f"�͍��F1Oc" n���%�T�ł��c�RN��p;,�nmB_g�$c�J:L��gJ�3vk6'.�����02:!ʺ�M2*�����/�dԣWP�b��UQb�,�Ѥtg9Z>G��I�Y���S�Yk�j��,�Q(gau:WL���N�4Sړ	�U%�#�^��Hp���-AT��u>w=i�JQ�$�"�����]�F9���}�A�*�XJRhr�zA����%�=��1�� ��8�I�TfүQ?4�C�w�œ���*��C'k�V�-?���U�����M��/�p�uV(˛��l\׉��6�����D��jq#+b||sdrLX,����K��,�v��'R	�j�k��D�	%pO:&4�9��D[��X�p�aVWdXaqm`r_�O���ձI���)�ؿW$>�\&�0���1�)�f��MA�r��06	�ޤ���22��t�U�=	�c�0����}&_�P�)6_ʰctz	g.�`~E�x�o����#�c��	B!C��^������wo����au +��\�����eIV��=ر�_5
J�S6�$�P,�l�:�v��Fk8�1h��&*/�}�LQ��6�@�s�΍�.��"I
�W���pg���+�(�4U3ِM�D:�m3�����^�!���a�F^"��i��x�Ĉ�%Z������{�;��>����`xNo�� �8���	��W��G?�|�G�q�����������9��$Dy~&�A�(�╋XX���x�AI����Ec��v�	�ㄅk��	&�4\�=��o���H�`�T�8����'|ʑ�ٗP���2«�Or�}�b󦍈FC8�F����u�����%�ޞ~uͫ�hll~���H�hL�O�A����f0r�J#���L�Y��+��g��c����C9[��(��_{_��7p���f��A"5'���nç>��8x��{�U<�կ��ٳȦ�0[,h��(��3e���ø��z}b�7!nNg<T�S�,��|&M���J�q�f).n��i�I�,$�LOM`qq��_��_"P߄p$�o?��L��4���o�M��`^O���B�1��5�@�uȧ�M��"��P�5������
��s  ��*����꽴��k>M�Mżx��h���K�O��Jk�XGQ�\N}c~��W��-/�X��7������R����/����E��`o�Y#�]N�Nt�{�#�c�P3�f��i�~��#M�Iv:R� �)ae!"�*������9Oť��/��JY1���J�p�Ri$Rq�+9�7�aÖ>��86����q��65��\���$R˓0Ը�I�R�D6�S�)���.%����$R�{��}�#hooG����2=3#݄���e``��꤂f��BO&R�0�DɅ��Dss3::�D堩9��Nk!��	I��/c��$OT]R��!6=������!��K1�N`zn�ύ`lb^������R<#�4t�c��}(��OQȗoUD�X�V��6�	�(W1?:���`I'�4��B&� �C@%-�Cf3;�twUP en��.��h�dC��;qv��8d2P�����~5�b	Ԉ�5[0��*�!���B����
!W�S��ps��u���M�dsk1*�j�YTةgQ��v�LQ�H���)��)Yo�͓��ʝ�A����3A�"n��#�#2)�4��X�f>�THF�6�aM���������LHHٚA9,�XUY�#|3<n;~p9l"�⇄�|� ]�W#Q,�C���ɧ
���@WZ>���)��Y�d�h�B� ,x��u���1>�Ϗ�>lڴYK����&xYMa,&V�b�8N��.*S?���0�S"���*�L
1�Rqم�L��8	4����r(�ePٝ��������]qv���DH�ZH/��I�$R�@Wҡ7<�x��T�D
�|�MMqd���Ϗ�]��!|(��9��i:?A��L��G����[��25���CU���&�R\F$���*1���ˇ`�Id�+1+�4RK��2uRRlXׁu�:���/
���b�ӌ�����	��xvy�(U3�W�9,H��Hgk�;d���Eh6���n�$����4���4kk��~��Har��H�
(,��+8sqo��$r}�wl�ƀfC^��UY���N�A�2'�����|�ӭ�JB�&��J��u#z!�:��u�a;BbU�"�E�Ë��(�^����Y����qx �nGO�G�L|�]ÅKQg�a߮����B8���c��%k���܍���@�[�Q�O��Fo���Lϭ"Y�!���h��_�
��)��?B�y��ę���B$:)~PS2��0�*���S֍�"���\�BV`�TB!�>��b6��g�����J���e4�YXb�c�@�(}U���nkQ��*P��i����XRX��sWp��ψ���,�[Z�W������RB�t�*r�em��x����t8}�mqۍģ�箻������l�������я~$��=���$���$�I�f�)?j�{�`sX�07���l��o��fl|x��8(x/#�čݻw����O���.S1~}��ߕ�G��	Ŕ���ʵtw����]�l�Rxr��[g�g_��k��X���f
y�E�00Ё'{�>���F������s�.�I2+�ӕ��"�߉O|�q�߿SH�4Z�կ��}��v�k�$�G�gVIf�:��^/�˚���a�ҍ̈́(��9��K��O@�Z��kE��7!�V��c���``�G�Ŷ�۱��ɧ� ���p��4��&�k�F^k�R�R5���S"����ޝAq�����f>`����@�a�	�}���ҡy��)��)�B$L�/�+�zY/2)�{"&s�����D���N���rBOc�Jfmn�@��x��������!��^��O���ӡ�aw���Zf�r4Dk�j[;��#��s��tU�y�Qcg���7p��<��>'|�4[���!V��:9��ٴ�M��6�&�k�iL.�I�F��LR\\;�����!$�+�.cfb�Deh
	�w5��K��hne&#��xت�tCs��.x�#\�~�w�y�o? ҍ����я(c5�Ǚ䳂��}Z�����<��ч���$���[�lBOW�@�l�XX:B�Ț!:��&���N����8���XV�*�Vĕwdl
�/�#_��O��"�_�"U���І���x��͏L(�ɱW�x�M�=�Rd�bj�.���Z�$�"�,*Q����V23	NS����KB1�;5Jw�I&>�n��@Ȑ���w
����M��ۂ`vn^:U�ZY�!;�$#�.(Jr��+t��z�h	֣��>�C�޲��t��i���S�]K��;@D�+�XE�Ȍ��2r$1�*	��3a��T�@I�fg�U>Iv��xX�$	SC��k+�n��c7[��eEs%9��Ś�$��$5Ĩ��&Iz~�����Ex�4��]�\�T�dR�T�lV:ۚ����^'�,|N�V�����2)����0�W�8-��V�C�S} (�E��M�=ݦ6Ԇ�9���
A�d4�b$�<��J���_'�]�b&��fZ��
���8幭�����Ĥ�xQ>G���ia�HWS�1�	��ߪ/��.5����/ѓ�=vC�U��V�[ʱ���-�3��	W�$W�|e r�T��,�7IM0���]��p׭�wJ���߄	�Uu��F���E]I��\N�)m"�)e!���j�6���Z*Sa%+� Z�4�91�߂��&�fdk�Ob�֡\�`j"����XY�(7M�e�2�L�g�JS}Ë����J7%dRqx�fl[?�ގ&��@�i��Jq4��ڧ*����f3bi�G�1�ǹ�ゟg���݁��Vt���p�d�=�@"Y@���V(��LF%��ǫ��ب�b��O�M"�;v���UVi8��X�~��Ҹt}\x[$s�l�0�������,��$�før�
�=�c�V4)�XF,[���Wp��b�6bǖ����ˢV�Y֜TS	EҘ\�ڍy$�8�]BM    IDAT�0Z)�L�#-y�r�I9
��*����ݪ l����,��7S���`"�4�t.%M�5��шH��P����+/!��
�6i��r�6���Pn����40�R�!�x[M���#x��?�m[ש"�?������3��g��ć>�>��G��R/�%����Cb�c�zrb�7p��[�|�"ҹ>�����O�:Z��Z�V���/��^@,��{��&L���8	��LS���d���I�Y�3a���$����(��g>�)<��G�v�P*���˿�׾��$�w��R�S��۫�x)gY�	oCrX ���K_|
'��2���E�x����x��G���?��_,�����'��O~������OAh�H���Gp��^|��Gp睻�Hdp�̛x���091.����Q  )@ֿ��cr��?���c!����Vdn���K:DS5'T���d���F���{	$�f�R13K�*��������y�c0���/}�z�D�i���K!tJ�����zgS��	�-�K�y�o!�,bՙ!�F��Y|1܍
.D���VL�/SU��x���ffIG�PNFa����3P�g�1�$��1�&�E^��}R � �B��:���{>����;T�����ߏ>��J���� i*�TJ��-R�Y��c���.�}�\�x	�j{v��Jh_y�)�;Q~�T�����;cxp
i�����X�N+L�6kf2e��5������,2e�C�z������&�>u�r��0������`�T���G1����gQL��\��d�*�;�N&W<̫顙F����÷�Ё}(�3p9�����ի���3O�&!�^�AZ��6����(��j��B�����@�t��Q��`m������GTA���/��%��T��aq�(xaq�3�\ހ��G�Q��[��2��$��&��mD]k7���&�ǒ)��Y��|0Q�����5,^Gfv����"��a4s_P�J���P� ��@MѡYMY���bRV-R���#�Q���#��ӽ{�<� ��XX\{s#Db�U��;V4�'�y��8'A��b�]�A��aag�p-_��4�%��C�hD<�)J(����������t蕻����ٱr�35�.��92V�Lu�u��l����tb����N$�n��+:۪�t+F�	&1�"Qk���I��C2�����$�|�(���j�Tu�'�.��ь��4xB$ʟR��ԍ��$���5Xqq|Y:��BQT��E��3�6��r*Մ��L�����$k�\�v��;1�ó�cg��v$�xv��I�%!R����R��$Q�8i>����ȸL�o%Q��ўUST�F�On�GhE�~ 	wA3y�� �%����4����	8}n)�0@>���H�c��⇒�c�QM*t�J�0�R�
iPS�R��oeQ��a\�L+7Er�d 	�s)�b�����Z�	z� �LJ��[~@8L6��"M�x:� 0Vjp�-���@w3Z��i@&F�UМ�$k��
a~6�|��σ�&�@``-���{����0��WV�8��I�=v�ݶ�*���L!�2�R+���B��U�	�R�B�+�Z��j�X
>����a��"y�$Le3�*ɲ4o�	f�kN�jf��&��:g�A��ɁQ��!
O��_�V�&����_��Ĝ@ٲ��n؀#� 賋�%u�/�-�¥�k��;����ʖ�8w�N����Zv��� n۵�=m���
���b���,�8w������5
���1˒��!*)��X�]Y�U�`�O�x��5l8XlF$S1$3q��ɕM�,Khh{K�Jo����'a$�����J38%#IL���j@�{�FZ�Sµ�C���ģ8�o�d�L���p���p}�4��h�����L�DK��W2�M"��\�g;�@��%�����H�{�{/�˟��:�d]%�i�8~_y�@��Z���Wj��T���X4�HL(%'KN)���b��t����Jgd����9�ݻW&��R'O���'����Il߾]x�����E����P<�섳111��}�Y���)��Q5Y
OG�P������c���=#b�<^>~/��g�pq�f���B�E�wܾ{�Ql�0�����_���2����|a~�{9z�Rr���I��)��:z�87���	x�>y^z��'�z�;�K����,�dƶ�4���f&'�c�n���/زu7^�����~�H$#�sy��J ȧj�*gu6'!$��V�
�ќ4�U#�?�f� �{�+8<~x��a���h�k��>�,�J��j����W���J#Y��>�H�L�lV�/h��?�[�i�7�[M�K�4J���Pw��>x���N��c[����I��]��(�kȗ��X��f��fF:���˂�� ���n�$����ۿ��(�p��d���C��w�%� c�R�N�F� �{&R�XF(U��\c�i,�ʈ��9�v�f� _�b-r�`� r�8�]��ř	��!4�,@:���K0��2!��h.pX��%��j������܉-��1;5���i�w�������҈����{���tTĠ��.Gmbl$�N�9Ew�*1%�R�(���[����$����䏋���<ߗ���L&"���M�|���P�.����q�r$�91�A"���,��Xe�M=�a�>��E3HĳHf����5`����8४N2���iD�gQX^B-A-�TÀ)-ң,�b��7���UH(��	F�Qk�`팊U�8�z� pl0���m߄w|�!�|.��	���9�fAŮnUU��pJ2$um�q�$�Cr�͂&�5��Q��c$݈��3��	Cz�����%�`��Z*��Y:3�Dn�$$�o�T �]�l���y�D�\�:H�s-����ʁ̓KW�aA�u�D�K��$!2�Xt��=�{}�`�n&��Y4�.���'YD#|�Y��q�$�T]��8�g;��(f8���廬���0��^�'R�⺴��]�ʊG��g�C��6x^7'1�mUj,�TrR&ԫZFP��*�4�E�U��f1�q0����3r�W�@T|�	3`�����
._��J�\	�� ��D.�k��%�*t�֭��>!��f��w��u~L����ؘ$�A����F�E������XF�5!?	���aГ0�c&Zͳ��$M?,�^Vk"� ��̥&Jc^�\za�s��p�V����n��	��l�Oe� +#'�=�}�"�uv����WP�|Zby�d@"������V����׃M[��UdKE*%,�$qedc�+�:<����f���я�[�a�#k��jLU�Y�k�Fv�Ua�j,&���ˡF�q���� ����������I�$J���-Nl!r�b>�N%��%#,E��o*�M����`|�l8�	A�i)HN4�D�3U0����D5��%�عu+�q�>)�f5m{��^z�%��1���Ac�W�<B��}	���(���QY5����"����h��	�p �+��K7�!_�?�f�Dk;������%e�:���V�ʤ�e$ɂ�j��jn��bq���YX�5x����#�"�Jh"9�`A >���b�Â�J����%�}�A��;���H6W���������Hz66��Ԁ��.�^'k<���4�>(��	���r��H�dO������������X��/���B��_�?��'���.qTȱ.���<s�7���%RP�����$r��(���/p-楓Rtuw�����7r:쒛HAp����{��|�::��#����Bdry)fX��wv�qh������q��P�nQ�aA��݂?|�1|�#@�P�"2�*��'������W&P(�Y�,�\���A|���Q�����c\�r��:��e�ຽz�\'?���?jڠ����yJ�x^r!�g�p��>_+�q��S�Wb��i��FĘ+��<���D���M����p�{Dh-��_9��(l.��%�Pr��3^R	R��y��'<����M�, p���oE���� �yzXQ���v��0 6��\L'Q)$Q.)�+*c^�K�걛��N�l�kh���@�R@%�6����o}`�O?}���S��������_O²��Ԅ�YL&��~���L,���l6���{�/^���|T0��Y4��}�>ܶs;|8I4dG����i�A��	�\L`t6��ł��>Z�`5H''�M���[6uS��]��Kg_�BS�	K6���8��E��7�`�T��#��@P ɡa7a���رu3V��E���С�ص{����|W6�ء�7�d���~>���2�g��>'tG�4�I!��t=��W�(}��ZX�gu9$h׎ݢ�R�"���c'p���0�=0����#��A�lB2W�b$�ƮA�o���E8�N!��ưP]��v3�n;�6
��'f�� �V�| ��F�A#�b��M̂�Xm�������vjf�W��@
��d���q�R����]�:�t�s�tIEI�0��D�&���4����C��`��uU\�]�smfS�G P'�ⴡg�Y���(�t�I4I��lN �BF,W�S���aI�v�]�v� �q�`0<T�#\)���L"1�L�x(���_��Xt��n�HP�O.��"Q)�8�11ɏ#�%�,ȃ`w���Y��ES��,v�J������؄Z~��M����E��.<3�v���d09�/ٰ��e @�2�b���F�3U�t8�t�4wT�C�j�M��X����	7W��O��TOqK�!�hqu�t�!܁b�[N
~��	D�Yx}A�NK�"�Q�	!�P��֤[����ū��H��>���q��~��v���g��U�^`)��t�nr��4�8d~�I�ӻQ�$A�\�E�t�Y s���,�J����?�E�/��)�+��D�k���I�E:�2ANg�PŧS&4�BNK]m�6���C� FY�l	�3��A$G��Q�?���j*J,�D��\g�\��|
�:̄������{�m�@�O�.Hϥ��F���OL�=�3��Xe����kYL΅D4��a&�=�ص�M�����-SńqIA/v>�Ћ~�
�χ\$��>{Q�8�>�	9G\�*?�Z�lH��*��n`jn�B	[7o���[�s��zʕ*���i!iڻ�n���*�-���z�$^?y-m]h��9g��B������@w;���t�X�"������Q�4�G�L[�x�3�:�\q�Sc����Ҫ}��9�=NPѫZ�Љ��&x�lk� kkaL�c>���%�&��aw��8GwUY�
'DL��me>@j����n��~�|�?<���Q� �?��/�W���C�`�{���ߏ��V9Wɩc�X)�(hJ"<�LJ�I���G�m!��}����?Cog�@C�>s����o��8�e�V����|&�.]���֭���"x"8{�N�<��Z;v���M��at��y,.�cÆ���R��+e�:uO=�N�:��"������4x��(	Gcr��t�a��M�Y>����wp��(�%�L�yru�����x�>t
����������!.\�&'�|�)����m�.ix�u��ˈ�W��l�s�M:��˧ϠopH�<�������E�n5���Ƥ�ω������o'581VE�ݽ���mS�w���آ���j�i�p+N����oC��p՚�tFd�)��u�lZ�A�!�ߌ�5�ݘ��o���M���&b�����:�5�#K`ee&��� \M�8](��Ȗ+�B6��&&��'���Hi�y8m�wC���^��8#�����Z^;����lN�.���
��Ԗ�ݟ}�{~�ٻ�d�.����wS��wN��篿�L�j��l�'���I�X��b��hڐL��m{p��Gp��9}�i����u�M�loŝ�nGO[\v3�4qXa�*WE'�H����lW'c�K#5�dpIA@�aq�#~��~������+W1r��Ut7z`�&�<q	��)Ԩ�c�Tr�Z׌֦V����dri3��;�o��X��ĸ$�w��Nq"��ȏ�C��kmkFWg����"�i����v�qR�����i���XL��(b MV�@ilB�
��vm߅]�v���M
�_�t\��*��V��C�bez8�۾�v`)�A*gD4U@.S��<�&-6�U�k��1D痑^ZDum(D�R(� ��	9Qg�8X�j$��:�]�����q;�YgA@Q`*vX��,�jD;�J����;����G�Ey�ȟA�;�l��ž4�A,�I�0��L��CbJ��}"[�d�N�7���UU��Ē&�����
���+Ja��Q��/	";�<��ꋺ����d4�/Ovcu7G�#��R`�����.3�%Jk���@�F�@��H\=���N�T��Mf��0�#	gs�b\������nd�K�1��9�$��*{W��r�R)r�jE&CGV-���m@b���U9���81�5O�����p(.u�Y����nB:�(���+��e�D��ؔRa�[4�& ��Vp��Y��py�ů������&���֮���$>;~>v��?�������F���nJ�Z�vy�GT�DTV�DDi��(� �����~
��_�$q����ݚ���k�n�^���:��V��^��A<E"�{wg:�Z�2�{�n���p2Wʣ�O"�b�`{�`5�d���I�Ǳ�1�298شe3�&�44��01���ό!� �ƀ�!����ni��MC�mi��Z���"�뀜��481)�J��If�(�������arn�Qd�8,tb�^4x,�
��:d�A�J��!���m�
�Z%���
�;)σ�����XD(ia:�R�\H/Z�L��*2E~6�*nL-����^�lZ�����r;��p��eї߻ewܶS|R��ȕL��{WF��c���Dts������z�]����ND35�X�����1�����b��@k��Zԓ.�J�<:4T�Lo�֘��P��:�7k�67�pS�~���L޸�lZ C��y�e��,\Y((Y�2���]���h��{�a|�Æ��g[_x����~A�\�=�h�lXMoϠ���e��T�;���}�)�(ɥS"Б��ݎw����C_W��}��I)�Z`�:04����~���yG1
���7������k�n��V�?���7���] x���{E��d����J'�+_��l�BgTKe���x�O�T���X���.EC{�2:�c�Y\^�u��ٻo�pΞ����~c�pz`��NƑ��14ԅ?|�q|���%�4����_9&PB�ss����y6q��q��mۄٹI\�rN��Y��y#Jj��wzb����/=N���
J����<xPރ~To�qR��5���).����M�CP��H���E#IF d�fS�C4�@!_E[{/��zē9��/E�ٶ�����Ć�u��=oF�]N(���k��_����9X<�0��}���8|��������b�F8M(�(��"�J����]w@2��\���x4������hn
�I!���	��#��4��f�����#��2:���
O�Q�ҹxlz����>q������T$�������o����/}��o�Kƍ��z�̪+��A�:.�\
�M�X?<(���	����������'1Ms�G��[6��ÇD�i6�=X�z��}=�8��fE�FW��^[ƕ�(R,��`'#���蓴aur�R�ьx4���9��O�i*���S:��k�[G��T�����Jx]~Y�\�R��-��jÎ���a~vZ�-��.�*8u����I	@�䲛��"'%���hkMbnn Ը�uB����+���߹)[�� Z]Z���,B�Q_ZB��uuX�~#vl�%Z�WGn�d�!�7at|��O#����D����<    IDAT�ܴ�k��a�!iW��55%��F��G%�G>�Dry��
��y���!�*qR�a2��H7ْ��@kK2���&d&l�$��CUMjb�n,��m�َw<� �u,���c'#m�N�e(Juꄛe��H�	��("��)�aU;�,��1����]pk�;�4����#$���?t]��nu��ɩ�|�K&�Kͪ\O�T⯺�1Ѻ$z2�]=qf�eW�E&��k�ȣ�M��&vQ�e�seKT�����>��Y���y�R���Z!AOafy�ʕ�\R�3U�l�յ(����SEp�3����,.���pJ7��{�'��-IK��Eau�t�h>���=Q	*� Tn��� ����*P�h�]��tlI{|�ʮ^ܞU�MDi�j�]�c�B��E��B.��>��g1�<�(DF}�t�Xq��].)8bVE��ܳC-
lhhR���ov�4���n��?kdh�P�z�u�/ Gl�2�ѧS�f�N_��� �$��f':ۻ���$Ϛ
N$��J<+��^�����uaˆ~����ͷ�8�d����`�$����05��k��ǫH8͍�`, ౢ=�ǆ�Nt5��m��e1�KgYq���Jԕj���,X�ep���O�a1s&&���mط}:�0����P̪�,8}�T]k�x��eW),{Oa�E٥�T�xn	�S�@��JG&�B�)O3�����5��ӗr�y����؍��)���J"+q��)���6�Z�T�����2���u�$ߕb�Ks�v�
R�U�{h����z�7R8u�:�V�R$��l�PQJq��"!��9.���N�6��&�Z���G�D)��K�}#aU&3(���4+��~��Jg�8��ܼ�>��oN)���[���N�<+N���6W8rh��3����I�}�?�7��.V��u2����@��L<	C�$��V����T��P������H��k�������>��;�h�p���������ŋ�8r�J#1&�w:(��k��*S�|P<��I濳	Z^���E��M�S���s�}�1>�g�}��:)�a��~;,f��o^~�e<��S�Lfy�|_N	�:;TN��$F��ǜ� 44a���9�m��Π��N��L�b����?x��>X���%�*#���y�ΏHA@�L����t��������!2֬ژ<3��W�ɸ�^3��G�ϒ�DP]M�@��䡇�&��~�3;���Zi��G/�>����dG/~��l:��&d���xͦ�Z(
����/	wR���ط/����c��}hj�A�xI�����<0:6���;.|J��K��{��'�����?����#�<l� 
7*�L9�HG��x��;�G�� �2~���ӟ��+x���§>�0Z�}s���X�ʄ��B����2�<s��<-�.J�%�iMn[��W��]?y��aus����
��={b���~�L�b�`�סfQ
�L.�S�9Lvoۄ�>�!�ש(u�ө^�ɿ�؉c���]o6���Eo{'\6���%��-(,H�Lx��x��l�nx��RX���g�ჃR�F�yqt%�+#�C�߆j,����]�����f,�Nɏ&����C�K[{Z����D�\BGg+n߿G�+.]8�K�/`uuN�CF��L��l�B1/���� ��RE�&
����4�W%�c7{ppP>5�~m5$cS�y�=Ĭ��7��=|u�B(Es�|m�ώ �*#Q 
5��Cؾ��e��Z�p�`�7��1��aV�w��=��9s�7f�M@��(V+��c�5�)�)�yM�ww���11�1�^�DT@Q@Pzg�齜^߽���$��~����s]s���|˧�ŋt>�D��-�䎦_�GZ��t��fezQ`� ӫ� H���E
�B�\op����\�jѱ��T�FQ��O��\(7����`��8��ᭈ����=���$[�
�$i�R�g��*����|a"`W��u��y/�$u �9W�G0v[���$�Х��d�ϧ	+u k1�شu�I���v�CJdv�17'h	�7�{�^�[��"<��6�.�Lz��U�:�Ҍ��.u�V��c@����֩Md`(!�7�5r��&�~d3q�5fM����R��.��\ �Kt�t

�����t���\����\Y�ѯA]C��ג/$L��J-Z:P�}�\�y���b(Jb�ۜ���Ak]�=�й�p�+��fUi�s!_�2�� q�@W� Z;��s�A�u���	��+�0�.K�Z�����݉�:�gc�7%8.ڎ5���]�s4��&��_��r��#�
?��T�%��|�"A�����
��`�bÈ��X�Fɀ�����J�D�t�x�Dh���l�!n�x�6ـ'�ƺzT�W(�Kfb"�˞�8<vo�)u�؈i'����zHKU, �0�i�%�'�<a0$�m"]��mؾ�	mm����EA�*��Tct]9�"{�tj�1�dB��'�L�~C���ۍ��4v�>�]�����5��][V��N���'��;���DN�	 �j�߼,��0l��N]@9iS��T�͹ynm�\�ةS��D4|��6�Y��$v��4	s��D]enG�x�$��F�u����?�e�Ł�G1�|�2c<�4r���9®ql�SF�@eU�L�z��΃ز� ���9���@���O�ĩ�%�T�}����C�" {��a�@r+Ut��EK�Q$�QIZV����I`˺u�;v4�Б�db�+/�D\&���S�E��&f8����ÙsN�������6�xk1�����(b܄�8�$$3Yu��4���0�����U��t�x�a?��v\s�%z��ظy}�����2�cR��p�5W��K/�����K���?��R<����oo��6x�>�����/����p�5��x�� v�G��#?�1,X E�t2�e˖�OO=��7J�K*>U����|�&r2�7Я�����Ĕi��}�װn��pKPR^�U²1�Y���7\~��O꽽�x�õx�/oc�'[���=F"5��"\�'tc��E.��~��z�1,�0�hko5\(KZ�S��1�}O�~��ș<묳0f�|��g�r�J�1��R�B�1�2�U�_�-�`�44�3�8��ᷱ �9�vQ��.�Q���{.n��Vuw�g�%[�`8(�f0��`0�ؾK�.úu�Ȼ"����+���c���Б.,|�m�ٰ��<�$t��������.�O~t���n��/���{�����ŷ�v��
�B�Yr�ƺ�|�������_`���q��N��m�'�ix���^��.3������XB��?�{γ��x2�NpV�b�倏��
Y��N�?o���<D�h=rjkQS���^�ڻ�����"b�$|� jʫ1n�8=$:.�T��������V����M��;��F��v���K	�7�iW2�q:P	���G���|��/�d�14�ڂL�!�"ʎ:h��r u��|4��NdVV��oP��|g̨��0q,F6Ԫ��*�G����[��-9�(R
��#)�P�'a�ԥNK�[�ߑ�@%
�H,fRB>_�P3HĢP;��}n:t�t��v�:o�ZП|��7lG31߱<vjA�/����8㼋�F�7��@4��aFޏZ&�!!�g��jjF����v4�(7�B������!("\�@�=!��X�lĽ2D�c���2K�u��/0Q �?C��^&�>�z-�5J�H�R�M��8)�X����dF�*�q�%N�/��U.2A�$ٵ'e$+Kը\&�"b���2q"f�<��w����ު*�����9�܈s9%w�(d6O���]:�T�M�"I�,>�Q�a�c��.`���c�MU�Fq��Q�u���@�x����9�w2YJ�L��֖"9��~�
��TT�,@�!Ǭ^N�؀j��К�(��i9<��8�30dK�YX�X]��_8NH�&T��1;�d� 3(q(�7�\,��� �1q�3ƢHgG�:rL�i�N�b.YEe@�{��R4���H�L�$��W�ΊH��y΁�(��&���A�-*uP�TJ�c'6��S�g��o����6tmQ���_E�	⡋�*a����s\�Q�	���E^��_���ء���q�v��4��Y�U�>���������GRw:��I1׶�z(�.�3q%w�s�j�y�21xYU�G�V����%$V�	�
R�"'ճ���aAN�������%��חBM�(�Y5��",חQ]����\n�CJ]�x����X2��Ã��!�>x����g�xs��2!<��=c*B�F�Ѩ���8���t�l���L���K�X+X��`�Ɲ����s��H�qʘ
z�"�v�Q�q�m�"����`޹s0a�з(���Օ]�t� �C1������f�g�'1��1�Ա2MerN9a�s$I[�&vJ��2ز���9���#����	�v�dD&/*�~�~�֍��5��}!��7�s�aw���^89:���H���ի1�|L�h"�s�"�_��NnV�UXrt���r��?�^�~�t������S/b ��/�x��)�>�ƴ7;΀��\�D
ϐ�~��)�f�=*�F���}�߄;n�I�i���ٍ�=�8�Y���p�ӧO�5W_)u��-ë�.DIq1~��7JJK�ǟ�����5N��_�[6}���G�妛�����?�0��.��\;�o�~�Y%)*�x�����ʐm��N-yJ�H��!�_%���p:X������s|�H2� �)�F���݉��_�b�2�������E��H.�]u��j�1y�D���n�X���\>�ѣ�h��r��~輸���u��y�X��F���,����w�w���E��e��9���8BQX*O���jOe� �I�!I�k�r���е�uc��x�Gp��sU�!��϶��ہ��J"a%`#Ga��PQ����;���/a�*&\wõ��k�b��jm���z�����t�^�±�^uؐ�Ó��K��_�_�탵�����`���[�ݯ�����$:{z���k�e윳h�0{IMm�޿�%�%���5��wp(��ӳg⨺���w.���)ƍ���K���,|k�_d�#F�a\{�,B�"ԕ�p��q�Eg"pc��!�?�3�����*�2Tx``�'SR�8��e%���n�\4|~�iII��z���ջ���f�ODq��u���E�U	qU������O��D?{Z�G
}M�qt�f��� B�D�>%'	?�GPY^	���r^Iq2K�>c*Ə������P	#�R�p��wD&bfzƙ�c(��"1�|�S�L|H�%�6� &�ڋ��}�Ed�	��!�D�pw:P^Vf*�4���W�ISNA�P6���k6c �CK[?>�b/�i/������Wq����s�I.����@\-e�X�*�f�{�=MMH���(7g�_vB &y:�Qe�ݖ�������Q(�&#:���9����7]}]D�$�ǉ	�OǼ[�A��ݽ=����j2��
���S����Y����[4�!U�YэU3�F2��	cF���]�8r��?��e�B^,B�-%Kx�ԂU��hr�����!gGBH!C��Tt��8h��@2���Γ�g�<�;�diΠ�����vttu6����\yZ$F,1����`D�U*=��Q�r��[h.>W6��U%a��B2u����LZ2��bȩ�{ &�&%� ��Ta�G(EA���)B�@G���I�aV�����/XQ*���k%���B�4K�N�3�y0�crH�ʌ�P$JݕJ�L�e��ބ#�*�����%y�����qs��o}$�5Sw������U�;-3��\���n�O\(*ѯ��g9�Z�Xv���d j' ��Z���$c��'�j��7�.�������=Nҹ������*kQL����	d�rHfd��rr���lg
~���2�Gף����2��f�����;���4j��574u��/v���PUW�4	��"��x	�1���U%p�#!6(yf�ǃpq~�SN��Y��ȣ�c ���F��@,�?����ȍ��:i<��	��t	\�"�,9M���wX�f�Ɓ��<&{�/(��j�̦

j�5f�)�ۇh��G;����%��J��3fOWB��*��t�D�T�@�2�<7l܎��j�t�$�1{&��ڒ�7�%�K��B��I*&\h��Jő
����c��	�3���YDbv+	�J%FVB��N(�a�.�����̲'���b/b�=X�r���p�����!�A�d@��1��k�,�PȀέS�^rz�n�<m��5�O=�2}�	i���b��q�6c:&N�,��ۿ4�X�huE��ȋ�������)�����rӵ���������;��?�o��5u|.��B�v��hQ�O?�K���]�w����������3�>��`��s��������[�!���E~�W��t����~#j��Y�Ze��!`q��q��;_@�[��*��;&�s�Y��U��=x�/˰��5����w�ܤq�q������A@�mSx\��'x�7�i�.��͈��R
#0m�I������(*��<��)��FiY���m_�Chǎ\��tW7�����)�3g��D�k���KLr��M]8��5�T�M7��Z&z,�x<:J���l65,a�99s�P�1i:�/�/8WEe�W���~� �S�ǥ�C����\�y�͗��+/���T1醛o�e�jqY<М��n�����c�B0��ʦq������X�����3O���&��=���w �b�֝X��:�޻Q��d�����q��K`����{�m{����E���xl��ɣ��ew���J���K��t����F����\\����F'����\��3�q�N���;?�W\p!F����eB�VŌx<�C[K/z{��8�(�Hz��!Q�v�1#�H����~v�v��zxH*�2A���A�Ji�GIꮀD��8z�ñ=[��k���Rz�" J������b��jkkPR�IS�b�sQW[��Q	��r�?ڋ��v��S�i��ʤY�`�g3�G�����_�v��S�NU����s�pQe�L����H8,fyYDb���G��8�/V�r9��x%c�cO3>ٸ����i��YsQ=j<��b�F�2��F(8�������2I�t*�:vm��=�(�$��S�|΢�����@g��^Ɯ,/Q{j��]�f�������)�$��4�J �� F�N���n\�p]z��?��Ŗmᒯʘ?�L��:�t3&����~�eśDV�T�Mݐ���R� ��Ϗ!�@��z�,�{C\D��{��+�
AuE��|@��nu����ݣŐ�q>c��y��S�!���=^Ub��Q֛.�Ȳ�aHX2�	C�c�`��y=���<	�߻]~x�AU��]p��x�'\$G�����j�D"�-�H �u"R�s�C�qYvz�p{���4���JN��i<I�Ӏ������Xu2�Ξn�r"%e��ciU��0at���) R+��$Lg�:��P/�5�bDukx}!���5+�nNj&Z&d�@�4n'
�E�:ɠ���|3A�1X�v��ft���܈�--7	�)y-v���i6L�p׵��U��{�^c��of+?ِ&\O���i�7UL�I�浘N��ü�%e���C�/ Ln<�Y��yMX�#�F���|��,��0fT=B�^�������#�Σ��[�Hi%2�v�ڇ�NzP�8$gp���1�b��b�6Tc��Fh��(���X�˰/ ,���w��������7��*RP�V�@�T�ǎa��\6�p�O���{ى�:�Y�(����    IDAT���Y�Yj�p��^�&�0&�^��k-qA�#�/�.t���������^t�j,�scҤ1h��R'%t"��#����D��׻�����ӏ��A�W�a��31s���=�O�P7��9���Cq�W��o<�e��c0�A��т�1Ȕc:;\��0yV�2�Ŀv��^a:bL��{��N�'�Q�&�*7%�VQ@>>������c���s`�˱Τ��y�8��&���q:��W�+.��o<x7&O#�\.�g�y���o3��bǽ��F"
���5I��\�B�����Te��I��v�C�PS����\q�$��|��#���?��wi�~���n������k/c�͒Kn�����C�Y�.|]�·�z+��C��/~�-�6㡇��;o��֭���'�섀����)%A�����5� $@ۿ'N��S�}��A� �WV��Z&�1�'aΜ�ߗ�o,���#�}��E2G��´ic�oݏ�Ν+u�|:'.ي���O>'	`vrY���"�oĈzL�:}��رs+b��]��O�v�[�~�}���^���-�� fd���K�K]c3�(�����b��dix}|缺�4�"��]k븜�<%eY�g��?�k`�܌ع.򠺺�dZ���/�?���sѢ7�b�*��ׄ���Hˋ��TS3<͹s��Ysσ���G�?���7��}�M���;n���#U$1��g;������]���������ȏ�߽�b�|�i=ւ���*�}�}kyk�j���8xL1@oO��-�w~�n\}�h[�����X���xkkˮ����ӂ�.]����7z�����X��G_Z��;������2#����btC�?o6.��L������Oa��-�j�Ÿ�����<��ŗ8�Ԅ`I��R��E�(�8b ER�$7u�0�zB���r�A�޴�B)�rd3��%g8/I�I�bR�*��Kc��,��=�q�P��.t�u�(P &ԘI1[#�EYi*+�d�#~�<mο�L�X�^��U��6�߃];�	;��Ձ��#��NGb���ɉ���a<&]v���UY]eE��ww�6{b��h��F��P0�Gf�#Ǣ�v�&;�c�E�Pɬ�����Ŗ�-(1	��R��C���P"��Z�sVL����g�2�n>������v�ri��g�LaBN�NG�"r%�)��g��R����Ħ��R�HT����j.a>�2�4�^�t�G͘���e�58�z�dBA�L��������C�CQ���S ����i��T}�@���(�Γ�7U>?.��"p�e4j��~� iY�E�l�KyPXDs�ba�ǒ�����*D�ڂ�6�^'�2���%�����g�RI�3�������H��f�I�Ɋ1I1ĉLLs�Im*1���N��X�Pe%!H*�l�{x�Ib���=��Gӱf%-��18��k� g�`�#;6|�5TuVp.��y��X�WBg��=,4ϟ.ڄ*ף���a !����<���!�"j��Qo*�v��3yB�2BGh�dt�D�3n͇i���4_�U���t)��%�nw�o%KKl5ո,��0�8���^��m�$���Q�:�Q�����ߣ�;�t�0X���(�K"U��kkQWc�'�S�X<���
"7L�����y�3!�6\F�PK%v<��(��Գ9�Ҋ��A�B����\ԍ7�BAƏGI�gL$��_�)Hb�a�~�k ���VD����W		��$�t���8PUA]m9�K#���/���f&�y�TUk}�z��ծ{��߮��C�t�СC8|���&��)+�%W(B[W7��܍M͈%h>H���G�et�e��Uե�(���-J}F��hk����G�嶹FcF�Ĕ)���Ơ��A��U�<�� rL$�|��d�5�q}4��/iU9Uҏ/�&����*iS[��v���� ߟJ��P@y�'��OV�Dǁ�J��y��:��PH��.���f������]����&���2��/.ģ���:-��74���3f���L
�2�0K�&�LG��&�^V\�y�=H�⨮(���_�[n��U�2�\�z-��o���u���U������_l�/<��G���~��I���G$�SN���s�UW)���/ŦO?÷�.n��6lٲ�?�8v�ޭB�7���q�R.����ēO>���ujx�5�5!�q ʣ&�TQ��$>���Q�8v&i'^[�6}��'hd<1�\Q�����߸��;�Tao1���X��JA�v�9"�	�W|F|>L�Ə�.�00أ���-��Q���@�,�1�F���g��X~<V'��k`��&"�Ѓ����@�z)��Nv�G��6I�!Q����"�������3$\,�q!�Ȣ,R�s[g3���Z�������o��^~�u��Ӥ=�<Er\ȓbу�4ʑ��6���#I���=E����p�MWcTC5\��zء����>���G�6Cgw�܈/��l<��;�K�d�[x��g��Ջ���*��^�l,|�,Z�>��oFt ���r)�5��1q�X<p��pɥ#�.��V|�.��Ѻ}��~�����o��o�K������t��N�ت������U[&��9瞁�7֭ߥ�����V\q��زy��mm���?P��Í�#�b�gb�8�ט`0L��&���z>�D"|��Q|��n���ȻK��+�nBS�z0��RwݕGmU5�%8��K|���p�S����k�6 5 O�!'8��L���GK�JDJ�5��%~̚=	s�9��p�#jQ!�²�����/ɸ�D��a[&
�\c��9��Ĳ�ʿ-+��fdOy͚8Ɍ���#����F_o7��f�z&"�:U
iڇS�2��hɼ͝i,|�c|�n��#���#(wL�;$�-�^�=-��s+�D�A�#�Ews��E��.U�(3J5�+�S�!���%6�[��9�h	�͆�1�}�*_.+ $�E��#��g��+n���bh;�!+�,�kHL�.�L�3�pV�Ւ�$-�J�=�%�uq�P�gt�,z�ɸ!9)He��V0A�u2�����(�Ӹh�:��"���Ua�2��
��uJ��M��j]_ow7b��8*��LAM�C1�s:�����P��Ug&gLv"\�zg�Y��	k�ګ$u�3!��\��Y�i�КV��Dc���}.���z)��E���lZ�AIq@U殞~A�5�3�ii��0��$;c�}�k���=��zU����cI��5J�	���c��I�Kx�BV�H���Lʟe���������Ҟ& ��0�L6a����G!�$]ָaJ�:8	tS���݃��V%��0!`�$ZVD���t1AR�eU���&�am�Xl�]{�9|��Ֆ�'�Ƽ�Lh��pT�5��DƓ��-�0��cѡ�CŒ)�?�F�:�uͼ��������=g`W0n�J�s�P7�fYY�J����&:�c�W�=��O�|&�H��U�S��CF݃DV���n����,#1�vj�����ćןQe��bq�~�� ?��bP�
@UUN>�d%I��=�zL�d���L����V����"(�q���Q��
�Cq����8������7�y�)y0g���(՞���wt��څx��
�}Z�,�#�
�=��Bn�ݿG\�X���PG�$�|�n�!���G��/�;`'z�'��+'������T�x��楀�Õ� /��B�vlX��H�$㲘�΄�ݪ�K=�	����g0��]�������1i�hK*��_\������� mD�H�4u���]�h:pP�T�^1�zV�@_�҈"0�#l�	AMYw�rn��F��b$�����գ�|�稩��w��)�:�k?Z���v�С�
D��w0n�x|��F��3T������7��M�y��`<��SR
x=��O�o�Q��D<��{A�#�	�����`�6����͊{�{^ZZ�{ZW݈Q��~���ؾk?ମd��&Li���W̟����B� �,[�7�y_l?�������*!�z��y���C"9 H;�,��Ք����C0"r�\9�U a����xب�}D:�oM�m
&�N���ğI�k�&���!�5��㜹g��SNA$Bkg6~��>��n$r)�[�
m��h����.��~���)6��������a뗻147�@��r��ޗM"��^>4z#�?Eyy	|�^�z�(2� �2�Ǐ�t�����>��m��K��e���}�+(d2X�x1�y�Y���ᡇ��w�"������o���}m�YϦ��t��U@���յx���q�U�!�,^�:�G??������~��UB��/_����U�wx}�).�1zD5�̜�3N��Q�%8tl�<�:�X�&&M����N=	�/��O<)�|�[��$I�4��aܨi�(����)�$�t��/{���8ؑBA�e�xY��u���q���T�	z��Eˡ={�m9��V!�ӌ���4�I�J�j6%HK"��Cj�Qnt��I�}�t�Y�@?R��M�V,|�%|��G�(-��ֈ�Z�$����=����a��\V�G�#�(��`X_>�2m�ɓP_נ
W����Ac�(̘9(
����T��^�{L`㊠�+��Wl�K7�wЏ`���LQ�''՜�$k
��EZ���09Ȧ��|=�Y	A�xB@��<rE��4ظh��U�%�_US٥BMA�L�k��y� ��>xp���p��� A'��#�$��$7.>$�2�bB��,1�����$s�_a�Il���� ������� E�-�MYMG�	aF܌X9�h�G27^�����Nt��j�3f����5��`ժO�Ŷ���WTWicf�MFB�A(���r[�T����p��i*�F�ԉL�R#�H-gS}grgP��l`P��0�<?�u8f��»��!w^7y���87q��h��(�if�͘|�Lk�1�7]�����K!��um�yH���E��7�t2W:1�9��6URE="�9%6C�
S%�3$&$�2���/�;�~�Wk��::�dJ�S$����"Q[�y�Hp�~lL������[��Ц�ꮁ�0	_��.+�sg'v'ȾO$-��'JڪAQn��eJD%�2�YY>[ӕ�.�;P�J�e�=�� %)=k |L򕔐6d�f�9r�x0�KC���y�WN�OFL�LrXU���}�01v��"�d٩"������D���r"<�%��w"�a`pHssܸ�2Xڵk�B:�V��R[
�Xq��B*_ 	�L�2?�b4��B"���<�`��ys,0GzO&M���Ic��f�{�^��H���4{�Pz9�`'2+.޿}�ʸ(����B*�p���ʽ����0irM��3ɲ�x/-�!K��N(�!N���'F�+�#�.�^�|^x�r����܄M�V#��
�׃�0	�"�q4�`I���6v���p��W�_��&�T����W�ģ��
�xe���:�7A�u��-�J�z{��	\(il�5WL��18�+U�ڪR�}������0r�X���W�VB���M���p�M������e�E����_��G�HU���/GgW�>��֭_��Þ]�q��はݯ���o��g�U ��_��\r��8ag/���{�y�up��	���:�qk�g��g�1M�f&�#�cD�8ttG�j��=|�AJp�0D�^��ķ�s?\x����=�%+>��o��O7�@����R���&�<e�8��=��5��G�9��Y��䰲�B�f� ��ڬ"ϕ�K�>#=���{����������R8cܡy����W��ܿ��q�����K�p���������������]����j�|�t|���@I[��$��/v��p)΢��s=G��tI[��:�Cͭعw���_��t�e���A���.��$V�ی�_}����Sr����o߉\2�%K��S�<�c]�x��o���oSG��eaѲ�ط�]�*��3��NG[3�#a<x�Wq�u�@��'_ŢwW�b����{����[��]%�|���^{���b�xZ\O�8�ϟ���QUN�T`��_����8�ڊY�L�m7]�UUx�Ex�7�:�t���E���N����8r)�@���H�@9)��i������bKɼ?�>%"e��N�^�S�F�Bլ쓹���훱{�:t��C>5�`�!�>U���4x
��`R.�5�e8��S1e�8�݀ƆT���������=����O;Y"����
���HS�Ƃ�U9�ܨ(Ŀ#߀;�HbCQ#��+`)-����Z�+]���cF�Gq��C9m����
1-����(FG<��MX��n|��(�~�C�Ȼ�:�Z��! yT-]a>fr��@w[ۚ��h��A� FY8�X1$՛�vli?���������I�Ԥ籵W1��*��_�ўHg]<s/:OG{ڄK-ʚj7.�G�pe
&�@^���Ǭ��~,��$+h4j0f���z�2��a;���n��v�� Hf>��L����aax	w3�usL:!bĠ�c���{Mu��	�0�����/79ڂF�R=^�7&I��2�r��&��'X�sS�8d����d��x]J�S����<}=��'�<��@P�����N�H�9�@����{����@����:W%ml�� JD\��k��/]��Xdw������ �KBdW��g�^jY�-e\�T��:L<����"x���}�\�}}=rΎ'����K��".��b���A��-`�%�A�d4����f�ډ�̉ȗ��IE.!��=f����?����]�Ф,�;�EEY)�K+��Y�G#�,7k�#�U���o�[3X�hA��|Kd�e0��(XϚ�0�-ǻ�)�卻l�Tp��$ OiV�7S)TW��;)�R����4�y�,E'�I-��4���Ld�@渞y�#��D�;�-GuN!�D�$�� 9F�{�5�C�V� �I0RI¦!X X�h¸����5��sʐ�����Tk�����ˤ���͊N}v�0q�9��At{R�"g���%��"v��H�AI���`q򶊙��Z�m%
��D�-E
�Z{�zFH��7�o�8�[�b��5�w�}$���f�RRaɆ�H@3&i�/�C��t�t�����[1a|#�T* ����P�
��b��12������Վ�^��eyHX|)� ��F:�3��.�MW�CpG��iç���<��?Z'y���;�<m�*Oj�����g֬Y�={����r�(�|�rt��˩��#GԋP��K/�^�����y瞭�Axȋ/�(���Añ���L�$�zT�WB����0y�ɨ����!�\��C�Z��'��Haڬ���7�å�%��7���!,~w^��b�~���@�K����Yg�Euu����v Į����$�G���V��b��Ƈ]� ��r�L�ŵ�~
����o:��|f/�*���q���1C� U�~���W_+N�`�ݽ꾏7	���y�	%ܐkG�b����w��pE6o݅�7lBssJJ+�!q������"e�inH�^sk>�l��\)���^���8�EGK��U��(���>��$��c�ҕH�S�㦛�n�nK���'�}��S���{��������X���l��Ö�F�ABt����?M��ݸ��K$��ۧ^Ţ���z���_:�,�������~�%O����%��_t.�}��4^����CG���g^�K�9������ �1J:-~u��MA(\���>-�6�/8cG�1�G��Q���?7B(�t*M�h�Ɲ-�r!�����F���5OC��n}N�@uI�~ڏ�����z`Z�D��%>ds����;��RR��ÅT�����8ef̜��cF
���ȑ�x�OO`Ϯ]8s�̚1S]a���ZXoCT��6�jV61#;�	ĉŖm{�!A[    IDAT{Z�5��WZR,��P�����aƌ��2���˪1K�T(.F8�G��	�C��EP'7�t��>��6��ݝp�K.�E��3!��t�Aa�`�b}�hm:���f���J��.u-�����ˀ�T��+����I��/;���(�pz�!�WD0�sp�yg"�s���K*(�_�s`m�6���ؐ!;!�[���8Ye�	�9G#�i))�!љ�VV >�{�e���'4�H~ �$�	7ɪ�����A�9�xV�sUQ�����OHF���D��!��~���[���ꑁ �m\m6�A`+�	*�>; Q�&k)~�HيֳZ���!}qʼ*X6�;�2��B��)o>��Omz$�:�g���䢛o*����n Ckf_�m�f'a�;�4�	��ۉ�/�,�O���xj�G��@�z�}�&vS��E_�q����J |�L��N ���<>�0V��d��I�-��Ĕ�����y^�v��V~y��΃]���Y���[�d��1�F� �FB�C2�c�Ȁ�8l�]�s�Ԭ��D�������vA�,�
 ;!�xuR��@�hdg��&觉��r�Tq��d`���(,��PřfvL8�Y�l�<��`%N�$�M�p���T��ϕ�>K��YQ�X�"UV��^74��q�2-v"�K�I!q���08g��*5��Ò��Kd�!�����'�``��B	L@�"���(�|�Hjb"�;\R�R5�*V�x,^:���.;M#��s\��,)��duʲy�;\B"v�-%�AJ��U���t��çkW!��eL�lN���Q�P7ў�$�g�&�"�Gq$�[n�w�q3ƍm@��^z���W�F��DuU�x(t�f'�6�1�~*Rx���,r�Գ�QaJ}O)#�T����Pp^^V)��Ν����Oc��Z���!�1%%���f%����O�?����
8σ�9�G�\ ���;�D��w���3NW5���^I�2�c���B$R��$���ړ��5z��� �.`͆���bь!��R���p�Sp�_��g��L<��@���o��.�_���?
O�š���=]=rt�NEY	�}�-�Mȥ�"�WDH�eW?�L�0ЌHȬ�3�f�ʎ_���~�y����Sa��*���L���,���R)��s��k@H#�^_?�Z;����\r)�:�Zp���Sg����8���Sغu�<Q|�AL�6���fD���+?X�����W��c�y��6a��*WkOm،��Y��.\r�����KQUQ)�h�H��q��s0z�8���؏��}	���-�߈��u32���\��^U	���ނ��{��xi�*|��6nBgW�~��q:;�XU���U\}��ړ~��+x��[/�7��񃿯����.����V���s挺��k1atJ'H���-�����hiu5ʫø��+p�������p�[h�DI�Z���O?]x6F7V����O�1��n��^��>�]�ўV�ہM{ۑ����B"�EO7mʍ��8l,�E(,Bq���H�!/�(}m����؞�qx�f���+�=ۛy%��D�je�MP�ȁ�
?N�}2�9{G֠��(֮Z��.��ڬ30��^����,-7Z:���6K���ڜܘ�i�?AxV��8��P��ߧV:c9����ǅ��ᔓO���p��:%�!�R��Qm�\
�2�t9�z�a������(.����:	���h�	�A9!Y��k���]��~p�T>V��yn0��@�}��l=o�$�7尡VŖPu
l]��OY��7��;��[	A��<[|Y#�)�/{�7�&6����;��s��{#4�G�$�#[�捖�S�L-���Ҩ`Z�F	��7Ҽ�a���j%'�`	C�rI�A���lC<L���ʀD�T%��M%VU�\vmR �s1�t��Tj'a�SpCf�$7RS6mb�i�eAC�b��hV�p �z�|�ÄD���t���$�Oȃ�D���cd��� ����v��x��N��4|����'�v
�fu���xB��2��"dƳBj@&W1jR�8]Z��AH�]�
���g�#��H�r>����e�;=3�[�cs�q�W�=ޕ�B��dW%1�"���x�����؟�@���9p�q#e0#l��%��Z�ɔ�1�U��Jؐ8N�
'HSrZ��K��Y0^�}=^���-�#��T�i�F�����P�0�,uJ�]��3�����T����s���I���[҄�r�c`:v`�HȜ�( ��H�OPVQ���"���	��5��p6-����]�-�Ǚ���o��y�r%I�M'��s�ǍT#��R�a"7�繝��p���g�C�Qc�$x�e��@T�o�����<�d_�~�b�#�g��5��\�)�`|r(���Zōl�\�A�[����e@t*HY"�&���$̲��Ɠ ��V��*�����߂������sϾ�����E8v��n���#\Z&!����_�KF.K2���t��&�����ea�Ո����&NИdg�����]��k?�r:9[6���J���bu��{��!l`#욒+AO�tR�Bp��a�������'M���T��~�m���B9�$r<9W�l1,v�X�`�j�F8`�U���+���/v����XVh�ljH*V��N�׾~�y��(�%���ko��g^\�#�]p����66�=eŜd�]۷����"�������lZ��@q@�%)���d���p������tT� �$�'����Q��~�r��y�ǃ��rA���%��X��'̞1K�)&Rq�m��O��Mx���úui����٧�?�1F����Wb�ʵ�b���~̙s:�>k���z�PWF^U����I�Y����/��矍�.�X�����0��{������Nbْ�r�w���|���X��*,Z�G;:p�M7�[wކ��$^\�Vmځ�:�14�?%�	uv���>@��� �7O������%2�-�7�����ǟX����Rq�P(�ޯ^�b�ǿ��ƫn��"��ك [����U�b���Q;j܁ ����r��t.{���e���/!��ǌi�p�50���dT���^�n�R��:�:X�ҵ_�-p��7\�h4-<&'�H-�b�� ��TJ!&���~����(��c��vx;z[�r1A�E�G�ȶ�P�p���Kr��'�k�ĕ.���碐O`Ųw�y�:D���6e
�*��g���bi�rq�2��;w�@wgH�>��99rj�qwL$Y�ۃ���c�޽���!�֍��/��s�'i,�@<E�Ј��$a��l���4�9/\�J|���.ބ%+��f��;��#��"�l�$,� ���Zސ_�:�VPj�����:t��6�p��ѵ��v�_�!L權����ϤK/K!��`N�\�#a�v�\�}Ʌp�=h�iG"K��S8S��+�I�"����p�تX�At���0XWࡊ#����ɖ|�00b���B\��KN���xצ�=@�UwvZ�A�� �L�o$F-�H�v�Df,V`W%k���3a�p�i�&�� 2'��5��Ov�e�	�)&#3&���G�d����|�����	T�.�@�ץ붓A��K
�����'�-�$)��2βǃw4�z��9���l�G�Й`�[�[����a3�B���_'�v���A=;�L�>��Y1�a>JY=�|�ENg�?0�#����]���Y�!���4�W�`��Zɑu}
���"m>��Ngg��W��� J��^�
�P5����,*�e�f��N�:M�s4!�!��ɨ���l���*I���[�)����/U�������YU�5&�ڙ�yRb9���rӵ0P-�e�G���5����dë ���Q�,_D�ܴ`t������j��d���\�)8�P��&,�;�����	�gJ�	IV�",&����mu0�{?m�Td�>����:s�)";Z��G�LA������ʿ(Z�w�8�'�l���<+Q0]�deX���g�<��*!�)���(�._���Di��e��R�!)s������_,H2���K����+p��b��FdS�3��/�g?�w��F�BUu=Ǝ��ѣ?ٶu��e�>s�R��.�$��~P=���Ғƍ�SO��g����:��ءommǚ�?��M[��b�+3w4�ƳsVP܁/&���u��@ǿ��UJ'1y���G1k�LU���I6&�xێ/M���ֹ��(u��}ɝSJӖ�KW��/�Ͼ؆�(�C)%9	��0��)x�{p�ٳ������;�W��g_zM�:��^� q�k@e�8�������!�!G!�X���|r��2�$���Z��1ޤ��_b���	c�y�,p
fSU����!x��.���{�����Ҷ�V��Ӧ��t��g�_~�̘rRTet� I��.����;����	,}�}A�2�N9}6~����x}�2��b���`�|�#Rt#��O��\��S&a0��ҕ���3ω�v��W���/FYe6o;��_x�>X���|���ŗ�G�@G[+�9(�����!z�{+�x�2t���[oƽ7݈x"������ԓ@�`B|�x�R9�{{0��_�������e�^����Gc��/ϝ{��W���(!x�Ppny�/׾�h飳��������z�;�n�Z�߰{��g ����*u���.Ăy������K���O�3�V6hp��z҄�j͜<i�HKNBC2l�S�# �R����?ޏ�[!㮄�_%�5jlJn���.��'A�6�#���绰m�G9�(�d��v���Ļ����Q��U��>~��3�1�ÙÅ���7,�)3&���0�ڇM?�`o/&������͛������knV@2}�L\��*444�[�@�
l8r��i�D_�]{vKW��s���-<:��nC��{Œv#n]q։��I��|�.<��CtF#�j��t�ÏAU�(���8�)$A�o�Q�a���ٽ�--@gK�"���߀��l�+\���J�2���L%;oȡ�� w#�ץБN� θ�<̻�8�>4��1M�m��0�ª̶���Ą�N�3�)���V:�ɉZ	A&o��(Y�4�G�9�b#�'�B�	 $	?�ު����H&d��`ᘭ���Y�[�^�&)0R}�9��|1����K%��*����{�x��_�'�����f'!�
N�d{��U��`�-�ϗ@V�U>�"I�$T��>�w� ��^���e�,�K���X�u
�qq�c�$�<X���0ؐ!�,lWD�.	�!湛���!W�	���I��2�e���wB��� SI�U9f�Ī�%�E�Έ��id������'�3�P0�	�`�aTvg�Eb-�Z�T֭`�F9�V�q&6���0+��us����*7j��K"Ad�q)K��������@���)(�:lLtoe^��7<o�����uK��m%h�9X�9!�g��Ύ�p�k��1�{�J/ԏ�h�ˀ��<3�������7HS�ά��9iا�a�3�%�e�=�8��x�����M�p�x��!�؈I�ԍcBo�qΐ;�s�����N\��n'9&94	q�Q6�D<,��4WTR��3���|��q^�M2`慕�Y�>?��X&c;L##i9�G,C�&��4FV�!�Պ���E��K�>;�<&��>��L�,��[@9R�D
i�{��W���܊��G)qa�C��|C�	DJ+��8��v:�L��CG��sۗJx/�eOg��Z).��NsT��¸1�0u��;�LL?�ͭ2Iܼu֬Y����LJp+���s����}U��4�x�}�I+�n=7�"a��:���������^z)J譄�DU�}@�ev�8cq�&�k�s|ѫ��gJ���0r2Y��؇�"��D4�4y&�Q��Y�o?���?S�b�O��o��^X��d{IӠ��l
�rea��{vlCs�a�3�&�Q_[����2v�1Y}c=�����pW���/<w;9�c�ߟ(�¢D]�%�;L�\י����AΧ[�!��}{����&�|���� c��A��z�T�,-�����g�[�Qq��g�z~�دQYW�W��7�Z��M=��R����>w�X/�M����
.��D�9����x�O(����;q��#
b�������JF?�Yg�����Ξ���QP��4T���^,^��Z�݃Q�u���-׉���K����q�s�l��T����&���?p7�/8C�4�%,{M�����y�����_���C��Pp-}��^}k�ϋ�K���R��C���V��>|����Z����#R�5W����3s��O~o��&J�G������?g�~
ʋ�H�p�p��y�(r��I� ��i3>�l?z�~�]%2����b�3��Y�u�ȼ(��XЇ�{�z� �C=h(���@���hۿ�v��#��IS-<� ʫ�QY]��d�=-�2u���J\0o��BȤ�ر}+�|�R��$��7F$,�����ۋ�h=��b�_|�8��yzB"�y�>_<g¤����@�5�}ͭ-8��&���)S$�G�K.dL|X����G��xb97�I��WW`���(G�b�D����.=h~���~�A7�˃�o�����AwS����[�D4\�ʍ\��M�s|g5����j�+
4��ˮ �;i�S8\�9��s/�G�G;[�!0Ҕ�?3%���w-c'�2l�;VdH7��Y�$Z����GU��@�	O.�\:i*w��h
�m�3�٪V�ؘ���
���b �[�S\V����O�Y�'��$;'�O �m����W^��dd8� �$�m%kZ���@Ql��`��Z��P�Z��dL�ѷ�"�ֿ�	3��snv�۪�RԒI5����u�J�,��O#=UǏs(�����@�Qѝ�=X��%3ʾ��x�FɈ�s\1ˆ)�����Cb`��rL2P��dp��ň	`JQ��~��$ikY�2;A�q���j�)W�b��*�q/[����o�Dy�:K㜉`4�/x��	0�ټ:_|�fC���V����չ��@�(�ء�� ������r��b��z�jl��L��/��(Q�������q��kw�l�Lb,�LV�� \�Ҫ����{�Z����tP&wv7�x�݆&�5��cun�����9q��SR�cဢ�s�����Es.�5�/���c����@�$�C�a��'�l�	�����4H�L+��)��Sǜc�w�}]p�R][�TV����v%7E��j7�z��� >k�Ӆ|&��H0	:8�rÕ����1��V���y����2.,-�Ĕ)�p��9��I���,RkL2���R��0��$���K��(��`d}��rN=e&�i��ի�*L/?SP;¸D�6�JRF o}�C��oH��+�궁���Ĺ�N&�����Ž�~ӦMG6S��e���W_ő�G)��=�b�y���!��K#U�ǌ�Ƒ��>ڰyg�M�n�t'�C���igL�7�s�%�U��>�sU�4�3ӣI�	�"
HH"��%�1������8���Y���`���L0IB	( ��2J�0�<��9V����{W���|��^KK�QwW���o��}��������VVQ��9ɭ��>����15��*e��c�voO?�=�\Q����2%���ߛ�ԜڷÇ_A�V�����d(��Ţڙ��ׇ�C&�/��^{����&V���N@L
�A!��x��{�Y!���7nx�u��2v��r �/U�}���Ï>	���i���\���������wމo�r;���~�y(/��Z���2�O����+����܎��/���!x���!��O{߸�6���`meU���+/�{���w���DK˫������;�م4>�[�'>t#j��v���݇�s�u�U�`��f���w��g>�	\z�k�R��k߾w�}o�P�?���.����Ͽ|�T0    IDAT����O�!���;���G������V�?��ɮK33Z�,�C�8�tu�B~d�|��p��<����ރ��4�	�Shwlx o��2\q�E�E�d�L��n�g��t���E���A,��hz�h��5%�-*N%l_h��g��a-��r1+���R����1w�9 ���c#�=��!��C�� B�(�V0>1�7\�:\~��8crL6��f�=�N�:�ՕeE���Jf�L���Ռx�t,x�ފ����aju��i�ڔ�i-鞴�1A #�}��C���$�#_�}��P������t�>|w����-���#>8.G��h���|�AU!/�� �1
����
t|(-dqꥃh.NM����t�ڵXkSD��i
E3T1�2�:�t��&`'��'e�t*��/�DNC���֖Q���L���I�� 0@Ͽ���H��`q�s�o6<��ak��1��[$7��>�kjUG�N�(�&:bt��:mjrT1���R�F`CA Q�-|�,X�4�FB� ���>ǭ��6<�!p߳�sꀷ6��~�kd����v���4DX��(���<��1��l(�~��g��Љ��c�bBZ��n
j(0暻߳^��z�7 �!�"݆�f8��Vd�bvTV���R%��*`�Es膺�,6A���h;�ZSn#���3�Ü�0fQ(HL� c*���N<Lrm�L.L�{h�LJ��1)E�B��V@��4��*����l�s|fy�ҝ��6-��m3���b�JA��{����+�MC��u���e'����d%t�p'U�il]�_��m,��	��!pC�u��Wwo |�B���W���Y�,����V��E��,�Pǲ��HJ����a�0q��Y0ʹ�.��E��CpM�i|��6D}���2����oK��dsP,�LD�.�m]�e^�k��n�FX��n�=ϫ㲍���u����3j�Jbx��(�u\��Jp]q V/�طu�O�/����UD�0Բ׏�ỲǤ9s�ƽ����J�$�!|���>p��*ܬ���_��5|��_�����I��{6�Ln��6���S����T�a1�p(%53W�z&�=�z_�X�\q9vLnE�g��EfI3�*�g�����K�J�z
��X;wO���s�R�١��+��m�u�^�w��@'���O��_F�TB<�Y����L�ߋ���Ӏ��g``���<p���?y�z�;�2�<.��|��g睵"Z��&����N�z�qrfI.C�P�ZK�������s�٧��8�p�k��pЋ��Q� �]�2�0I�&g�����k�K�.Rij����w�ܭ���?u�l�H*��$�߿?��~��������k�p�t,��&
�y��x�l���?������D�������x��s���������gC��ՀV�ٳ����p�����[�����5�|���uo��H?�����w�P��&�����nx�����n���~'ݶX�1��ޟ�����}��'>�i\�v���w��K'f�"2�k�c�Xۋb:��/�����q��c!Sė�z+�}���Jz���.��O��������=|8��y�?����	F{����`��F�OnF_��ǁ� �cd�_p�>/y�a���K�����	�����׽o{�5��A�L8�)V��8|� �M��'����c�BY9�O$��%5�.a�Sze�H�5W�!�c|d��*fOB�S����©�(M�S�jZe$B���6�#��"�ka۶1\x�Y8�Ha��14U�i�>r���߇�Qd2e�޻�x�;p��stඨ��Q�|׀?�J�����Y<@|Y���jF��;&e�ǃ%�c�^m�ӎ�\�u�cx��X��P�&��7�D��<).��%�ۢ�O h��@�EB��A�������C�Ν��Y�ذ���Nn��6N�ޚI/��=�m1a��)*�tJ�{S��Ej"I,dVQiVe��Ô>�r[��4+ޥ�k��a^�?*�jdh?֎���e����)�J�}-V䤲��/�`�@r�m�����q��gu� {s��}�������4*�'��l�u�'�'��N��Y��7_0� ;u����D������Ы?YN��������\�|^��\��u!j�sŻ@w�XZ������66@�]7D�Xskp�8�x�6@�D�g���4�/����o�#o�R00>�%�m�ᶺ��\&���*�
BkE��_z�9I�����L�bd ���d)c!���z�����4gY5��	y�����g�i��yQ
I�cG*Č	����l]#��2��HK�ͭצ�6e����'�lB���k@��p����	0�8�v�x�b6![zl2��Y�\�ހY��EO>\�Ca1�3��u+n]u��͈\��z�u���1i���*чl�s>�P���Hw4T<�����uǤ�M��}����|+σ�˼��84�.�a���8��Mۆ�5�Q�2k��|��z�b��~FRQ�f%*�峈���a��Fq��C�6�t`#��QA>��T2��|����{�0�
m����O
/���ر�L�ر���� �����e:�6_����B
G
)����,�RD�#�i6�\Kl���ׇ������3��Y�j�����hMm���
YKBKhM�{35u�|F�T:%Q�� �h�����
�T_J����aQ�(��T}ppmo�]�܃�Ba-�()
��,.yݹ��?�,�ٳ�=��6����㶻���rQ���T�bzz�H\.C�x�<��Ve���q��UGuX��}��pl=���0~�k��}�R@�*iXb���Ie��Ф�"
�٤-��
!��y˖͸��{t�>���㒋.D<F�\F"�� [�5e�/���ȳW�W�ޑu�_�����^�B1�'�z
�P{��Ț��Lz��&�\y�e�u�>��fq�w�{�}_�C������>�쉗����˘_��^v�m�r�99����o��F���hc5�QB�?{S���w������������㕩9�8 ��]�����Û��fl�9��l_��]��?/�.����7��O����=�ݣ���?!x��ӽ��;�����?����b�~��m�ţx݅���wD��#/��󷨖JZy�X�����AŒ�6�)N�/:w?�|�58c�fM"��&��B0�?�Z	���)<v`��(���fn�&n�p�t�yR
|��N�f�f�C��:>*q��F���h����i��!�e�B�Wm�(���(z�\ULn��=�14؃�?G�Z�@J\�c��ŗ�ñ�1=u
�l������9$5᳼W�P�P��P���,pR�M��h�P����S8����%��{���o��ڹs��%���g���|;��􏟅B;�N0�6'9�6�3�i'�|���|55D�C,�*��W�p�$�s'�&7}��FRv�]����i
���m��{e=�¢L�k4zU������W��^s%=q#*��z�>z������ɈS��\�g�5�:N��с�\��qf�EA�?:�4n��b&���ą���U���,[�����(w�?Q���y�2��\��ޛ���u�Y�
d��\s�bd�ּ����n�\w��U�,bAC4r�m!�ɰ���"�z�������[��|v���FUb���Z��~��Y�[q��C�����Q>֛�.EҺ���v�Š���Ϫ.�����Sa7-������J"�3��;�!E�|}+,4�cu]�J6���kݮ&;�2�
�6��r��&C4�p���R^��!xS,�"��=�O.JJ��@�h�Yz��J��O:
�B��SnuΪ�W"�S�;�AW=�ƈ����s+�y�[TvcA뮗�k�:r��M�M!l�u\ӹ�9�^맭�a��7���w�4�*ǵ�A�)�r�jNC��k�=�K�8�#S�.4%� �'6�����knE�v�r���lZ��5>f/s���{0����p��ה�/��FP��QZ����4	���}X>}\A��E��E�T���X�2��W,���Т�r� �F)����>���}7]�͛D��s���}_�ڷ�$(��������&�.8�8zz{O�Pm6�+��{ﴥ��O�y�vP�eՐqP�g4�wt��{�037���R�	�iiF�eSvύEe���s"CM��J/QgA�|��$���:�{�z��4�H���	��)�Tg������z�ʱSx��d}�YZB�ZVH\�^�ŗ��?���b���4�BX]]�wo�7�q'�Wr�S�@�Z���S�9�h���{�����"2�j�:ф"�V��B��:������	ˍ���*-N�}�?9�O"���*�=A��j��� <�<��8�7��شiX��U��}.���wʹ1�/c%��/~��
_kyȕX����މ����`d4���U�/.��&���HH_2���Ѣ�e�́���?���y^L��|�{p�uoC4�Ľ�>���_��|^Oo�lQo�\q��g;&{Mh�j?�1�w�8q|
�{�M��܄�x��Cx��#X�N)�m��Zj�.���vn�a���Ï�~<�Hin��׿��?�������>����!��������O�y��O�l��5g��AO4��y5��bz���o_@v����^�� ,�+�2r������d�K<C_�gl�*��Bk�|C�PA��	̧�x��x��
r��/ʥ�
3:�p � )D��چ�UJ�ZC��I��Ϥ1}���E�=U�y���P�-��2��*�0xz}O0�R�V,�P����>��]{�U��ګ16Sg���n#�_��O?��o����7�x��GWo�)�kMDC~��P�mX�ZXn�bK0�sϿ����Q-�Ъ6������4W��w���K.��{Q* _��;���%�Fv"20�J'�"���<"�|PPʩZ�����H* O��B�Sm�!��d�|�˳�4�d���3�Ąd��ɔ��1N?`��W�a��<�EoaA����Z���I����������9�u���M¸<��8����eU�`"�6��In�W)�s�U&vC}L�RZ����2��F���F��nD�Jb%�m��F���,2���[<��y�4�4y�<�c�:=I��|�F�h���ˋi2�tԐ�L��r�v�f���9�FBԏn7��m��"�rI]����&�N��S���&���fZr�qT�Td�P�~gժ�M���e�?�~�Ud�!0�װ8פ�;�!;E�M�l.-w���Y�v�o��˙�7��+>X�7uDER�I�愐u�z���]�5�H�6�7�q�p�K�u\�H�]�Hb��i|�ke]�4��-![������� F��DZ�P8�
y6��p��s2����� 6 ̬q�
p0` kg���E%��rt^��w��n�`�{�Ap?ǽNZ5u����_����-2���g�k�G-���P"��t�(��̾blo�3V��Y��o� [�06�������6\hX�`wH���zm�����;:�k���t{����5 �Y��)}���ϳ!0�;�m5>a�C^��N��Cem>".,��,�7�C�(�KjՂ�A{��O�&n�����/��?�_���ar�C(W]��⠾��e!����'��NQ3ғx��*:�:"L������F
F�����.8_�Z<������XI�ɉ�띃&5��y}H����3j;f����D�kA�|.�s@�Ki�����׊߇D*��Q���ӊc�@Q��e�波fQ���(e��4p�E���ػ�}ޘ?���,n��v|�������꬚�Yz�062�}�iL�:�F�"�����X�J�J�����^GKS�7:@qߡ�
Q6o�y��b�� Ɗ��1���k����1U����G=��Z�4O�w��{oz���<���<}�y<��a�I������Op͵�G_?�.���F����{<�6*�2>��� |�1!}�)���?��{+���a|�[��J��f'��7��bc�Q���w�C��$�����?���{/�+�x����>�A�1ڧ�U�mH�]k���ͬbhp���>���s��S���������ţO��]�������^��i�{����}�{y�S/~�g�d4�A����ҋv�w\�M����)|��^9p��z��Mo��PB�:�+�U��a�%(�8}|�J�^����0*0��Xb=X̚��c��7z�����x�I��hW�Y��p��h2E���J>�|@����shU��k�-����Eu�@�N�y;(��G��O�>���Ɠ�Gp��a�]���t �<<:�P�w�Źe	��d�O�]��j�H ��<��P%�ڤ0%-T`ye�A!����<� �W������EL�TB�E�����mx��Ch��݁���&���r7ufX6���[B:!
��#��js��z�4:�Ex�LϬ�!`:��h����yaaUC"�lt.�I�^;R�R��h����o�������:89Z����:z��\y����Mw��+
�c��V���Yί��7p�:��h ��'=��~��G�)	r�qV���Q
h�j~v�����'g�aj*�.��)�{�uY/T�f�����rAFn�t*��l mC���U�ʐ�T#��\��/�_���ES���5@,�MQ΂�_]��� ����J�r�����t���A,������4��H��j��q��˭O�I] ���LS;`P!��� �i�,I[Ʒ��!򾽖�a0z��BD:���0��t`�fZk�,�DTp0��כ��Y�r,�b"(�(�b�M���\?\��$�5i8::���>5A�N�&$>t�i��TQLlhtj�"äYg���=C��Zfm<����W����)}������j�,��BN�:U���V�4D�
�m����C��d�
;�߈���f�͎C�������#u�\zVt�4`�=�f�Ar�(���}[�k�u���Ʈ_!�a5��n&�K���/ol��>�(]�yx����j���L��`_�|>�lQ�`�5$��А��h	�F��*�<��(�R����̰@�F��F�TQ�ٮ��F=��ާ~7���1>ү�f�ߐ�Pn1m�؁�Va�c�`7͐��zx�O��#X���&*x�҉�\&ԩdZ5���1�B����|v��-[ә�y�ZD�:�H �T١�耆�G���+v���b�I�WS��}�ӑ8�5�&��2�@?�F=@,��k uA�3asʡA��G0чP���W����i�5�9朻�����ۃ@��<X^���������:>��DRMN.�E$�UW��#�x��p��!�+Q`d�_|Z��у��#���g�J�6��!�A�K�]Q�;^c�+�I�JH#S3ժ��J����	�&�s��n!�5_9_G4�<���Iϕ��G�h! ��B� T*��ګ���W��R���� �k�af,��ԓ<�����Ï����h+H೟��}�;���⎟<�\�O0�H�G{&��jagl���S��׀/��o�+~���Q)0:2��~�ݸ�u�a�?
�,�"�����ͤ�����K���'�E6����Jem����᭿�����_����_�2�����������Ƃ��N�#�2F��\p�&��Cx���{Ŏ������#�>��BsP#=F&����O�	i �7�3$�o��|L7m�#?o(�\͇�:�G_��Z9�b+�[-�������5�&��_4[�����1K�9�����9dW�P�̢�_C=����QTWf�JѴr�@1I��?(nn,҂br%_��;�k���#� �'Fq�Gk�    IDATÂ�<�����DLLL`߾=*���qॗ1���b��VֲBX��
er=x�A����lx��ʞ������m�Ė�{���P����A���	S��A���LQ
�{��Jn�@�'�0���%�8r3�@n	�F�4^n���s�fSpol�ͣk�ĂN���:m��<@jhH��W]�FЃ�K���+U��vиKFeC�����Fʅ��-�_(�)�D�V���t�&��"���p$(��]nR�
�@���*'`L'eA�l�\���Dt�Ri�V(��B���x@�~dy]j�}��d�фL�b��~����n�)��7S��k�m�Ҧ�Y�c�kp6Ѵ�c�J1�q���QR�,��D�B<��i	���6�݅.M�6ۖɼ+^��JW�V��i�/���`4�;Hf=p�٩�j����;�E�i�u��˦���fUM��N�b((|�*����;[G�(+��EE���k�_<����L"�4jR�x+|�7�k��g��ŨiN�]Z������]a��]����r!�V+ISD=Lќ,E~87]6>|�������+�?�~شf52v����bUG�q���u�Nos��]Q�͵pz~f�����b�6J��H�[�눁��p(�-�F�5,��ߎ���T�
)sRss=J`֊A��IC���y�v/�M���X���3��b�hKa�b�*�?���?�>�iZ�G��V����>g�L�Gm`& Q�]
x��F�^��E��t���j��;��VUUY?�!����U!��w����R_Լ�zHѲ�Z�&m�gUЪ��{��O~7���<1"�r��G~_��o���i�t��)�@h"�J��(?dԬ%��%D�45��&�|_��) e�z�����g��3/��
3|��'�	<���`1	F�3�����ب�z3ף�`<j��:BX6���.V�Ѿ���5K��̸�� � ��U��B	�R���� �YFqaθ����}x�U����w��D�^������wo�M.CWy�k��C�\E�'�+_9FF���O��WЬUT�0�Iz�:���+Y��Z��i��7o�~�5��o]�I46a���ڭ[��Z��JSZ��^3+E�B����~x��jU�NKUm]�r�Z#������
�
P��	��K/�5W�۷�B4��z,~E#!�,,��_�/�=��Ss�z��@8����o��R!?y�!<9�v�� �MT�����r�fW^y�y�[��������/E��&���x-�;g?Fb)�ǒ��IY�4td_#�ZË��Y<��A<~�=�4z��Xo��z��~�g���O?���<��������_��^_�w!O�H}�6�l��uo9��;�\�>�<|�0�9�N�P�@! �VK�ey ����5L����g����;��d*b��C���`�?��7���r?}�(�4�	0b�|��oZ��ׄO���@�?��(���]Ά�ը��,��^TXY#����q�LCym(f�d����ޝ0��N����I)�2ݱ$�Ѷ��ؼIH��v�Ã�D"!M	�F�q��N��b5�CG��1^"A��
Ut�1E��b~yU���Ilڼ��aK-�[~�R#(�(4=���Hģ��˨R#a�kv�lhB� r�,��*�����bX�^�̋S(-.��2+�����j�7�&�<@����\%�4n�F�&��P7��.8:�}��2t��/E'�����ͺ4F��.T4���kr��Í7M��&/mӋ�2�"���9���7�욒�Ñ�x�##C��P(���Q,5.M<p����A4���˴,5
�7C2��e�ҘA��V����'�vl�ύ�5�~�#��<reo��d�g&��E���w�w�SǫI3�k��1i�(Y��)�T�u�a����uC�( �OU�f�ɯ�m����6㦙�s1��,��l
.g�h���b1�(=J�����r���J�N����=6��6�>sC�FS��QCc���.�Ѫ�H�k��%S7E�-bI :�b��_��v��m��'����h*�(����X䄔�~�x��3���b�;�~�c}�Ɂ&rf�s_�Lνe��
A����h	g!%��&��An��Զx�)p��_�ø�lG92������FKϫkY�Y�4l�r\q��w2�5
n��m�]�WNVG�YoƝ�)_��V��ܾ��m��XMg��(Xm�gQ����Ѯ�>��Ym�}�.@bm!}�n�k�&��#5�r�2{�9f�����V�>'���1H�	'4��z��&�r����m�GBr�/��Op�4b���Qwd+��\i�&I�{ =��B���w��vLNn�n�hi��?�$��Ew"i�f.��v�|߲��L�_�#d�L�-/�
O![�_�h�L�LZH;�k��+۳y��M��@�Z�����������{ H��x���y�tl���Ů]�q��-z�ڝ�
h�8�dB���鼳ϥ�p�"WP��~�HI�KyRg8H
�� ��aM�i�m4�9$ca���}��{IIެ�:�a-��-�߁o|���_&��Ui�1��K044�G{�|Y�T"�@o��n�r�r�[����H����4{������;��Ќ�0G�Yr{��HR����=��9(*��H�$�z�}�BZoD$�ggt}z�G������sExAt*E��>Lnٌ��!C'�h&�:� ��2f��Ih�(��A��$vm۬=ujv9%��h�8@�ˢ7ʡN��z�l�=g�C$�ZzǏ��Jf�v��}�FԹ��2b� �z�������H*u/��<w���VPny���ͷ��'���W�[���3�6�]�4�7߸��x�����1�/���B2B*�ǖ�8��p7>|��HR~���]�+���i�ԩS��3Ocnn���G<փs�:W\z%zS��8�6n����a�<���q���P� �ބ�$�(`ż�B6�"g�*Dڈ�M1�E�ŦC�UC��A*B~m	�Diu�R�)t�V�vh����4��GSa!
mȵ� KS9�lKh�4&bR@ٓ�G*��M5��d4T
��� ��1���B���o���!���i�Q.���oɞA��[|a��w6F�7+�P����P_ z�2-7gB�L��I�!�D��� ]�(��!����CS(�̡����QF�C����i:���<�;���ʟ3jG���+ca�/�9�I*�Ӄ�/��}���r*ԫ����Ħu��֮QG���"�c1%`j����fo���'���/�A8A1�E�UE<D<���q��1	����9,�dp���V�G���?)�G��Zc�C�<@$���� ���.t�k~z~�B�z�kjltYǺ릹�O�m��f��9�S�r�iSYCS6�~U�4\e>|om�r!N�B�E�4CI�����p�r��|&tG���D�\4u�ڲ�[�eP�4���x�� q!Z�ڤ��S'ֺ�����4=�bh�}J%%�O���$J:����h8��I��
+R|A�y��x �}Gc��C�M4Tp`܃����k��i�7>U�=�\�c�H+"�����F@Ȁְ���3'������H�,�t�l�)5Jzn��I����Z�뿮@'RX�G#1�r�����Mp�hB�0���}�FC�[R��Y/r��x�l6&�¶�ʽ_�4�����UMQEPf��S�e�b�V�� n|M6�>Ni-�,2;�VB����{�"�a%���<���0��`������1M���-��1��#W:e:tfP��Akok'�ZK|ߴ+���4�ؖ���&I�\k�
����!�aG&�ۆ�Y�aC�j��1ٕ4�Z>k\���i�b���� O���3�qꐠB��8�٠�4���ƦgB:"L�Nv���ВZ�&�.PMȔ��5�xZ�Ƶ޳���䱩7��X8~��u�����O6�ȏ̢4\'�#��m�������KNC���*�q�U�"(���CT�����T��E�Ը4%&כ!�b
X�z_o�z	~��V��+�3c _@._�iG�	�,,�?�=�4D&����>I�K��'�)�J��qx2Ʈ[p�%����ئ��q݉VR���˦�Ke��ƺ��X,+l��%]�:�ᠦ�J��Z�?CDC�sh�a�Ո[r����l� iE/���W���-��ͷ}���t�~i��
E�k�p�����g8q�X�Ac�a"�}�:�l!#�h���4E���xM\�+C�!���y(V�{ɺV��.p]+(РTל�GtMLsGףx(,-���f�P���76�P4�ӳ+(�k@�Lv�<��j��U,{�S�ϡ?�j�)�y"\�q��=��6��2����Ec�V�?֣�s�H����^Z�?��Ƞ��XO��%�baL�8�p K��j�X�p0�(3@3���A��F�Vњ���4�i�ҳϾ�͗~����{���i�x�-��������ٷ��6#��:���|������ކ�&R��pr����"ۨ*2�B٥Ez��P�U��oۊ;v!��1���@�@�Q��!8���e:�{S�xC�	�`����]�)�'�z�^�!Q��&`g�1�͡����8y���C�UC��D-����,*S�w8�(i�c1χ3���4՛�S 7RN�+�`.S�;����0`�A8Ef�C��� Z��9R(:^��!N���^�#K"K"I �7�J�p��D�@�RC�����i�| X���ll>���Q��r3y�m��(�!,X^�"}rk'N��[��Y�h�4��5+N]��s<I���2BbM�Xh8<�d�$ܹ)u|�z�p��W�+.C�,e�Pcp��� �4_�Ym5"<$�*���CJ&b�u��d�OF�xQ���Y�ͽZ� I �c`K�*ӟ�8c�VLn�@__BM��J��W�M���Yx=!m��|^vzlz#�$�
L���b�X/&'6iBQ*�������
�VP�(:����v�-��G���f�ˆ!Dn?Q�F�H=�q�%�m��<>3�$xPV�p�fخ#�c&�>�N�z���jG�lG�*m�k����_�X��(r����=ɔ^[HM�%+@o��g�"���Ȝ%���c��܇���:�O��y�T���+(3s��D �3Y�5�(���e&�L�#��m�h ��9Y�sa�>LC@{A��H�
��d����X7�VIlg\�7wM��M��Ն
�F�]�C�|���L�b�A����J�c�Di��'q,�L������'���n<��3Ң�	�)μ>�}�׌�k �T�FS	��D�Zcjz�[d���r�C��?f6'"fѪi��K��)�XT��&zl�����z������7�M��ll�F��>6nS7&lBh
R'�7���2�v����ma��jz�:��c�,� ��,�Ig5�~;�����%r,=�-�y(e# t0H�Ѡք� q��	�I6����R;��iK-P�j(c,��ZV����]H��	>�A���UGd(q.qYT'��@�O�c���2�F�ql��҉#���[Q�d
�9�P=�Wr}�R����ڪ��ˈ%B��} z�H�Q)���R�:G85�vݘ�qHc㧉�"�Ex�Z� ���Q��G�-f@,d�/f�z���CS�k��n��.|���ıc���\ ��#at��>�u��������s��#y�=�Ll���w6�B�8��}�TzN�Zs�В۳�c����a��`E���d�0���E��Brpb>���P8��ͷ܆�o�3+i!�jv�MsY����k�<�aiyA�/���e������b���_,]��Br�q���4ו�㬀��a�!�a�=��jp�:e��������rKՊ����2!r+����}��,���6�Z4;��M�9Ҿ��{>v�Bi��U�b#�5E�3d~F6М!G#��$�&�����T�e�i��~��%@S�j>'[^�*���ZR,3ǡ����5.\���E� ��?;����̳7������_�����yb�n��?8�����&��	�y�u�ba�=L����o�o��L4*U������I�w5�"�λ��F׬u��0wzAm2�2�PQ!�s�^�a���4�|�y�[�h�R��#Z��L�-/+A�#@.��8�}Hp������?���d�h�Oaen�R�zY�Q�����9�fŸt�8�Q�?�ǆ�xȍ�֡�<�PK+k�4qz��Zr��������<�4ĎP�b��w�D�|u+���n�.5���g�w`�Hm��6Iu`�ghQ\�b�+ѹ��}1�͈y����Ʀ�`"�`4�⤚�#7��գG�ɯ��!�$S��[�.��[�lEmC�Z�$���Ɔ@�<��3�	o|��p��"[+cvyQ�,,i=ǃ��&�u�0�F����gsAc�NKLoJ鐡09�5}�l��cG��ϔ��TL������ܳ�(�u��|����Vs�7$a����5�]7��q��E�"^l��p��kjW:^L�/�0������qj"q���d�:9�!�����H�\RZ4��w��?'�,@�h���>t�z��a̯�9���]�A��>)�5NЇF�t=���i
����
N����J�JYt�h �T0�h0�����y#<�:�4k81uJ��,XY��s$z{4����
żx�>o�@�7����|aY�-�7��@h�^1s8�e1�� t�Á�h8<���5M'}�N���E��!��:ņ$��\N��ZUN~)(���o8$������В��͖��{<�yX���B@[�H�ڄ�y�t�!
D�	Q9}[˘f����Q�L��$K�mMC�R�WǤ�j�Ɖt��\.����;=n�C[��X���b��߇MSmi7�����d��VC�t��;�&u�%H�z ��B	�r�j�hk�""�����4+�5T0�.X���)$ח?`t#
x�?MҀCG|�s
L�E�;����+D�;i5j��~y<oD� ݔ��F'To�T �3�io��3k��	��zY[+:7E!V�����P �}�q�ZU�jpy�щ���-�2t�g����.���m .k�8������4�1�r�ʹI�9'Mf��v�<���DB�2�Bz�����*¡�������z���!�a~qN��-[�c!��ߍ���{�uS�ɕ�L��\z���&-�����ֈY��L�\�i_���9�0��"f���+�Tqx͚�F����}ߓ���'<���#3/��C�I�u!�#�w�i>��\�f���wm׽Q�T��Cg��$�7͜���GF�n�$���쮷�h����ǃA��8=I�C��w��V�-Df��G��+��[ο~���ͷa%[4�:!�@.����^�tû�ӓĽ?�����-�%cIY��xMi�\/�9]K�h��f���Z��3�5��!�R@-5Q�M��RsmB�|�"D�y���L݁ix�B����pO�땐?����p-SD���^t��K�꜄l�f��}rc��N[j�a�Ў11�$�fW��I�d�X>"�(Z
�5�<�U��ҾI$�YC��C=�������	M��H.�e�-����L���!x\]����7]�'o��>��C��}O~�?���'�ڤ�b�&}j�:��U���ُ��l����?<���-�[�w�YHF(�1Zӥ�
��ů����T+�z�w?��� �{l���,r������=��ٚ�I%�Z��p`��*Ӎm��D*5��< R�8��<���X�?-�z�d�NbꥧPJ/�Y���q�#2� ��W�d�8���%R��:���-X^]��'4�
�a�Ý �K��4�����<,y�E��;�X�K��Y� ><�g�C$ދZ˃t���xZL�s��b1�		�D�'O�Rz7ڶ�'j�c!5�09o���'i�	�    IDATO�%�8���k�ƴ�8�3�"��D64��7 �!غoy�u���X+�1�� Q1�3r����l�)���@cm*^7'~��z�כ���6�#����է������0}j�HB~̡P�wL`��]��%��o�Z[-��$�m��Qv-���A�|�ٴp��&3�m�/����ą�����J���\���V`����e���ڻ HD������PЃ���n��� �Yn�-T*ᐦF�^o��_���	��زig�ށ�����>5J~�����[J�<|�(�?��m��(�ش�=}j�}q��@�+M�8q�33j�x���a�]�����0�8t�ZM/R�a����f��in�^T����qyR��/�Aς�h�'�?pzɅ�1�/!�-�FEw��[K�B��ü�<���0{K%EO��܎�ӳ�. /@п��ds%�--�J����(�sP�h��Aڢ�	��b�k�y���I9�⵨j�����CM}�O���H<5��j�Q2.O�kJ�Φ��k5Eժ)bCA�&�rh�7M���"ժ�ժeT9�k7���HX�-S�V��[|Th�ĩ��$���'_��]�^��k�ʎ��{"�s|�*ބ�m��i�+��߳�ea��ǻ<g6�����?(|�hTB����	cں\�~�jd�Y]��>�"��I���+����I^g~V5�B0IY5|�ԩ���ɽ
�.�g
E~VҺ�i��cr"�AW��Bf�dT�����+�?I[H]��"�i<\?4��� d�g�T�;�Ɇdn�q,�]N��'�OW�i�m6fbk�o�/��|�}D�ZH��0���>J��f2m?'u=NG�uE�(�wW֖�b�Q�	5�2��6n��mx�E�c���$K1N�Im5�?R�8,���^��dK��i���g�)mR��d�4�̝���������S�ͦ�T�@���Rw�s����㥃��ǵ��>�A@��m&t���p�^���\���䇱w�vD�^���d.8L�趨!F+D�g�&+N�r͈�K�2L���)���A�!��A�I.Ąe@H���jA������X�6��fC�B%�E�� >�ɏcǎ3���݂�����I��	�u��YN�2z�0p�����<�Epv���h��$�����x�g�q�gQ7@"�g� ،/i�-i�G�Ѭ�0=u�؜���#(�<(׉*�iH��I���tfCĸ�yY�9+ӚU�hB�I��k5��C�!�J�������"�)��(x�VA%�
y�=}�?z�8`����=��o��2L*e0"�@�{T��zn����>��?�ȯB������·��ҁ��D��@fC�i��+jVs8w�v���.F�p�]?��?��NO���[�n�y睏�����G��vp��q�r����%'R"Qn42)����O,����G��\>���U��5�P��b�r/��+W H]���[��ћL�B���UTrk��3��En6���,
��Ȯ��*�K��b����R-"�X�����j�6�oA:WD�B���H�4J�4�8�
U���MU��oaph#�[��4P����7��M� ���;�Q��	�A9x��;�ٲX�����d��C�qP��M���W�@ ���
f^<���<�����!��(Cf:�6, ��Fʐ2ℐ���l�ѷy׼�x�ůE�Q���*ʭ�I�dҫ���cS4����.n�"ޖ��F12ԏ���ka/�aP��<��Ȯ�ėd���5�y�(�'F�;Oe��x��� �����
����M�BؑBϱ�l���`
�HH|�h2��q������
�Y^+�!�"�K8���-H"��)m�lX��4֏���(8|���p��]�������Y/��O~HԶ�۷��s���h��r��r-�2
�
��E���+8~�<(��s���ޝ������D�hz�b���f򘛝�����&�L`����ݡQ7�
���N �@����:"��l�Ǿ�;0<D�9<��G����*���-c�ܶY�o�}�`i9�^:���%M���� @nO>�kK��12��9g��c
��7���*6�Q�3L�� S)� �KDυ�����i�1ב�L�:��W�c<\9��"�$pOS�9���-�zzz�"GytD<ja6*jf8	�:�a?�׫��|�݇b�"��j4���RJ�TC@�G��2�ŃrBȽwnn�j�d�&�|&��¦6Fr [��F����a�T:���'M�H��-��P�T�(��؈�Xt�Z(9�7SkY9�*����YB�*��B��z�D�6���l�l�} ��F�^��X�>���&�����N\(��6z�G��T)�̠7���C%��Ȁ����X���8�y��>YHFb)��E�VK�1	��;�~0��d3�ω�챙d*g2�!KU��j��]��{EL�,�#�Z݊���]�s����tǡΉ� Rg�稵6�,�����}G�E4�41�
��0����!J�4��3��XSf�o�bJ�tS~���2<�ʟ��{��ޥ�r6��`���}:�Y@��V�H*���`�H���Yi��&6#�ߧϕ/�0?;'����(S�qV%���)�8�0��tO=�<�i�39�<3b�}h�`�F�$S	�$��ƶ�Mص{�m�d,2�]ON�I]M��
�=!�I����ԩXZ_(7����9H�П�U��
"� ��FԚ60Đ���AQ��Q{��C��wo�=�?�pT5��!`����0������2�v��x��g104�-['Eu��3Y%	�-�i�M$��-��M�6iҮ�{G��k���LC@tJ4_Q�l��+����oֱcs��w�vZk�:N��JCq��Tj��s��R�_�)��k�ͳ��&����a�8�:�>�� �T;GBc���-��y�%�p]��K�A��F�y�j�<�ٌb��D����n���ϲ�נ��Kg�L�V����Õ��k�|�G�}�[?��cso`�0(�̅�iW�M�ć�w���u
��җ��g�{N�������Ǿ3�Ƶ׼Q�����<�pƖ3�!E���6GP�z��K���T�a5��(j_��� �0��8QTHq�ڤ�� �1�|[(����"�����Ԕ*��t�i��v!?���e,��`��14�VL0�8��p�O�1j̍���^� �;�Õ�)��墧��dڧQl���TC:�D�h�;�bǞ��
EP�3�(&x�Dt�IC�0FZS��X��!P@V�pr�h�)�a��oq��JO�X���x� j�-���P23�������f×�iVT��*'.�"6��n=^`h�V5�.� �fMA�VQC�F�
 9��l��r�%�*�x�it ��:��GctT�H4v���<%�}r�I�;L��W��zӧ�����TO?��<�h��+
��B�!�=��h�E?�99��vn�P*B]>/��6҅��#�,���Mڗ��Vd(!<7N+������@_o�������x�sz$%�VV2J��3�b���c���Pss�k�㒋/@_��F;Y��k���i>�Z
ʛ�Y���G����c϶1��f�U��5��e�o��)�10:�3�ڧ���\#�9r�$��2�79����B�EX�U��=۰{�V��$�=}z/�t��Hb����<1�D2�&�gW�cO���'��GOD�SY�j�XG9�������_����
Ł@>W��\�"6�@�XF��Ǒ�S89�d���vچ{���R0ds�P;#���d��5�)�����*��bU=cr3�S��P�1�����Oaa%?��Q"!:��W'�ǰu�V��p)�
�����9<���ͯ"�@ 3�d���V�@����>l���5=3���9diL������t�����v���}ƭ3S�L�e��B�G�/>�uC�k6�=V�s$*hsc����5dҤİJ��҂��.b�7�-[T�բ+騳KK�9
�Iu���#�c~%��E
���"�<�����d��8�l��̊8豈Ec�M����A?Qܒ�x�N�h�k�Ƥ�����=�{q��I4�2ņ��zE�A����	��"�T���,������x�a�S=ƴ����4(:�"uv�k�M���0�B���-c�-��5�X7-
)���t��y=(WK2"�z�N�P���c�#�t�H�ؓ}�mt�Z�R�x.������RfU&iEa��x):ޅ��CZ+�]�WP�D�~�6b}�<���shx|���D��Wã\���E$�QL� L��ty:��*j8��ľ��B�1E�Ͷ\��8�����"r#r�
1޼y���,�Mk@�i|�d��Kjb�mۆA�VuC{4֟��>�i�3��.KȖ�ZF�͢�B\?��e�p���1&cQq�stn��=?�!IU��'�������Ө�f�ם��F��p�����n��z��N�[n����0:4�5���82<V�֔M�""zDX�p0655��6d�j��{�Msh��5���f�Z섞t.'v7�z�k����s�P6�7/.̩����oG��SϾ��'fQk�4�a���N�Y���q�2�5/Ǻ�)�ʚ��k�����e@�:<�P&N���ɉΰv����K��E40�Y�g���8���h�aW���܊@@�N��Vn���������?�����������Ǿ��#;��;w�?�+���ܳ�7ЛD���,��=��� z��������E��G?����V���A�0~�Cƙ;����^��Wa׮3�wיƻ;JI����1C���O�ŏ:���X�%gX��T
B�M��:h[K5�hŕ��)f�]��&��7�1ݼل�G����U�x<uQi����_Y�@2�x ���9L��
VfO��]E��E�����@�\\�?��/erI2I}�_g�vn�w�K�l��R�I�p��(v���;�D�����$��JNt[
C����0�u�o�y*��D���~y%�'?��4�U�z�QX�`��a����k���nt2�J��~���-�i'�dq��/�M|��w��[~�:�y޹X+�1���L��"U>�6H��27qM�h��&ҏx$�T<��TQ?06ڏDԧ@��y(�gW�92��j	�f��y8m�7�X"�Mze-�����,6�M���/��X/2�&�٬�L�ϥ W�f=�(��܆�۷"��O��k�^)_�ca-���,�L�b~)��7�h��4t�fSB7�/K��5I}k`p8���&01ޏ@��%V�(�Z��V�Ea�o�z�$=�䳢�l�y��32�\f1ST#ݠ���F���k95�k�Ul�2�K.8[ƒz�:L�b	�J�b==��w<:8N��� ۷��̽g���]�y��6�Mo�2+��|u��AH BHhF,��a'6��;�_vv�O�΢I�Fȴ��խ6�ږ�Y齻��n���Rkbc?|P�tuUf�{��y���1a}��U*�O���<���(Vx��e��.�>��o�#�E/I$��8�O��MЇ�zq��$b]Q5x|@QN����*�ϯ�0��!��'�v��az��Go,��G���?Op|.�YzJ�$̻Pk�ƽܼ��2��!�xV&��������m�7��5���	�%}N]��maI�<n��	RM��*޼z��օ��E<�^YJy��������� ����u9Af6���*^|�g��_G ��ˠ#땼B�o�z���jC_'b1���VW�y{�[��4<p��N3�!b)�������f�$&�A���I��^ش����X{;zzz��̴�E��1=���k����mayiM����@ �����p���bC�Tb�h���X�_�����(�X���(bvu��Ϋa�Q�{U$�dWV�T̝=3��[.�RP��rB8L(��F�g��4�W�â�}*o(�h��K��t)��QV&N%�B�hݝQ\�tgO�#�,��/���s�:m6js�˸7�Z�N����(�O�J�3�'>��8ԆF�)��6�I�m�VC�ϭP,�x ]iy�89��NŉC�nAOċ���|�G�䲺���d^OS6e�ff	�6V<�`��f�hpQ��4��)�䆉`n��PK���0iKC�|��nܾ ��=���hs�M�\I@eK�2�	* U��80k���Q܂q�L���cT泔E+%&
�lf�0X���=�]��RX_[F6�ԵB�T"q�?���.93�-T3�r�	�ǩ��̻��悹:ST*H0�Y4@��(��Q�#�ΠQ*i[jmTQ`N@>k|D�fP�Xյwt�^��Ck�����������i��g����2ٶH�~vj���T�(o��ʙ�4�4�����p��n��7	8~��$I�,C+a�<�Z��V�l�f�ͦ�"���R�?ӊ��w���|k[q�͗���w�Q�sJO��������Lp�h�V�b"č�������uS�7���s�5I���q�Nz��"Y<��%btI�UE��{O/��(���GW(7ٔ�����s��ĨZ�չ���S������3J��l����J��+�L�������#�����MO��(�!h!�4����B��B�RF�PB:�eeww���?!���ӟ�c�����yV��'�NN#�L)R\_�E9y����X��V�O?�A�T �\3��#�k6N�i4d1.?H�]�7�49�`a�u���
�Xw�n%�EK�&7�3#�0�^��X�Rhr�%�H�lb{}E�����,�D_��C*l��k�iza=�.��'�x�cxQ�]cm�~Db������,����.�%jr6T���)7�{���5{k���eQ^�|c���v)7�J�������\C�Z>�:J�U�MۭN�2ؙYFb~H�57����2)�\�����_͟�o&�(Cz�4j�ǯ�7q��i�g�j������tRAuMZ�:<�8=!����XG#�]{���
賶Z�(�rҔ�(�_\���v?&Ƨ4��2��Z�/h�������p��֗6tp?��#�SJ"���ں&����Fq��	c��z;#P�O9��&.i;�)l�'������#T����~P?�W�.q�,�jeDڜ?1���^P6[��QΕ������E����0vlH��� y}^\�1��k��N��P/8dB6�w�P�o���d�f�|frO�@$�F�d��Xm�� 򭳽�Qjn����lo �օ�!�zԨ�Sx��Uܸ=�j����Ń>BWW�}�c<H%�(f3e\�~_~���n�??��� �N&)W�g��1�����T�.؜>TI�P���P_�������I	|@.SE�����b6o�4[�v��f���~�ʛ����V��x�����7eG&��Z7zw� &w�h���<��*�-�����+Dwg�j^1�ę�o_����ؽ>8�,L*�
�1:ԯi#ϻt2!���U��9��+��W�Ж���j����uH��O4�\����N��討��ܸy��\� N?j\r2���|7�o�{���Ґ^JitD��XP�16�/�?S��B ғ_�Ϣt�n/�:,.�����X��B(�.��ԉ�ho�p@��(W�DKu8<.dJU�mm��9m��ǎ��1t��(�ٕ���5��%��GQ�rBgP��3�o����S'd�.�/=99N�7�s�S��E&��'[���3�2���RX������"m=��RH�Q��c���(����<�F�`���t�Fg�ω���No߼���u5�@e���6���!p�]�~:,�\Kr��D�E_�������J^�ܔ;�� 6ŷ�R^�V�!�v�!8X[RR1�-�U���
'4aeƟ���?�J�J���B6����hN����kV�4�*�$=1M�L�T�<p��K�a�\
��[M�Y���l�TH;��s�,��    IDATŉb��C">����5�H�����K�l�!�E_;��JF�cH�
U�
W�qq[���(R�|-v>��4��x~F�t9=>��mh8H1��=���dճ)`���2�e�h0B���K[4�acT-��D�#�."�Y|Q-�	y�{��;����1�A���_������/�`�PϢH(�����!�T�\[��a�nZx����5����r���<��#L2�J�^\1�jn<Z��P.s~��:���x=����t�?��.>�g�{_��3�r����v�O���ϧ�G������6@�ϩ[Bz׈6�S�⽨�	G>�$CV��f#�� 
J������	^Ǖ����]��,��dP]��F�A�����J���h ��Q)��ޞ��_{�3�����e�/\�eE��Ȇ�/�����?�BW�����󟳝��jZ�6�	ݳ�(�-"�'ll��4�����D6S�����l��?������1q|\F.�Y}�}��� R5+~��
���Tm1�8]C�P�#։�#5��i�S�\uױזB�D�Q�G���S%���P���!��hj�5��\Es�K�I�XD�i���J�T�z��,�/`mq�tN�;MWҞV�:��s�:��}/*��._�ɳ��׏D���,6��J-�����pƄ��� ���C�!�*&M��o�2��y߰
�ƕ��:zn	l\'3d��>�]�
�r�$����YY�va!���'����j�|C�	��͛��fB�~˸�d"�Yl�
"CC��'>�s�?���!�6֐����uܾ�����vc�hBA/z�06؍�('����m�q�|��^��;w���D080���Ǵ��ح�%_�֭X[�c~~;[;�����sg���&���+kX]����^�CS���A�t�F�)�zN�O�b݊�����po~�IN�c������N�e���;��]eǄE��p���f��p�>ҩ#��G�D�8�$����I�Ӆٹ5��ڛ�h����/���k��.����5M�ؔp�BC;K�t*�����pj|	1Y�l��#ܙ]��^��1�:u
�v?�i������
�:&''0���	d�5ܸ{��.�0QD�N�O�%���x�{C8d��nJ��\��;wp���tG111")��Nb����R��3�g�dC�d8%'�:*8y�S�`t���PW��א��sT��F�g���� F���3��E._��ۗo�q	�
D����h�-cjIŭ�ӄ!=`��|��c�=�a��$@�#���d�@��Prce=�;밺���9�*az��c�2�J�vx�H$,�+�A^�	,�3������m$sd�wj�n��:d[ma���K��?І@�`j��������puh�����&gܬ�p�07�%i��U�Y�g���<��%tF�ȧz���zݚ�Ո��e�u�n�f�g���:��W����	���#� �'��*)���l	 �ˡ��&���0wo�N���sgPB ��p����Y�#�'|H0�V8�� ߏ�N�(�=fQJCe H?�=�K&Ӓ��mJZ�v���L	3��1?����}�1]'�ܑ2{&F�1�ۉ0�]ng��0&K���9�*���`f}��Fn �aj7�_���id�K�KC�7�\�9lfZd�w&a*��І��V'���തDĶ���ZE�eG�׎�YI�P,��Ӣ#U�	�,�%i��l~��aqY����|nz��,�V���Mɡ
s�r���|��&l�67�`܌J1�*�!��rU� L�p!���>*%�ahm�8��7������O~�d�{�f�S(�U�Ѡ���|;��&/�$�7L��
�,��8�in!i�Đ�����F����A�X@��*��5X+ ���jY��);(A�ՉP���n#c1�u#ݡ$�gn¸!(gS���o?�g������5�q����/ൟ��3�������� ����K�Tƭ %]y���C�-BY�P�b�k�e4��������b��6��Mn+ݛ��N�m�^ÓO?�������Ƿ��|�+�h;�/���	��!)�?���|����[��&ZT�}H�FN�;�x��>[a�	����$�)�(���N�,�M���!���Mхa����g�$g��#���(�U�QJ���?RJ���O�ٷ��~�_�����i����Ǿ���}�n�>���_[�>���'����� �.�Z��c؊׍D���_~��'5���x���?{�4z�{�R$k�M��D��\�[x�'K���/�!(��p21��Ҕ[+F�U����g������7�%m �����<��9�2�J�l��N�J�."��"CP�7`�U5�aHH%�j5���*�����wy�=�HJ3��� ¡�X�,��t���(���'�8bL��!7�`���UB+fN�>忓����Zaa�rj�x��f�z�b!�ٮ���kY�f�STԹ�ce��iH�����V�27��a���DJ��.k��j��\x-ِl��Z�bB�!O&���Ga!��}}��G?��O=�d1���u�Kd��-M{-�8?#K�LT�2�GC^�t�K*D?��C�f�I����*~��7��ρ��:�c�;jH$T��Խ���[7fD����(\��a��Eo؍�O�8��]x���w�ڔ�&$�<�#�d����#�_XG"]����TN��Vc�f°L@�}K�]a�����U�ְ4����Q@,Ȣ=�É�R(��s+�~��::p��Yt��! �._���u���1�Ƌ|���E[��σ��Mb�� l�M?���=ܝ[����BC��N���X���9$se��a�#�P����}Xw
�ُ�%�������h}�BA�!*H�������M��GG����#���/�:>�lE����#'H	����@�g����06�	���u}�f��~��,����I�p���泄@ȇ�''1qj��:~��elo��t�t}��+ņ�Ԗٔ4�T\q"RFoOF���"� �B��F�*��vP�r `��;����i"U�W��Yp�X/F{� S�������_������hu=��3��;ʁQ(�|vknJ`�.5ݽQI��a��^�$4�o`~a�lEÖZݦ��𜚦�1[,���V�-�����Ŭ�MadЃ\��<"V��(�8��ʐ�Uʉx�qz��~iyC�c�x�H]60�(ݬ&��,�T��e�,�*�����߾�ޮ^��>��6�κ\��������R�*�V����+���Q�wj���Hk6�,���Y�Ͼ���ϩ�? 9�����p��"
5�HM�Zc�x��菅Q��4]��:�t�XhJ-�\�k���b����aW.����*l6?�.n5��{$i)��f)	F�0�^x�D"���)%i���5�/I ��]1y"|�C��xm�Y�ӆ�Q�k��BJI�J�o��Rg�������HS-�(�0>0n��Ӗ'̜{�	�n� I؞&���=>�H�
�4�%P�N�h�!�|�R��S�!�v���t�u���������oG��ͮgu��':��Us���?��
v䦟�4�PJc+�P^S��X�60�2��HM%=���=7�p�����������bwK��M���r����L�Q� ū+W��Θ�ϖͥӤO�������"J����w��~�_�:q�,.��_�"^��+�X[�$=�cbbB-�A�� D6�l荴��>D

@���2��țB�dʩ���ූQ_�'�C�i�г�8���k�F[{�ȇ�{����������7��Ym��
Ez@x>�"���6�Me���3R�Mӿ`Hqv�\y~J���%l�9P�{���[c�'"tU+������ ����`�tB�}&.���%��x��M�u$Շ�-�.� >k,�����O|���|����~i�ZY��?|�/�ݸ��������'�ddƀ��"�NvH��F��`�����y�[��/~Y���|泸x����)�|tx�PP�!��"ժh8m(Y�(:l�ދ+��．�-��%,�9o�P؇t&!|'/`6��H�`��u����`i"��Q����5x�4f�u_UBF+!JCH�vb
oNL�+����e8,L9��"�ͮT=�*qZ�Ց+du�p��%CNs�0+�����@L]T�o''�l��(k�⪐ &/��F�qS_ɡ2�s�+r��������?��<l&�� drm���*�$y}����f
؞]���"J�kz�_J��ʅ���A[y'�Tg�F�!9�h�Hk����}��XO�}x�=�F�Z�����J���CB���6M�NNA؍T�
/��d�m����h�� �r]�m��O��_��̂��S''��#9d+j(��X^�����51B,���;����G�P���v��P������@�z�([�RA�q�=����T�� ����v�2�7\�X9�3f��x��sj�T���I�H"�{�(��ۈ�Z��ccm�~;ޏ��!D�V(��W�I�ԉ	LN�5 S��*z�9RX�s�;�0o|���N<ya
������,�7/���^�I�mp��	L��9sK��ב]�jas{e�~��mlmH�A��R���>\�x��$������z�6���Li�'��9��cCGgT*�4,.���\�yՆ�����>�:���Y�<1$�>~[�9\������G.�l�>�n�(�J��`���&__���hH��e ��&����dnK>� -ª�Doobr���&��a�����į�m��[3(T��J6�Utw�pz���vd
%�W�74�f�*ϯ���9sFM��AK���>�A�<�=�88-����p
�544��j����t7o�be=�
�r�M0��� )��׭��g���XtB��ݎ��!�>هz��"�B^����El���X������α��Cܝ����&��Gp��C�:��{x$���
R�b]}�8���.*nm�q�˰�\?6���6�~�����*��_���>�6���:1K�-�����ɉNd3>���Y�C^D�^��fNL	v᣽�s��{�,x}�����-H��Ś���E\�����3�ù�����)DCV�y]��d8 ��&�q�{�(��� ˦��*�ݘC:]���#��J�Z��W�)*GM)�M>#u�0ܭ�",t���Xk$�FB$�cS�ϳ��nK��h��_�׆��Y
�@,����P��MA��BF35�w��>�?��Q�l4bi0�jD��K��j���)���v��NO@��i����0o�XD>����$h�k����%��v���TJ�`3O����P�
���9m�4�.Ր�a��$���"�X���!?���}����af�!j�+���Ϗ�˃2�{*P	1� �
2�8�U %U �tk�s�͝��=J�!�C#�
�#D#~����>���T�:�ޯ�|�+��~���E4JUX\v�={�]����h��+M�2�'}��:Ww*�M�MM�9���l~�&м,鰦��A��4����^�I0va��0>���~��(�k���=��~�y�m�T�
�ͤL+'���Uo�b�\{������V)���i�4�V�L���P�H�67�8�<;ʵ����!pZ�Y<�T/7ݽ1���X2؎������i�YɎ~>��,J������>�����_���F�����_|����i.qh����@�/����F?K�͵����ߏK�<�@0����÷��H[>�[���$VW֑<Jall]mQ�䥫x�󋇙Ӎ�ło=7��?���~؜�Zx�[�t�?�U�:0�'�\"�/)I,։��Xx��UhX�Ӧ�I�m�.(=^eN\�nbp�?�|�����!�$pJ�鉌������n��j�}x�P3ȤV���ժ�5I�QѮ4��ć� nL�ltlV�,�M*`��E���7�щ�1�P\�	�G9�a�.<J�x�rE�i���E'r�"��
�X��|KW�a�� ��l�q���0l���jF��������T��CpC ���ߋpg'~�Sx���B�e�F|�\N�o:>T�`c��|��AyL���˻� Z��c��`����v�:b] t���č�E�:ur�>�P�!B"Q����X]�UcKiGԃ��v�u�����pa���ʠ����I<z���c��73�	����pq*ICdX^�cii[�t��T��Ԝ�rZ"��[+F��s�a�KՉJ����p�3�J#�F%�X^�������LNM�P�OK�]��l����eI�
�{�~_���@L$��|��W���Pʧ��Cx��8N��"1���T���Gow/�(6v����/�`?�k��I����~LNG{W�TU[N|���p�<NM����h[4��l2���Awo3�	�w�Gp{\��VGoč�'hp�@��K�zk�o�a+�Ն�Y$^�M"���f��=����m��"����gC��2'���eУ�ѕa�|D	��	��^�v����a��R/1|yI
�eVV��qgukH������ ��;��݁J͊�dF�-q��r�12܏�}}}���b}s_zU���k�#}P@�qܬR6
G
G���p��"���H�Pf��͉
i!�a,TL�^o�lf�#`�����\8;!�%�ɣvwv��0�T�@&����i��S#���!w܂t��0y��C~�}$�n�U�����'N���p�2G��r��R���s�$!�R_�v�3�{	�P��
�١^D�m�S�_��d�<%{{�ً#�+bp�}�AT+LǶ`}s;;I��(o"$��`�fL�O�>��W��R��յ���Ur�k�+���만��],�l	����Ї���'�pvz�7�Vȷ�JTe��ys����	���΁K3��Ŏ)jLc�$�fa����S�5�龦���D�V�!���gM�����PC���`6���m%�Q7O�7�9���Yg��ƃ�s"��E¬5�)��1r4e[/�JW����De��B	�۫�)�f��Xb�R�WK
$�~>�q!t��gF0��ĉ�������6ko�LZ�*C#�ڰooo��`0W8Ԧ)��z[�G�x|�3�Kj�eifJ4ͤ�7ZFt^#�B��8��q���a�3�\�6�?����h�S��9�y��e	���#}͡m�ڜ�{H"b�������O��L������~���+�bee�<}u��< �c�k��:�;$)�5�<"���Z�M����5�5���3�tV�����d୛?ϯI��ֶ`Ʒ�±�Q|�����}����|�Y|�k�����Rɸ��ҡ�%``��Ɛ|�&6)��&[ͨ$D-�s�<��
�c�D8w8*"_�!�LL�c�M%�;���ys��GT�<N��v�6U���M�g6B��m�����������_�5���_�����^��'��z��O�ҩq�}nƴ�4o*�s,Vmv�wv m�������ܝ�������޺yG	�;wcC��sm�$ZP�Rw8P��pX���߿����6��a�=�h4�
��ڬR�(¾��}�@��|&�N�s�O�|�؝�S�{��@g{Tk�%)%�0�ީ���|2�j��DU&�r"C�J�alN���3M����H�k����6ӌi:���a/��p��Z2ׅ�1�36#�y4����-��D��Pi�%}~�gq�ˤ�I%u3��n\G;H%�D�``3��/��X�v�6<H���66	nd�X�����e� k9/�7���A��<��]�@3�J,|�����{Џ��z�8��(;,�9<D*�7Rŗ�K#�knd���l0殪����F����������ԗ^~[�+r��z�!��~JU�88�bs���{��M�@i_gcc}G|Hd�X�����2��I��v�x��i���g�oyu7��Ӵ������"?P�Ģmnn��1CY&��d��=6�${��(��6    IDAT��Z��=c(�����g���ˋH�������iP�i��V6�T���crbB׻M�
�ٌ���p�\+����a�8�mg������ݦ����`c7��^�V6���|���$����Y���]M�'G02ԧ�7��Q/��S��"
Ӟ��XトDB2G�r��kWp���� ���S�>5�4�%P*�5���ch���Hg���},.mbaqE����8?���&7$m�'�꛷p{>��ŧ����R@9��.���4&{A=��<Ә&L~='cSq��o�hѽ��%W�#�3�(�|�ʠ��2����G��簳SD����D���@oPj�-N/�9\�ys󋚸3d���ΝB[$�	^�b�V�s�H&�:�-2�k���"����!iG���faqe+�ԵѢC2�fւi�MC��N~9�Jt�KoC���h�����bVXZ[�R����:� 1@ο05y}���lXt���a/~�p4���^x�V��d
yܺ;���+�t�w���NO��G���2�7v�D1>9����|kIm��ߚ�7�y�sە��k���!�wG�Ig������%�r�:y�F��k�X�XZ������e�M����}z/�-=�z�"4�E��m���Y��"��4�q1L�Xwq��mg�5l4@�jJWgfȩ�S�vA��Tx��2^{�&r�Qjhр��ʴT*\�Y�j
�c��?'��D�kN煫
� 1[�'�8����t��,hCP��F�&C^�f3�b�9eU�z3��5/�̵�:l��ՖD�u���)���_xq��������m$CT��`5S�R�R�b5��-h�	�rf,���_��ӓ�$S��ڔ���P�n2�骻�N�!�D�mh�`�@�_���|�y������@X�5��+`��+���pSρ�H���v����J�<4:��g�<�4r?�G�%�v�e�V ���_C�#Y�Z�)��K�����A�\Ѱ�4��$l4���z��<�^y�4l��2N�;����tOB��&������2���Ď�8�{�@<�G|���!�AWW��	6����z�2�KTl�0E���(�ğ���C�>�ׇg�"���o�ƭY�J�d:a�d�S}�[Z���(�*T5��V��.��2�F뚓쎅���<�(���h�����J�-k�:�+e��Lz��gho���䐚�}meU5�6z�(Rzd3rT�c��J����'~���~�/~�������翈��kW�N�?��������C�N�_��GpfbTd N<-V�M+��T�R7ig�T5�,�3�l�����^�)�z�2|?{�1�����
��|(S;N�É������o,����ى�4�c�A�p�׆�X�V���]��y8�^�Ua��m�ڲ!���.<��Qb_4 ���O���)�|1�:��1W�$�n����L�~?�*$l�`mnJ�7�Z�p�T�=><@ü��C>��pju�*P��p�'���Ѱ�k ��Mg��4�h�̈́�*�_0@�پ�\oQ�X�v�*Cs�������>��-V��9���&
[{(o��!hm8M0�!�!��_���/5�T����~k5&��j���;<�'��^L�;�L��x"�l���XM�śSH9��)�4Jē�Gji��T1趢�͇��>Cm���d����Z��r��'.���g%�� �,ck3�����]~/�F�hj@�= 2��֮��G�I���pf�8�>���7�0�����ɓ'��$�0������,�V��į��^�!�3����:�&��u������h�,�x<h:���FW�=݆��U��������Vd�<q��C��@�Dԕ��-�5�H�9e"4�͵M�8�d`?�C�w�7p���%v񺶠+��vL���������=��:q��iD:���Nf��v�6gWP,�1�é���B�V����e?{�0�׃��zcc�җ�Frr��M����Gpb�\���h6�����W$�ů>v=�n]?̄�����E\���Lن�.R`�	ΠV6Ee'���d<a�4��7������㵬�X�2W���v*+]��B�u'C
�x��)�#�2I�����/!��+L���al��Fb�Eð88�p��],.��~��ڂ��n��԰p������;8�?����H?eE�h�R���t�� .	�7DO� ��+X\���;���;�u��ǉ&�$�H�۔=�Q�\��;�T�IhbM�1�(s�S_o ��+��EogGC�*�3����[;;���bd�_�E^�2��-`u�@��Xg7���b�x?�n��17�$:�"'ϟ���)�H��6�����7�!W�!���Ǡ��NL��O�� ��#��H;���ҥ�8�'�9��4n�^�Q�<�$6A�� �u����qD.�H�#U���'�xH�4�͹<.��x᧯cviVg NoH@nR�b��� ��Ch�h�p��{��Nh��I(�=n���"+�Ԡ�5!��+�t}������R]�&��Ak�X���͢�`wy������*��8�3�N�3��K��-9�f�e>_�y����8=C$~G�c��m�FlprLg�An54��+}�\��h��r�v3�u(���f�
~�Wޅ}���h"u��<�M1���qD�"�������8n���tbo�������o=��e�!�y�P�����j���{�7d�6�k�f�BH��kq{%Tͩ�	+B>�ڸ��R*	{S������@4����Ã���4����ZS��-���?�G����� <VkC�֯~��x�籲���=�yGW�NMk��a*�$�pI�"e0+++j�+����狺~�K��c��l�l�]T��Ә����a�����Y,/.a;����5�/=�?�>���+����n���6ů�'iS&*�ZZ�y<�z"`�E�C�b�(�T��E�UC)kW�M:�-����Y�8��0��k�t���~OX��pr G�%7%{񸨔�YГҬ�4�̱��s(��>���>�������i4��_����+'������x��ⅳS�����}��2j��y��d3P�^��bӃ�:)m��k�y����|�mqo[Qd|h0���F���~/��|�Żx����!���2 ��4�`g{��!�>;�ռ�47���h��cM��!A��:��Y�i�L)N� �j�Qb�ȋ	��f5�Q������`2҉��k���F��@!�	������;��o6���dh:T�z���Hē8`�r�`̵���ʼ!3�4�D���:�:ۢ2R96<��#�u{�S�ce5���m���P!O�ON�x ����H�!>��)CĜ����}���7�C���
~s
g:M�0�����͂��	��G?�c��8(d��L>h��'�����A|`jb�Q��v�TJ$ a����%��#��r�|��uM~�.>wv?|FӢ��Cd�5loe�4�� ��۝�ƺ1:C$ꕌhe�@��s���ՍsS�:6L\�8��"{�(	�׏�X���u]%�Y���J�}xT���)�_#��4h�lX�Ħ��5�a���R�c���!�}��v���D"'��XZ<D�(��tN:���~�	��N�kV(�j44)fS�S�@:�����p'Ƈ��E\cM&♕8f�v��9��z�q[��ab8��'�`o�03����6���8�:�ȣ�102(�7�D�޽uG�}�����$=�� 1dus��y]�3�c�x��:L��raq������ǧ�����������M��g�K�qvb����;
d�e�SY�[����&≼���(7j���W�z��gpX��Ճ�'���2�)fX��͗6 ��>6��FQyv��5��m��=��ް
N�g��bn�@?';[g����=8������%�Wn�`ecK?���@g[ �C���0b���o���[wQ�������8��&`���*#�I`aqV��P$���Sh��JJ��r����D�0	�7���9�x�7�&]��e�&�9��o���դ��&��۽�.���
D��[wxt�x|�K�*N��V�-M,.Vvv��=�F�B���=875�����4��𳷮k�~|z�/�E_wX'Q<Q�ݙ��B3��eI>تe��n�Y�܊˴��c�x�Ho�|˫{x��%�492,�vw�Q+eqzj�ΞBIX֪��ܝӄ��^�I+�i�{	���M����֋�գ�6��ͱU�1S��lUX|p���ho���Rg�tⲞÒA�Q�&K�}�󠶿Y��QMͷIG6������(�T̆`{q?{�@�����hZ��rj@9�/��j@zSf|�!���&@�$$xϞ�t
6�ʺ�ܔ�z@o3L1�3"�3Q��"���+J�H�K�<7��%�k�^��� ����p��Y]W�~5v�C�,X�n��nL�v8<���������G/���4�v�R�ai���2�:4�^�w��𬠜��:����n3%>�a���D������B)��@��A�����#���N�{	2D���j (s)����������tm}_�җ��|��r���zǍ��a>����V-�"||\a�-)/
�s�G��=���3�A�M���V�a-C��0����w�P���kv����X�X��G/�>��9~L����o���޺��"���-��7�AÄ�E�����ͦ�l(Gk���~�\+^�u^l��	��T���R������ZbTK O#�^�يЯņ���=�G2nyy��z"͍~�ԩ�qy�!SM�>���>�̿�%j��/���׿��T.w���㣃���b�S	�&	*��*�-/��?��C#hF�wx�L���X?|!/^��x��˚f<r�a��I�Q03��EZ�-���.���Cf|(;j� @�S%G=�����.� �9�+P+hb��)��S>�5Q� �[md�MK�N��4&�Rfo���ݝ�p�h�����j��2T��W1j��ACfeX,�P�2!�'�I:�6�5�hv�t�J�ԇo8�4%��{E�*W�d��kr�̤�r�gK�)i��cՍ�-�[:�C�'��Ӌ��u�P���c����p�p�- ����چ�A۳+��-²φ �Mؔ
ٸFf����	���_h@�;c!񎇁�hl��"������9����O`����	�'�dx%���V���4�4�.

o\N�؄�Z��3��X_a?������.���b��#~L�Źs'�t�t��s��jC@�e�ZD�-�������j�!�`�8����r|d�����������~��L��/��U���&q��]��m��
��� ��8NW�0mM���kwN��$V9=85>�XԫаX��jI,���-���a���f>F1���twu�\�a/�0J��P8���^�4�)�ΗAgl�7�}�����Y�ŭ{�8̖����������G��<Jbyi��q�ol��3�����a�"fss�����^�'O`r���	��q��,._��U���pb|�U]v�|����O^���*��G��#O*M�����:^z�UMg�O��'?�^����L������\�Y��~/ie���T����0�=J(�������y���Ws�k���)�&�� �z��L##��-Ւ�����
j������"��h�|(S���:�����B�l�W�`ckna�]��j�:8�j׆������z����喧_�*��G��~����~��G��?��.��ͫ����Z����@�\�4���;7ഌ���N75��vEd"�9�cp��]�p��P�+u���Z����{:�(#===���[f���M\�1+
e�>�G:�875���`���ǋ/����m���!��#S(cqyK+����&�Pt1bu��;�q�8GRU�;{"�<�ԣx�l��v�K"8�umV�9��qxs��!��c}x��S����L���.���M$7����֍{H-��b(T��ȋwJޒ:<@����U�����f  ��5�,��57���+*Mj�I1n&�d�M���ޓ�Y9� ��V�+�Ѕ\Vt�؜��O��>l���ML����<0��!6�b�棹9oM[�cA"Z�{�;�̚$�5u��z��4'�V�ߐ���W#�ձAa��`CYʤ���48N�{{:����^���Q��駔���$��b�aDmbc�B�E��[0��5������=�+��		�`�N�*�c�:�RI51
�YP�e���5i�!�U�@X��*Q��9Pc.���B���L��m��I���K��,(T���#mj>3��9n'x�����J!�Z��]���������B�S����/�!�XY��E�?��O��W~���I]�;vL�����5r!� Uj��1[g��M"9��X���to�OT-Q�*��,+�P ��a
�n�B�V�G>���G?b��j5���+��/|�n��~����d�[uM6�!����~�X,FY�rɚ	��n��ٔ6eN��T�[A���fC`��qϞ���a9��<0��t:�`{j6E�g��Db�M�z@D�3�#���[x�K2������o�m�X>�����͂r��`V�Y�y\\�X�9k���Z��^���,�I�������.���?)Z����k2d�C�y��i9����[y���:��9�^څB�#���i��RC�Z�����;{����)�l�,�L�� A�=O�c�Կ��3��&������g�K��ЦL�t⭴҆pw��+̃)���x�.�����2���j��2Q�������s��[7}X��IKvXu��Z�p�K(��+���S$�t��=���:�x����4�6��Ȕp���y�7P˒��!(�f��*L\��U����r^��`y,�h�+f�#O�����)|�����ӓ��88ܓ_�����R�u�6%G�5�|?���)&R7;<�H_D�Q~^�W�ͮ��7/���h|��I<t�$��Je��Nk+"?Qk���ر~�X8ȼ�@2��̝�nn����B,F�0�]�JՆ�˃n8�&=1��h
���+�{wQ�ѻ�FQ�t�� U�W/5E�U۵r)���c�8>܃H�����tևG\����3$1��%i���ѝ�-N>����a�Ϧ������G�rX�a�y�8:�U�-�4劚l���+�'��3�8>ܫ��L��ٹ%M�YE�N`d�8����:�V��$1%!���� z�{u�om����W5M966�_y�1�,`�9=n5���������p+�ukk������
����w=��c(T �Q���x������&7|��$�^1I�E.�!iZis!���(��)!m�Yܐ�e�,fͬ����F���K�pa�S���� bm
�;<�a#^��f�{i���*mC,Ѐ�nA ڃD���._���:�?�����Q~U�P;���y��]� �����W����L3��b{sS�������pe3���}\�YG��LBpF��V{�Y���7�(��
K��Lq���@�ư��6ż�b�mDgg7�,��ҶW�y���`og�Ϟé�,�\B
�����El�;w�ΨO��ҹID�.V��_��{j��Ϝ� ![*��������	�p��$.]8�\��H��z��^��@(�}�x��Q��[y\���{��8��`qF���l�r���0��t}�`�2FR�������YX�U�y}���_� \�����LA�7!V�2�,5���Ņ�鐳2f-�&'�Ҥ71�|�r[��<�[���P�%�� E �����S3�0�hr������Hw;�3x�ߑQ�zzt�Sޣ�>��+���-������$�s�h�\���*�˘���dv�!^?�uE��)@ᚤθ��/���v�	�s��8J�!���    IDAT��yCUv*�����ꔃ�14د GN�w��a��q����>�铓pY��Be*h�V��G�S����ug?��WE���ϠPj�!�k�{��$
�|��߫X������bq
e�r����P�"U���Je�# /����L���S)��2K�p+Iw�h_�e��pJ�
%Vf�^����K�+e����S$s��=�s�H�����5�rK��P3�������`����C��I�VR�Ӊ��#���{nml�!f�̕��0�+��YN�yVpk�Me������n��?�,Ǝ��{A��w�<����)����?�{����n���eά>[y�s���Ys�k"��u��6xn�-pP��g>'�nX�~�C�(��!��\��(]w{%ie�Q�4pV��<�ʥ��3�3!�Y ��oXل;d'Y���MŃُ����~����;����7.~�k���J�~���A�=u�~⒘��2����9'�􂫺F���+�&��_��7��?��᳟�oP�����?UCp顇14ЇZ���~�ˉ�Ӂ��2�}q�]��~Ƌ������o�{�k3o �v��!0]8��N'O��7�F�җ����n�Ԭ�l6M�[���-��ea�cv��hyZ�B!#W_bN�.��������dU�)G�D�7�~�dh���'/f�Ѻ��?;oLfo�А��WC�烝��C��I$ꇤ����7ڍG�z{�G��۰��Bie�p(�l��������7,EԸ���I!Y�|�h"�{����R`��J:�8����|��7QCxt ���`���&���#5C�x3�Vʭ��/�<lLC@+����1�߁��0~j�(���Z����E��x�P�>qbv��G����VV�����g�ctl ����F���x�g�O�pfz������hB��M�.$Q���i�v�YL�^\��[oݖ4)����t�ZF���д9�K� )!p�=�E��a�DP.$�)��}}�7n�aq� �E*H�wQ�0��ax�,h��A^��D,�<'4�E�A�����z����D��A�\A�(���x]2��h�� ���148��� r�f���J��l�*��p��$b��(�����B*��{e`x �h;�.��iܿ7��S$�{��$��:��At+�2�;z�����ۧƀ�{�ܸq�o�F������Ft�3h�����^��x��D��p��d
l(�9�"�8��τ�q���!2�����6��y����bN�m�xj%l33�[Vd�<.���81؏��6-��)�5l䕬�MQ(��g|r�~��`�Lů��6�V�Q���ׁPЇp�'�_{$��n
׮�D&��X��}��P�b�??1���-t��q��q�hf�Z݃�lw㸽�.|)�ԡk:�������w���`������G<w�
������N1���$�x}���҂Օ�ܹ��Յ�g:����7noȀ-iAvѠO=zR>J=���Wp��,� ��O�ы����&���Wqx�����E_oD�$�L_���윶���������N�D	w��p��
�"��n��W�0�.�\zǆ;���itE�!"�-`e'���������=�K�����mtt� U�i�g���0U^����h	���@)�]��g��P=(�U��YE	WU�2�����w��zF��<�!�/s�%�u�>�s����'�03��"1"!�� ��(ﮬ�]yW�l���Z�D�6�H �A&�t�L眫�+�������o��sp�&���������$)�4� 6�d��B6	S%�]=m؜��K���T6�"�G�T59��t<3������jh	x�Ha�q�Iu�i�㸮D�'�J�$�Q������؀�W\���{���]QQ��� nq|Ϯ�.�%$b1��.`yyUt�MM>��岉/���M1��hm��?�a|�GGk�4��P.��މ,���e���୷/alr�H
�
�NZ�k��2Pap�����ň\>)���$�2¬j�hdbG�<�
�^7�^?r#�6\���H-�!��c��f�[,Q6�4�ؖ �����[N�mlP�g�$����#��������㏢�g����˯����FX�����q���U�@YY�۬J̆�����\N�'i��~qi�v(9��ó[�ԙ�d��F���k�^�DJ�5�=�k����Z�����x�/ICƠIRn]���[��qR��E�i�A��9��	��	Ko�Y,Ek(q�[�0�|�wQ5�bE�M��d攃���Y���0P����\Xm���Q�Y-���u�wZ��� ���j�&���Zm�W�(�W�~��7���o���S���"*���=s�O����J�=���g?�	�s�9�x���1�tb��$U�ʎ�q�x�g��+��`~�7��т�.^�i���+�E���*��:T�A�l�ݨ���q��2�7`r�̉�pU��o-`u�=d6oAW����`2%g�EK�'�J]��j�&,��5r�Tl�D��s��&!om�Rc+"'�q��l�{C�Ƣ�]њh��V"'Rq��^�P�U45}���e�e�6��`�O���	/��wUE��=I���LE� �C�:�8t�^��T�,�S���)��p3�cHO� LZ{�*U6[j�Ϡ7^��2���{$��!�[���'���^�F-��O�����%���*�Gn�x���9�����6$��.�]�ū�&�rX�!�Z��w�5n*����&f�W��E6���6�9Y�A��e�9,έcfv��:{:0��ͭX�vAj�70}k�Zw9(�`v�Q��(�ne�Gx1�B5�Ո�������7߼$4.��n@��e6rP�غ�E���?��ݏ`��v8�W���z#csX^��P2�h�˴6����Ƀm۶���H�\PR���P,�B���]"�#ݪT("Z���B0��d��-�N㭷����o�������m�\3��BO�@T�/��n�w@�0C�
1`�8����[�r���V��ъ�'�c�`������)�yҒz��4:r�i�Kh6��bzzV�l*��Nǁ}���֢,4�CE���%�si&g,���j��� ->&�Z�-%(�Y$���ɪ03Bk
8���ϥ	��>X�KR�%��d`�UpYp`h }m2 يg�豴��7��o��k��ۅD8��!�^����e���h�hA��&�Z���-alt\ޛ������D�����i��\��iŎ�n�)�
��B"_��jo\���LQ^/a��H�?ٻT1ǽ�,�yMnW�pq���R��r�\e2�Q,�Žj7�#^�����G��������p�LH�"���[+�dU�W2����{N��]�p�X߈��/HƇ�⒂p��n����K��[3�96%t����y�Q�RK����Ņ5�c9)���8s���nq�47W�7q���"8<m�:=R����WX��éc���䁁��|3KK2�س{�������obv5����U:���|�ZV���
���`1pk*���י�����G��B�d�>H�=�-u^5N&ox<����*dG9j�5yf۔2h���pc�����3��bpx�r��L��T!k��-��iѬFUCeV(13?�BA��h��EA8�q�s_6��j����ӎ{N݁�����h��s�?KL�Z��Y���z�nMH
6��ZZE��47���il�/I�Щ���W�v"��}��6#|�#[[���ūo]��K7�A��ѷ��)���R��m��Ao_;������]��-B+��\3!K#�c���MO���<��px�a���Q�ĐY^�YI����nT}#��	+��S�;J�O�˧���T��日! ]꽋�q��y1���Ht���P8���)��7I��h <lP) ��܌\Q�
R��P��(E���G�Y��<�u��O�C���9��U�188�Ǿ�(�臡�Y����O���t�`Q�R�X�����9)v��K�2u���T7�$F�re����7O��
,N+
d 8=09�(Sd,e�^��l\mn?\� ��*�4L(�0����I��sO�J�g�vlHs���\�8�*哴{�C�������w�)�@�g�Y��|��CO����uƽ�����#�CsqvZ��e^$��L�5���b'�Z�}��O��˯���_|��p:=�t�lpg�>��D�#M�l�	e�Sk%���\�jf����z�uLc��y$7'`�F���v�U�E	5d��q��`j#�yv��h]���lL�����qՌL�E	B�E�{MR��N�Q��h�h��N�&�\���X5K��v��*�E��~u��3�l���FJ�h�Ֆ�'5��T�L��8�}w܋�ˏ�D�bM,�t5�k!��Ca~^�E��SD.��5�<��IR+��W�hI�����6N��4S���MY�B�__�m�`+�BdsC��(�2�=�x�t�PL��$]��5eجftw���aC��+������1<%A&N'7>=��mt��a��I��ı���xr�Rxq*�⛼ϙ�YL�O��pុO`h(�J��X,!���)Z�eQ�Ä��ǌ�i@Z��"H�怛7�ƛ�P����D�^ձ�R�>�Ζ�y��q��^�����r1
yē	ܚ���J�"E�tqK�V����ׅ;�>�kka��,a}m�-ݪQO��=(�fCJ����2:[ZD8f�D�h���022,����.��6�����ʾriy�،F��٠u�E$l�	E��j�rQ�.�7 �ĵ�1����=]m��P���Z�z��A7�r��T2�d&-��r���!��R,z�f�O�U���tt��E�\�H"�w��K�]1����H!��������.��v���O�bbf�RM�E��[d �l"��)W�D��F l4��

�8��<z�8�k�ۚQ-�K尕�ar1�щ� ��:0��mp�)d��R����[X\^A2Mo�\���&x=.���%����� �o�AoW�p�C�-q���H�ak+]9'�\}�$E{�P�Z4��P�\C�b�Ѧ�h��2r��MMD��3MYL�FTJ*=��˚��|��L��S,�����Â��>����=��#�$J4.0�V�R$r�1����u+�zo���v'O�Ǒ�%_cvn�޹�P,'��j�@��w �����$��gj�;��꓀���Yܺ9�R�.�v`��9��ߊ��u3&����a�ce�ݭ��qldԗ��Ρ�Ɇ�G`����N(C�vВ��a9�\�Rei&f7`v����H�Y|��{.K( �.�@ǩ,9��x-e�O$�{��ƹ��XMt5��aPmp���g�& ʗ��}e�,:jHe����hs��ԗ1�
�/�C%�����ڔ�I���h�Ҫ1�â�D�,�*֢��S9
:D{G�YA�qRl��3��M�]�+bQ��O��>(�<_+����3E9��Z~O�É�%���{��	��l�1?7���R�-8,&Is��ÿ��;wI4�<�r��������x���$!wm3�V9�*WE|/�F��w�ß��;��	_�����އ.��\E�E��
��y�u�*�:�"��6P��`u�a�bb�O��RY�w<x�2���<C�7�Q��:��E�yqY��n�����#c��q�/(���$�#l��^�|Y����1#%��������!)��V((:��  f�e4� �l��i���Q��Ҏ�� �j6*2�Q=�+�G
E6�m� >�Gq��\�>��~�:��N�\%-W1l��h(8�cv)m�����QxL$��?l��F����yJ�2jْ�--�9P%���\�;��&�f�V��Sh��X�D9��$2���C|X��%��׃���TII��z�! ���M �č�}�����{�<�3/z�'��nkk۾��U���z�?�H(�|�(�~3E6� �ln�tv��'������g~�v�އ'���bO��ko	z��;���rI:�� �͎������n��Dpv
兛��XG���Bx+co#�:�C0�r.3$��m��#�%2��Z��ps���d#��:���A�����
�1�ol��B��=��F�Oԁ�b��������KWS���|*�N��W�|V=Q��W������&��_ţg�"ŃCw��g>�����h�����bM�͙y$��QK'�3r!P����4ʐ�[U���R��iX��K�n�ZZ#&;Sꑯ�оo'���'�هH&�<=��U�$�U�M-[7���u��K{IN�&�t���σ&���mX[+��w����p
-[Z=ص�GlE봬�G�>�M��P7513�R��M�#���������#�����n�B4����� ����*�M��1���G2Q�+���X<'�Y��)�5��2=���9t}8z`'�:���^�A*����V�["8d@K8��$c^3�̈́`k {���U�9I�[[_���M��D��^�|>yƦ��0;3���6q������`������Qq�ٷcz����"�I7���-lFRB�(�B�f�;���������:�2�2V���0��X���ؿg>�Y>/�G1�z3��Jr/'Wtㄪ�=��-�YR"�-\�r�l
>xv��G*�E�"�R7��q��-����x`6�`�W��s��!��҉z'�}6p��DcI���������}"�n��/
�h�ɘ8�(�p���ۇpp{/�����Y�o�16��x��
�i�����!p��LƢ��A�˫bH��@{��A�\��O�qs|\��L�#���LNnu"� #���+�KF��w��c��7��"�)b#����ElDsbyJ���tsͷ��[ziP���#g��5h��+-��fo@�5E�D�*b�@㝻�I�lwq�X�<���Ui�z%�&�+c|r3s!�*��k�GWlf3~���ɵ�yk.� ��[�[F6�^���-ڇ..�"�N��I_o�4�l��*!m��\�"��'1��b&,��K8��{Hf��CB��|���٘F[���y{�m������ξ��~��sZ�SN�^~�]��/��l��D�F�!�D5P@��sR�:&m��/�7�Et*��9<Pϟ�ݯeH�Q�J(V ���5��ze1��F!l�3/��t�":QC��s%���L�\E&{�ƙ��F�\hA�	�Fb1-����������ɰF�9��=�kK���.kں�BQ-$px�v���>�{O�@2U�&��E��*�t+Kz1�_�wo����g177��	3m��DC(����l=�Ǐb�А�#����B����n�������K#�����J�l�IE�K��]G��;�����KOڪPYLz�*E�&�Qm#�Dg����RO�=�k���jH��x��@<Fm}EQx��Sh����YP���2�:T(�=��L�*⛫h����;2������_��?"���yW�^��6Db�/t[�pTҩ��D�+s.J�V�/�#�^
��7X��b��Y�B�)�|	-�� pc&S����edQt�؉��K(Vu�046>�}d�5�a��TR�nh�a���Nh<Ԫ��D-�A+�c��4�0֊T�=�a����݅�ю2�mRF���v�ZD\��!�*���*� ����r]�LF2��r�-�z�	�%=����ԄR; L�'*�R2z��|�?��_��K���3g�>����w��=_��cf�ۀKo��[#�傳p#�A�X/U���@O{'�9"�~�C<��Y���?�,6'^~�Uy�������@�
ü�Ӟ�\�LHCpc:���U�M6�����$��4zNiJ!��yY�b9J�B�.��j|w)`9�Bܠ����p9�ĆM�?8�W�7�F2��U���q�рjU7�6`�ř��Ȩ�C�f����M����hX6?��j"�@'x\3�M<dH�����    IDAT���(��r`y¢�����߁��rz+��I�M���(f
���_YAfq�XHlG�ey�X\�@A����6�	e�:v��&�*Օ��i��*E�އ{?�1��[��e#��hn#3�.ioݠ_��c�#(�=n�]u��u�`����8��Q�[o_��jL6d~�ӄ�:���P.�a��j
�~�G��뢉Y]Z���^t��y�pi׮�k�D�oS;���A�P��k�Ў!m>c&�w�p�
7t%s1�5�Dw�3:�>l�oE��	N�zI��x6�l�
��)	�L�\�bcmM&2�v�ܵ�U�t���r�������I�A�ˠ(�v���#����ڂ;����6|���(�V��Ϧ��ю` (�D<�G4^kǭxN
x6S�\�8���G!�v�V-���aG:U­[�~����C=���@o>F1�.W���u
�Kkr��s������D�9l6A	ο�6�q�{p��1TJy��� +@Կa5���O��
��������6�f�:��˫�����V\�O,�8!b�/@�xkk��v���Y�Ǵ��2�/#�V}������>x�z���sE̯&pyt�\y*�س�;�Z�9a�ې˗0:2���i�����ıg��m��\���XY[����f�4�������BE��Zhu�&�KD�p�ОAX8�O��܊D�����ά�\W�d�w����ܖn�Ty��5�Y ps�W��:��j���͍���MϨ�T
J�Utt������ x��8bш&c������
nM,"�&g�D��߁�w�۩|�'��q����)�l^����س���o�զ�/���]�i�fn�/��{���[��3h�l�=��c{_�jxL��+���+�Q(�k�&�Z�Hx��*���ýw�`w�h������d������a0�
'���Q\�����8.D����h*�$J��n���$�RD��I9��䂨�v>4�W5�Q�4��k�-�����!�r���$U��f��ʟ�TD�C���.C+cø~���X�����B�SC'�i����~�L$����@~��&hs�|�����h�h�?�C����:j�Nߏ����q��6��]7R���_X�m7�=;��W��ܛobeiQ��Z� ���L"&~�;���g�.	qܿk� ����5�x��7���M"���R7�>��D{f��fh��=�F��݆���/�cy ���W2��ב+D,�s��3]�����$^���q�5,2'���9Ąە��sN�����t6t|dXC���Ei:��,tҋn��ك�����݊���C!�B__��+"��3�lzz�d\v������nw���p���dA1?C#�Q�2?$��*<��gcP3��<�E�`�J ���>�9l�8v�nt�auu7�g�M��%���CO_����sb ȥYQ�DMרb^���ڄ�[7���&���g!�K�}�w���<��^A�4G*��鐡vMg��k#b!L�F�VO�c%69id"!��p����lk�!�U����(&���I��y�vk�����~�#O��O~���O��/��OG����կ}���h��je��-W��>�诛�`��On�/ξ���~]}��?��?n��n���m�A��2�������t�6���g�qm*��)�WCf]�Vj�5��C~q�' ]^&Ŵ�$��vw��6±tJX�����H?,F!�T�7�Yj�kL��G�h�O¡e�*��p��M�͆���}�>$NJs@.&����*���_l7��Y�+!|~�jE�A���B��:u�>�w�8|XO �zv¹6�6YX@au��8��@�S���:��n�	ɗUb���A����EM�TCP���4�P��]�x;IE�7�[ÍV̈n7LQ�̚�֎PK!�-���t����jEk�%��|I���ܸ1�lA'M��u]--x�C�������N%=U�kkE�`���V\Ёc���) ��M%�l z���N ���lm��VK�d��������т�u����Q�契Ի2Fn�ԫz�z��j���ō6?E\F��M�c��u劸C1x�lb&�����WĲ��ptliiq�4�t���&�y4���+66|�,������HDc�mo��m��WO�����O�P)�r:�s{D$�B'����d�,#Z�es)�l���΁��,�0)ۅZŀ�o�7������S��7���"�,2���N��KØ[Z���R�&���b� �k|.�8#qS�|�
&f��w�n�:q:��P@�XA�j���f&�m�������C���L̀�x
k�a��q��'�eL��C"_MH�'��4'c"J&:VB��A=���8�c-^�.�0�����F�W'o��Z���mMp�������Ka������}����8<�`~yM����떄m"�,��069����MI��W*��6��s�rǑ����s+\���L�.��� %%Fkf%┽��`��^1�϶��vt��# ���bcSX]]�����>�@�`7�.ҩff'��f$a�#�.��مMIi^ZY�f
�?��{qp�)\c�f�h�<��p&�Oe���m��8xhP�@Z�2��]��I�/�w�.������C2�ǯ�='�aO�
˴ ����7�C�8��0ۈ.l�TL��1��{�g� ��T��%��ﾍ��5�9s7���h�;>�����]��VX>i��J���"�|n���T?�Q03�$��T:/��D+�F���h���Ҽ	������4R)�!bs�ns��E�4���u=vlF�]���_z�dT��:k.C��kv�U�sV���:��� ! b,�7i�����MJU�-y�]�4#O[���u9<t�	��>�];���G���e��Gi�g�Z3!�͋1�s3��uo���ZB6G)��բCoW;:�mعcN�y�hPx�D97����i���9�L�;��[��S �S*uX-HgR���h6��ѽ���S���ŔL���ᔴZ�x�6l��8�*ƗWP&Bbv�i�����*f����E<� �"Ɋ�B�WT2I���v�㎄v�x��ڱg�v������&�"!����t�ac<K�P�!S�BQ��V%"��N'���uww�����(}�����Jľ�g�\'J�%�ƣр%�8NS��t{]r/,�����h�؍2�&�������>z?���x��7�(�I�\�l��/Ur��FgO;���Ǳk�.<��g��Kg��ʬ+��}�_z�Ӹ�̽�t�m9s�XgP �uD��͙%�t�"F'g��B6_}�b��P�����#���%��R.-hu��,�E�ƅ�x��(��%ԍV$��r9��O~����׮}�����?�Y4l�}�տݹ���/=���+肓3���h%�Å�bE��¨�KM g�%`dl����`8���	�{m%���lV������B�h�dQ�����kӸt+�xՅ:S]Yx����YQM�a���,��of ��e0��<5&�W���-ǹF�1R��i �i�/LU�
SSih���0R��Hl�M��Gm�:�"E>����0X%��f-w�����?V4�	7f1�"�G󿭪	��)[U�����N�l:�r�ފĂ�Όz�&���`�a=�GQB2�bY�����++��B@�nK�!h������dr@�$e���p��!BҌMׂB�6TS0��/K`Uˮ!����ѾoB�-$�����)���̆[��׷a���&+��u��t�t&��ce%$eKK�m^�)��������&����N�͑��l��Y�@�����ꕪ��܁��vi�����7BX]�@._���W���4�~3�M6�#tu��U��L�s���)?��<��±�f
�hm���n�w���$}�zz3Ց(�M�Q�[�h��Lh�nq�ڰ�D��s����y�ZXQ9��k� S�X��13=���1����u`���fifˊk]7D���H8���(,V7bȗj���HhSW�ݢ=��m�欫�`����W�N��@{G'�>�@�V���v��<������bc+_SP���� �ž�;l�K��+8�9w�
�~/N=��}]��E0M4��9��X݌HQ�9p�����@�0���`umC6Tt�`�,��������L��&WW�Y��E�ri�����R�;�FXĲ��zo�7�H"�r-�C��;;��x��Z2�����6¢������1�bfa3��hn	����>�L�B�!98���-�������mª���݇�o� �KвA�+c�����-	ו�H���mi�G�+��2s`A�/���tw5a������Tč����H��d�����n�ua���������{�a{�vx�N��9������-I��7y�G~�mB��|jn	�ˈ$r0�=��ZLla{o3��؁m�ڑ�%����=^D"5�;wW�M!Ь�W��:�2�?u��P-�g\��7&q���SEq5a͌���w����=�r��e�OL�������,x�~�#���f�y>aS����x�Q,ą�`*��ӏ#G����q<Ҹ��.`dt
	R-.��5&����CljZ�H4@��:e��a��A�)bdAKr�r�a�{f}6]�A�ˣ���˿@)�]�,L���m^�����1��f��A��2Ӽ�~͢�הg�8ꅜ��R�&�6[���Z��:��=�Y�w��^���_�|��9�h��!=tc�PI��)�%Z�W%e�`>��tF]��Z�q����ȇZ˴8�y�&~��K����N�#�! �Q�
�v��QCa2��*���g�����H'CJ��z�e�3������x/��:�.�����S�a4���|�*6�4I����P���/
��/��l���Q��J�:J-�Pl�i�]D��\o�$������nh>Q��n� 	⠅��wH��1mH��d���Uz4���ag��	⠆��|N-��b��
�XGF �c���u���:���ƽm���k��Ɩ�lv����5N�s���xᥗ���.<6�l�x6�2I ���A<��7��_9�<�,����^�sF�7�/~�?��[[@?;Je�VK��_�	���X�%�+���R��S���<�}{�bL�0Q��o��:��������� l��J�T����7�Ǐ��4��3G��k�m
�?q�q�y�0��v�D�G�Ɣ8������:=`��g��ML����tvt�;�����p �6W7QȤ���ms(��<T�&�`mr��W.����������%�X�1��?����K�<�p	NZ���EE��/���	�G�&�䬑ʠ�?*X��u���dit9\X���H�@B�)�J$�܇HM����t������:�tg�j�>�Ǆ'Z�x����J4�"�bi�6�a�يp�?K3^#����п՚�aϱ��s��U�!��ą|���f��gf��a�;��-��(�C�����'�,7\q# mIkJ��uecC�
��4~`MMw�FT�u��߅ӿ�t؉X.�͍y_��*�!rT\T����dqjbl�N��H'���\\v�v��+�b���[�[䄑ְ�
s�X)_�h���&'��L9�`� �<9u�Gx+&N�bA��V���f��y-�0��H�łJ���Y��5d`s����*6�t+��2�1#�Dt�e�%�3q*�g9����>���Ď�\FFM=*W�#Y,H����	H&�*V%_���F�'ŝ�붣��S�{\^��4�~�o�^���'��x�*�B>Lx�twv`�A����i	A�j���E�1�/m�6#�(0L6�G6�B�6�u�w6c�@�fz��&��P��6B���ƶ�}r�(J1B���P\Rhg�ezMz���B�B���EO'~Z	��o�ٳ���78��N�ޡq?�e��N��"�FzZ~���Tsj���O���	fE��B3C�迯֧�f��W�II���Ct$+��+��I@_.b���ػMNZ6A��/���/�aqu���#��.7�i�)kޤ7!��ʡDH���KtیD�1�ɢ��Et!�&���+K��1���9�*z�Z��/Ҩ�3h�Zp����lU:��b�rs�!��`�;Q�V%���R�li�LkC��K��rB��8Mع��?<v����8nݜ:'s=}=0����hn�Cx��W��'p׉ؿc� [�Lͬ��ĸdT03���hmn[�T*���ez��Ed�ԗP��ఖp��p��>�3���;�s�Q���B[y��^�2�������#bhҵ��11���pL�CX𲁸��aѼ�	_�X]b��(^�=��u�!|術h
8a��Q�����a0�����&/��ײ��W�r9�
�y�1BC��i�"GPEZ�jnO,�X\�{АB*U-��x��̩@%nUb���'|-'�Be W!�͈N���Y����(��2�c��bM�@.:�4��60�fB~��������C�Q��_�����4A��_�(瑊�@_L����/}�RP?���ɟ<�����1����+% i����f�������u��$$8��Oc��G��{�Q�U� D�Q\|�2^{�_��۶���5�/c)Zq�s��!��kǼ�t^Y�{�.�|�ە�o��C{{+>�ȯ�#g���駟���?`fi3Q|\�.�}���W�l?{�E��/#�B&G-]d6��L��ȵ����Yϐ�]ʉSy�ܻ�oԜ�E����es�$P��/�N�E�ً�ih�4lj�*�%���z�X���h���-��'���H4I)��z�<�'5;���e���Z�Hg2�����燍t�"]֚���"M��Eٓ��?���(�|��x��W����t��B�D2E�,��?���G�����M|�c���k������`bbB8����|�_|��n����I`!ia�LJ�ڐ���Ǫ��j?~�g�r�*�2�N:�'~����	���X6��!�"�sPLOX�n��7.㩟���\IgF����~�
!`0��:��d�����6?�tK�cL�.�Gl(+���;���/\2
�c�����g��ѣ'��/M��8�\V|����bG�7��ׁq%�����"^�0����!���aA	�.3L�(��}	��q��i�A�i:m�
�K+�=W�f�&BU�詅$�N�IC`�0Q�N`T����	dՠ )�&���]%�b�5���U�<1�R�sc��NQ4Ž��t͎M�A� aU8J!@����r#`�b�<E� B�K'e���R��L���c`��:v,� b�:B�,A��'#qD����
��I`��*qA{�>�;(�_xq�P�_��D�WS���!��sEq��>�W��=C�h���*�!���9��r`aɄR��gC�h��v�����M�DƧ&��Rf�N�W�SE��_�@�a	ƣ3�#v�LC�������fz(��t`�S�)���N%�ҙ`�{Ul{5�C�={��kw;��*������2tu�=�A��hj��
XwZ�2Q�%���:�|�\�]~���T"��&�
�f�T����MeU�B��+Z�Z��R)L�,Hx�p��a6Q>�K
�րO,Ը��TTJ%����e��fKrh��+�]r�s��e#0�ӆ��&	��3\�ױ����b�$��Z�sW-N�@h-����2�|���9x�Za4��`RɄX߽s�:}"��Z��!�������N޹�]W��;�t@$����-�#Z� �.���&g������lQ������հ�����&��'yM8��J	�]�8�s ��8�� �T���-�{�&±�tKk���}�K�,���BO��D8��""������Lv;�D(��Q1    IDAT�%�p�S3��p	��1���nx��l��WQ�F�� ��ߋ�N��gRx�Q���(W����-��V:c(K�!��2�*&-������GoO����rzӉ�dP���Ĕ�o�l3��~}Dh��}}8�w/�Z�	����-�gX|q�5xȫ��1���-�hC���t�R�>����}�@�����>llf��ۣ��	�^s��H�e�G{�	��:�ަf�r�3��H�F�(�kiF��/��< Z�`}��.\E$�t�:z�x���1��+M�P2�qLO- N �ʔu�`?v�DS��-:� ��	���a,�D`4 e�Z2��7������~QƢCa�jb/z/��XM��XB&��c�S��V�^�sSx��O�^λ��BGj��(d��I3u���V�2-V�t���5��p��v�w��i )�F�V��b��U��9|��	|㫏�}�"��9T(�����M�ݥ
W>��&�Z�h���H��f��/�^%^c��{��ѷǏ��hP��jvf�?�~�����!����H�e@ų��X��kHg�H�Ҁ���x$YN�������'���<�),NM���ۿ�3�=/Ti��!((�ѱ� ~����о=�55+��#��29�R"�(����F��j��`R�C
�9�$O^�3qo�z�0A�v�Z[��t�����52�����RQ;Y�+��ަ=��QQ�DXÜ�rQ9D�.�<y�F5T�VV�����A+��x����#h
���pK����D6S���Pf��_��8~��x��g��K/au5�l��r��g�q31Գ[8vl~����#�/�q����I�tu��_������n�cy5��naf~Qj("��l.��؇p��	�,��R���E\�x	��v����<��wb�Bɼ�u�O�B"�%��K[g��q�w�zpa"�����+._�Z��rc������ׯ\�ڼҿ�Y(C��|�G/|o=�=h��D���1�PىQ�C(�`*���v;�n��y���F�n}��Ò�ZL�@��]�aW*�'F�~���l�a%��i���8
F?�t�*��&ԓ���22��W�W���h�*=h�0��q�7����S��\��!`�(���E����ȴ�! ��\���)'!� �8�Ҍ��T@�����ZxM�Ŗ�1-��7i	��A�q����s��f�����yHK�49��Y	ɒ���6�>��'�=ІD���L�lQ����b��/,�f)ǒ�{��+�Aq5P��[�#�5��� <Su,��I��*K��?��|�h�Տ�XX��8޶ٓ8ru�a+�`*҂��P(��:���T�!X'߷Z���Ƈ���[��*tU�PU�b#j��E(d61.��5�y5�)��0�M �.�cE���Wk
�b(��TEg�@��#��v9����˂&��ѓ���h=�JbQ�0���f�)czN�.M6�ן���{/mO3E%8���2�g>=�Mf�p�"v����d�)�şѠ�sڳ�q�vv�J��il��D� �t��V��t��0O�h����,(��ً� ~�"����"�
ŲXwwx4��L�K�[3X\Y�����,�F*.Eq�|^�Z��Q ��G1��.��^��dFoK@�C����V�Ji��<,��U�"I�O� ��B,�C,���d��*�ޒ�N� jOQSJ6�s_����F_��u��y�g��]nй�,��M���a��K�u�zc�=Ai��D��r�T�U���iE:15�D&�@��w�BWO��\�F\�x��7��@ǌ��"��lD�@dT,Z��ߍή&�٧B�6:��HR�X:���IB=ӂ�De�p�Չd�r�s��z�]�-��j��N[BR�r���i��&S�B��_��jq�a���mC��	�` n��Y�0x�n��XVqk|k�0
4	7�D#��a���bh�;��Hj9�x����y���0�9���,R���8qtz[�ddݳ���Q�L>qEj��([Y�q�ŀ��0.�{�+[0�Z��3�8z|����0)�fM�
H�2�PJ_y�O{<6INgA\d:y�t�&�|�]ds5��Ai��[N�3(�P��)�69s��{N�=s����N�_�l�	:T�[�/e�}���P����fA�ˌ��-��ܳ@,
��&E3�5��D�Z6��
/Iy�)�Q��ĽN
X���J��#q�1�D�\M=��
�0���h���Oa϶^i2I�I����ٗ��K�`#A�n@2��E�C��':�g�BQ�
"�$k�	Idg���G����q��y.i�I�Nb���~�Y|��G2�Aw� �'���Ь�+O:�t`d�%dIueHu(�3�\g*������~��/byf���{�h����G8����:��v<�_ÑSw#��`an#�cjt��-���1����,z"�L�V�I�
��6���et���D�q�����6�I��|?�_���3K��F���$ϝ��C
5m ���|ѭG���%�jq8U�k����>�|��_��I��l#���XW�|����������e`H}uo.��o����S�>4(���U� e}@��%�-��~����=t/�����_�)��c�у���~>p?���{�^y�"6�	�5,��"�u����ß�N�{
ӳ�x��Wq��w�݊���{�����u��fp��E�{�=�ܼ%N��;y�Їpσ���.,�������λ��ri��~��������q��~��޿��O����q[P7�$�������R�P �"��V�U�4v�\<�;::��x#��V�z�k�|
w�/>�
a�*��B�\G�`@8<��i����5j&��dn+Z��6�0y�U�Cs��"6&7�����}$w���#vu�SԐ ����@6(�վ|J�wr*���	���A	(�R/b�������,�AA8O	��e��>ŉC�����4�{l"$>[�eqſ������Uʤ[ُZ�vI��A��J
��g�a�8�a��K���$r�,6W�XZ�W�T�,:���)-�Л��'͈j䋮&R˾�_�_������7,j�<�ُ�>�q����ŭЦР��6e�*������M�?��� 	l��!W\���|fe��G���3��%	Q�A��Y*ݚȏN\^X��� E��K+.G�E��9�#�|6l�]�]kN��'�MM-�ZhYA�oE�E���:�yoMu �ΠZ��	f��,^�0[l
�����!��i��,`�(����CR���}>�V�Sb^�|Q=?V
���$�۲LԼ�ޭ�{=&:@���Y3"gT�nT(�6�dRE/f��$�%��(��x2#6��r�jE����f�9q/�oBo��M�%�uf�æ��i�4��[=�^Ah�'��q�^���:<Ru�hx�+��'���M�wW6��Ax+�b�"Sy�[��L5��1i��E��3�6I�S�ӈ�
D;�4V����j�Ey~O-EDdJ�3,V:���B�h*y�>��=�r�^�B�����1;��HtK�(F�wv�%؎`['�VW11zS+��雭3;�	5A{u��.��߱�f���cq9�X2�<�w�,��r��^�{�X����B�h�#�c��y��5�]�u���#�$��
��(�8�i��ffV�������&�E:�	�׆�}ؽg �"]G2�6I���R
�n����ˋB�C�4���Ut-ط�W�W&��Lbf�ϕ��.�!$����V+vlkCok��5
���`y $+^J&r���\��lyq��Ǳ������.V��B-A�:��79�`��>b�&x�~��PP%�L�TB��e���WFp����&�����\0[����	�}堅o$�W��R��Ybݍ�u�A��yf����{���1�E��J��f�&�f������$�Ne)٠�ؼZC0؂�;�K����4�Q,0y�H�Ii�$I��J����g#��qF�Ѵ�Bd��Tǝ�w�؁]��Ȧ2�px|r�s��q��A��>�V	�4��<��t0T�8��b1�=���}�Q[[ՐΨ$��xB���z�T��V�=>��A��ģ�	�+�$����B��"<���E��r���7���?�YTsy������߅�탻��X�h��#_�5��013���0'0=:���Q-I�%���Ј��Os�s�Ć���Fs���6�W�̩�Ƽ��%:.j�h��g�_G?��.f4���X'F��:)DH�gP=���f]�F��"��r)�Ώ>�|��ay��f�}Ӫ�t��w/_�w��?���|^?Lz��i�Q<��/��p��qi�~��p�֤��Ya�%-��l�LǏ�Ʒ~�wp��3x�+�����q���9��{_ǃ>(z��^|��s%�$��m��ݔZ�n���ѝw�%�����o�@6���>�1���~V�����?����E�H��*�g��Ϡkh;;�m{��f0�=
˧&�Lf�G>����_R�?��!��#���w�ݫSw9Z�0ڭ(WrR��HW�&���TJ������+Y)�yx0	�����I���=;��O'��G)���@9������.��2<���8wu�L
p1��iF6�(.C��"PKJ(h�E�5D��*-�M%�dQ�H1�&xh���o}%��L^��7_O'�w6��Ft����3`�"��WSŁ���2�{N.X�K�]]���{Ni(��MQR��2I����$\4�^P��r���*b@�L89Q"[.�a�{�=��<��قx�(".�3�$"��������.i��zA	��, ��AqaR�FC�>�
E�^<�T��3<T�pU=X��}8�鏠cϐ�.R�/]Y���>�"��a;�I����z���X�eI'0� ���L&�]"�P!�Ȏ:.u:�"�ͩ���oA�H�G�$>�174���%#`�YTE0����mK_S�6'�,�gM�&베�?�to��q=R�O"i����>�B�8�d}�O8�.r���1�Grڙ�i��W2����U\Y��U�C��(p7�ܨDcC��N#2Y� ��H;p��ؐf8�7��.�Ox$*�C���g���rr�C�Š���A���]�r¦�h���,�;�SRق4�3 �A��#)�D��*��R�u(��4�rU�!&N����t�X��'e��"WB
b�V@PB�`Ӓ�q����Č�i���(kr��FHgd��	zY�aC`"���Ǫ�l"x�X�kQd
�Qۡ3T����^/�����/�&�,$��o�m��]D��B�8�7	����!��!�ɳN��*L�Y���^"��$,�"�.T�5[ܘ�ץ����(6�����4Z8`U�V���c=�[��q�`2Vhr��w"���!u	l
7CId2��l��dfF&��z-���6��4��8�^�3\�6�d.#6�,l���i'�ǜ��y�l�^u�$uc3�յ4�
�[Q,0���X��:��	�-y�o�\�Ju$h���
�`fr�Qح��DC5G</�l6:�x���G_7Z��&o��
9e�ۘR��Fˡ-	mF�&Q%"o�Z��pC+����缑�9��U�C�sC �JKH�kĉ�m���2e�Nb6]m.�N�4��;s�&�Y���Ӿo���l_�]uY�-w���8W��1��IH���$�痄�pr 	� �``���^$[V��UV���w��7���o$��w�9��˗�-��~�y��ۿ� ��",�R�=��CI�RťW^�{�y'�o܀'�|�}��r�"��$�a��j�D�V��Nt�h��x((��穧���U-���a�s#�,�#�AZ��"jk��6Y5�݌r|w�6�|.NH�� Kd��LfE���o��ׯ��2�Wݝ������c'u~�]���ʎc�:+�ƕ�nD�-A$;S�Ht�3�)�����q9�<�w�{ߥ��]/���|��q��Qл����Տoy+�t�m�]X�d��2�siL�C9�-��ȼ�F�a�g��Φ
��Zرc;�m߂ٹI����j�i�g��#��%/�SUS�g���nQ��6@C#���#���csF�O��@�%\���V������lހz��1����I�\�[|&�>����?�^8ѐ�H,aaa����˿�4�]����#���?���������'��Jn
�،�����oy��?��O����ؾ}+>��_�w܂c�f���>���Eݎ��c%_D��S?������������`f�4|��q���� b?^�s������cs�6m��`������#Չp<+�p��f�����{n��g!�;���o=����o/�,X	�Q;�S�D -x��~'{���v�P�\y\K�ZnY~���f�ܱNz�Z� T�A+`#O��_��^>�E3< _l:��ަ
��(��8�za'��/$��a�Ž�D\/��VTz������`#��	`1���CI��(d���7�?w�

c���3Ԁ��Gw+Âa ��"�n]ʍ>S�ؠ�8S�g�r["��,Yl7����^䊶�=w��m���:� /���@V,�T���N�����z�!�R�]9���Դ(C��)�j��QD�F�@#V� ��O|��!j�F]�.���D����������{�6\��7a���X.�^Zԟ�͗����Ռe�h0��M����69r"��CC�����@�����hW)�����<����C��V�?�A�$RGE�37��L��tq�k�6+f[��~��C	�:=�ikZj���h0[=6�>�Q����hM8(��Kژ_�7����)��R�,�.U{*#���Y��Ay�Xx���,�Yf6��9�n8�Z��g]�4�b�i*@�����D/�3o��5��@�`A�2B�PJ�٠����C1`�&����O��bW��5�5P��͜o�Z�Lضy�Լ��!�o�{�:lft(�χE���hX��fiB���z|Q�Z)r��TQ%�ؤۇPb�R4�u�e�h֋Z��Qi��s���D���h��
<�Һ��{s�g�am�+Z w���
�a�7�h
���jF"j��K��B����T�'ت���`2��/%����A�9,M��� �}�HZz�,i5�w�p��&=�r	���P�v0�N���
��9�ZPL#�c��%�k+K��ٙe�Ѱ�.ʤ��DAp.M�Z6|�z	���������T��ߝ��N�aBi�+���YA4��:���PS%݊����J=���o]�l�$Â�؀�/��6�[=Kjn�iY^��2�����WVLNN+�Ո&�X��E�]f�p�$����
�j�8�
)����(��f3n�<��0�פ���(O�%*��dL�}������@PZY�Eu�����U.�k���|��y�V<��K��/|'O����&6�j�܁��aG#��eD��E~N��Ʊ��K��z6�Ә9?j���ֻ�s��t��)"�B��YN�%�O��Ԫ���a."���'Rf�Oa�S���M�OcrrR�i(Q���P.M�fqI�P`�+$���K���^�vѺ�[ai+�f�Pv
�����E\y��(
x��O�[?���et�^���ĺ�硣 ���̯�_�cf|5n�_DH5s�jN�'��̥IA���p�mo����������ߓ-4�wHEL&��H�+/�Q���12I���Ya�MD��"Ƭ�<T���ڪ�/K�H��u���/|��x��G�
�X.��ze'�V�ϩ�����ǃ�x�N��>���Ht�Q�7�~�4�l�7��]|经`zv�2s,��~��"J�)\�c>����w�O�x��G��_Ņ���G~����[���k��?~�GP�P�EQ�5�[�ܴ�?؃    IDAT�¢������\��������.|���C���?�2>���\��*�ƪ�u��l�Y�����!����6��̾w����ȵ�>��'�K��9v����9�y����7�>��|�2���ux@D"���j!�������7�;�߂Z.��-�!�j<���-�/?��s-�b��l8Պ�+]� �A$�M���-�r������&���]����Ã��M1�fڕ �㑘�����^�,A�|i**@����h;<�OW����F$;�$Ŀ���� �J�rQ�RKx�
�$��jf�D�~/�6d̢'�FOf�F�F�H�Q�R�B^/2����7<~,��r����$5��D����,&�Cyn�8�D���lhm^�	n3�i�9������m7-SM2i*�g��=������ʛ����M�V�Ȯ,�����HF��j)�nR�;�u����7h��6�-�]�����?Bj������OG*�zdE�&T�P�l5Wr���,5ޖl/��S��tP30 *@տ�Q%sr[C�9aT&Z�	��{�}�3St�	�ͼ�A2u5_�,y�������ὨU
J�֟%_���p5p�58��
?�&�̈́�������9��<�]uǸ��j��iX�6�����9�Z<0�Ǝ���61���2�7�7��:��A��f�V)�J���/�w��&�t��FL�2�B.����Y4�#	�9ģA5�eMDY@:Tͪ�pR�8��oy�%��2T�J� �kR��U�d���FjŇf i됌N�-*&ݎ?'[d"R�yZ������K�W/jlm�4R=	���+GMן�)z՗K��D�u��C�0?��^�&�����K%c#IosO �~4&����"+�j���I�(�ѩ�� "���U�+@�;�79��Z����0��PY��I�Jut`aiY֤P�H>�-�of.}$_�B7�,�in|� Ʀ���~��`v1)"9ʁ!�Z2��#���F�l�s�����iA[�@V����D'��� b�!���S4�����^i^������:���ޕ`�)�D{��kŌR�6�[��.�HM��p�GGG��m�\?�
�i�h�3��'��ҹ��!��=�Y�\s�Қ���i����p��p�s���gn���Q�I�i�>;tZ��#x�9�"�o�IW���@@ǯM�6�o�}�x�������͛���W~�� �\���"`	٪ɦ��gw��j�Z��Q�@�x�ב��@~y�����2�q�,�lй -S(���`���9� �p����-9������u(��������9Q�]Z'� -q|�9�ynK�@@�c��1���SD���E;�����^y��8�ry<��nL/g��X�����
�;��#g�]�ayf˳�(+��5��@��˯FӤH�5oX���މn��h�|��x��Ȏ��0ؖ���-����<�^�g����Δ����E���]:/tI�=.+z{�e�*������jUsN|����o�	:�q�O#�!�4���8�����?��#��hI���˽�)U�}�7n�����b���x������>f�P.q "�k ��WP�O���Ç?�x˭7��G���
���5���`�ރ�ߟ�J^,�}p�a�h�"3R�BY�B����Ό�vJ��]w�>���~���~���OK��G���y�#�K�#-���*ٽ���}��8xv��/��e�S���ӿ�����ɮ7{:R ���³�*B�e�����D�AH>��X��/���j�,��&��}w܂+�ߊf1?�l�hoǭH(�b���<���W0��b� _��Y��>��~���舲�sW���1��Q�,
l>XM�e��>1���R�ϰ�%��%=)��:mA]ᨉ ��酅��V:4�m0��C>�f{��^bB��5M2����8��T�qs�-�æ�֋��FtC֜��%�j F�PE���m��6�G�g��4�VMf}�|�B����ۏ�҂I�j9J��zk��Y�wؼ��D�ܠsf�;�4�ܴL>+�Ʉ6QCд�ܶ���:����ZI�$�)�Y��60�)�Q(���`T;���Wu��������G�� t�`Z%�<JW���l2���L�	�&�N@t&�AA�{�5x)�m�q��ѬU
���Ó(/� J�6؈����nW�M%���pN��y>)���(�2|�G =�2�s�.u��E���4�d�D)�dR���f������-n��F��t�
��/nQ��ƶJG!
��s��v#�� ��8{ˇr���6���?�6�Q�)*f<����1�RC�Y��J�!�G���6�<��昴lY�#����a$�ğ�&�G�!���Dzl��!�M0C&D�|u�||r�hh2���N�mӔ�TqK$G�6�\��׽f|�9PH���F���*����,�3:SQT��0�%d�M��IX����8�g�ͽqә�1t%L���=#-(�H�"I�%��DQ-��8M�?u!~ګj�!r�B�t�2�RB�d�ƻ��e�T,}~ۼ�u�8�R�c(gy��h�Z�]5�Y�#/j�Ic�P�)Jd��������7�U
�� �~��2�z�j�Ac�h�D�F>��J��VN����o�����/�֘�QU͓^�N�s~�]�.��c���jrP�� L�%g�4R��1�&*�jLc%݅���r6��@�:)Z��Ս�-FUc����G. �Vr�#�.包5���B�F����.����T�F�X��le"-��� ���:,`��a<���b�PH5���6��R^=����Z쭤���s��|����w�i�c��jlY���FXMf
|_��2"ޚB����4lߺ7!�YJÚ�a�u���;��; z�	qcݥ����BKf���f{yæ���ަ)�}gM�3Q#b(�̠�BJ�N�X@��{4*��϶Pp�XX��%��w�}���:�t��� ���cf9�t�.���r��&pjdss�H/d�O�!���<wGW'��D#�\���T��Ƚ�o�Ϋ����jى~�{��'�W>�t��aˏx<*��-(�FL,��[>/�Ѹ�a^S��D4�H<���3J	����M��$(�g"e��E�����{q�[o��5�ܐ�*�zz���gy�*x�'��?���t�Md'�X0*�����m܀����b`�*|���#?x+�<�%.$�{B�(*^F�4�+/;��ɏ���Ɠ�����������Ν���e\y��xn����	5�
*�`�P�YĺD��ɜ֖��&i6��߁�����x�����Ñ�y8M?�%G?�L�4x^r���	s�h�J�Vzf߽������怳��e ��}������<�o�o����P�mį|qՌ����.��/k��pIh�A����K��ý�܄k.ڦ�r*�e��1SbkMT��|��#84�E=����%$-�ZF�I{ <myEQ"��M[��\��BJ�r���E�A�mg�e8�-�F����~�N��4���	`!��M!���X��OD2�|n�R��-�K;��4����i��a�4Dq~��@��t.4�C�� �bLbW6ʌ����͇��ؐ:�@ej�\w$�a
���� ������C�����FDcnRi�l"�m�� /"C��]/y�/-*��V$z��7�cP$5w��Cv����[�2Եi-������m���W�#�%<��8k��4�E�Y@�y�&��D���}�f�����с�M�(o���0`�GII��2����/a��h��6_����E�
�3q���Dl$ƴ�`3xE�����jñ2�
¡����\�����s�g��/�r��w�g܍�l��ś>�L妵^-�Q�[.���d�5j�p�fЖ�����'�^���D��D�q�#��Y�}�EU�������j�Ԕ��7}z����cM]:� �Ґ�]ұ���M���������2r�� �_RY�G� �0)�D��8��b[�]5�VÂq&E�U���� n
e��ƛ��*�"���O�,BFkb���50+	��}j5��wL�B�e���O���7Ä��P�`1�G�
-r���L@	%TK�T���hu)��=#���Mɪ%����"=�iBP1�U���.�բ�il.:G���E�8���"e��9J�o�	�E9��z� :9Z�6�~r�)�� j{�/����Y�Y�09Lb9Yb?U�O�5ekɤ]��J��\�2����N�FAz-_�,��&:�
�����ZS2Z�5}O6�^ݢ�pT3(���:);<t,�0� >�Ǚ L���0�<j�jՊ���`(�H��_��6�%>i?�»�M�~Y��^�nO<~.&F�B�y�hv�1�d��m�U�]a�X�^c`C����ĥ�D��$,&������C5�F8е�uh�Q�~�py��B�I*Wv$�A�c[�J��Zm1�������OV�>w�݂�Q��aZp�RV�%�o��[Dve���,��{�ƚj~NC�j2T�}~�@�"�ڌ���A�BX�u6�w�j��C��2�kg���1��o�SNXv:@]4��ͥ�Y\{�e�붷�K.Eo� j��Ɖ�S�_�tΑ�r6W���2&�g$j����%N(w��Z�hB�H-siW���ǭ�݁ށ~o�M$cx���c?��,Ź�d�O�6�|��٬���4 �����}}}:G�]izD�;u�$fffdMg4"q��m�sV��7N�:�^���|#��ηa��u��Q	����O�Ңv��x��w���x�Ԉ44<�B�޵J�t�e}����OcÆx�����o>�م�B�P����5�[�B��᪝;�@p�U
����;��/�����k��Sϼ���×�o�1���P�逇C��l(M��	oÁ��Cqz
�f�r�����z?��&��{����82�,jhY�[.�嚋1�<=~�|�s�
���{�]�㫿��#?3��~�;���G?�T�m����j�RP�m�e��U��-k��bq�YL�`�A�@P��rp������7`�-h�����6�<��&0�m��?z/�A3؋���Z�ÄU��
q�fD|�yz�k����3�%CC+�~؄�gh����i'G����ni�ς�B�M(�Tf'03���k:I�eG�B(�M4�9&�S7�<�,�W6��@��B{R��M��-���V��S�i"�����)g!�A��1#��Km�4�fkğ���6���&e�NDvA��j����I�=�����N̂�V5�N�̽�/"R꿙&���6畍���t
����q�]��c� ri�K���e5.?&q�g�U9��g�-�(ݢ>�q�����/b���-_(W�Y�Àd�8�	�!���h$���k��w�i���T�<Z!��M��t���-�(Έ�9����CK�#�`�l���Q,�]s��J��͘�`�&���������,��%��-�	l�،r�d1��L	��@��Hػ�M�a�����(ɘ۠8�r�;Ք3p�T����BÁ�0�6���pT�!b�!� ��e&12����y8T�0iZt"e�Pn ���C]
t�j��<:�Pv2
� ��ߢ�ֈ��F�X�D�h��=�������X�5Ի*GhQ���4Dl�j�.���C���#�rCm�����3��
�"-Kt\�-�}Q�x._��<��5Ю]V�u��D���p�OQ�����e��P.ԋ[~�Z�~~n��P���t/>��A�:Ҍ���+Q9 �C��e+��>���{Y�kV�#�e�f��Ơ����U�+�C��;�>j$�`���"�D��Z]BL�ظ���AO�O˧����(�p U"rr�e�f���W�F�M:�ʭ:�#~m��`��f
4 J����?��Q��55k�45�&�rAx<uR|Ҁ�}5����Hq9�:��zC���:�BЌ����l��=.����k��eRp�DʀY��9�^��H����	��#*��[�Zfx��0����ni8faq�`t&�\�_=��z蘁 ¡���hP�d�G���sOʊ:	��s����-2jR�ye��d��J$4��+G��{6P��h!�%-c[�T
�䳨2JՎ�\+ �]@��Aw7֬Y����lX�w>��$�P��,l� t.��6�tv	�6����YR���~�w����Z� ��|FAD��6�A��p��-x��������r0x><|Ͻ�'��`��D�Ğ��|���RA)�o/ay���u���VQ�=6-�cA�^�+w�$Y���شa/�z�<�(B4X��j��V��"U�b�f�D�Y:4���r@�(Ut��H�3�������I�\V���Eijj���{ϻp��;���%D��ċ���{.�l�>s?����].�����������̧�oz�8v���_�SϿ�R��b�_+ m[>����8������ÖM�x������F�'���я�]q9�۽����Tn"[k�iZ�X	����0/�,P�
W)�W-��4�`���{'���7��#O����(��X)�3��홅�q�F';�A�P�|n��,-���{o���|������o��7���|���D�M����oӈ��_f��IA�om����1Y�ZD�U��7�o��m݈f!��y6�I�h��򂡧ˎ���~<�w�� |�N����-
%-����;̦҆����[>��_�L5Ww P�:�F�NN�o�P&��.2���q���.'�&�X�E���\mDCQ}/B�,��S�E]l���T��X.����$�L�ж��>,:Ylk乚	�nֶ'��6H��IS���Dű��%7k�>�!#������;5����&y�Z!�����5��G^�g��@��B)�m1�,Z�h��4�����;oEt��ˋpʴ�d!w��\�d��������S�\q*x�Q�{�}(U�5j�g\Y)aa1�f�R�'n�I7����>���[JD�G8L{�rYK+yC�� j���203}����.�� �E����%,,eP�q�ِ��[.#?=�_�9����"���������V�Nߠ���3�eɿg2uM�Rt�6�8�X��+�'���'%(}aa	�|	�B�b�\A�|n�
p�%B����ۍ�N��ְ�N�{�g4���>і���p�@�vlb�ό���y,���v�.�%�?@
�^��7�@�A�
*	���Cޠ-�B&+���r�=�j8eb��j���ry];�ъvh�+!��[/������p�Mݦ5��m�[�е�L�m_�\TN�Xmږ��,�D!jB,dO� kۚ�H4 ��=�_�(fs�ؖ�RY�)�P�旃�Ϙ�CG"rQIǐ��I�B.��,��C��?3+������3��q�i���|YK�Vԥb
�(5ԇ��!<҈��� ��aN&�]��H� IHȡ�KA�P!�Z���	�}��WZ��!�M�(c?*�*JԼ��6��2��K 9��U3�i�����49��iRg6�<_�t�i&�^R68fK+�����:æ�K%:�q����uBD̟��1�"6u�K�N�6F�//��P/D4Q�*�C���j�Ԁ��'� ����@�f��?g_�@�o�Wa��u��1p-BWď�SG����0:�s�g�J-�(�e3�e�h�^�C!��v4�`<�2�txF+�� JZ"��RK>٧��7GzGN�C�A�2����R~����Im�
�2��-�4h"�Ƕ�Zϔ��@T� f�5蜡��A�I�	�!���}874U����s�e�]K����	������{��N$�](ׁ�{^�W��6�B���8����Ơ���9\���&U]a��뇰z�Q�:�f�n�:�ؾ��R��    IDAT�O=��DXZ�r1�r!+����Un���'E�=P��ש�҂fa���8 R�H����0����,M7m^�o��0��X�zz{�$��".����!�aai�_~	�Sҗ,�s�aE#t��C����	�s��ճ=���k=��GN`a>�/n����x�ݷ���CCC���{?����?ę�q\��J|��~W\u�{�����#fV�(4�f ������p�%��o{eO��|��hd�x�]���>� =�_�֏�\
�P%jO��J�"Hi�;��,��"M7W��w�w�-��3����|ᖯ|��ϕ}�5v� �,���A��6B@�(�y>��<��Ig�� %����c���͸��mRg�5َ�AَV=X,��#{�̾Q����l�`�!Z*u���P�0�V�g�6|^�f��9Y���)BԻ���,ѫ^"M�|,�,�����Nӎ�'i
A���Uٜ1����P���k)tS���QY��ӛP6!0�l��\��\�1��AY��)6� �� ��F�/&�K�R�)�B;̀�CE�qE��^�M
6��J�%ߘ7v)(����/a��)̝>���	%c�����n��g�鹁@��V��@ ~�ִ�QI�;!��7�}�k�1�8�M�,E]t��1��3ĨPT��M6Y�*��tD��G2F(l	=bS���	`y��ӣ3�d!"�0|�:��X��)n�yH0y����<���dJ��[<I=
�5�,�R?�{��ۋ�nF��G0�U����
&g�w�+���M�6�!8k���I6�-#(�@��Md9/>.��"�t�I��G&159�期?[�"c�@��ukz�Q{��_(4P,;J��gZXZRW����lQ�;:��NX>5[6?|�l&y{��'�(���c۶��������!��`�c8~jT�.��b�Sw!����6��� ��*��
Oc��IubU_��z��5,�������	�"�a5��I0K�'�x|H&btm��I�Drx͹��a��,�.�X������*"��i�I�!o[� sJ��i��n; �nZ77�R���3FgGTHd�X�[�R�A$�a��nxP����M�\A*GwW�6�E��J��ȸ��4�
!�~���S
 [���Ɲt/�N�Ye�':
i�`-!��6�"ǥ
��&�\�,�0uGB@C�2�X��TK�����{ܐF���a���A�ؗq�a!DM��Bht&��7"q~)deJ8jw�p*���e&h��kk��%�Q�bFN��@�e�%��b���s��5)���f�^�	��>+��z��IdJ�M��l�	��%�d)f��z�����]T	]�3��hK���P�H���t�PO)
�&�K"�58Б�Ntܧ�h���p+�!�æ�H��<'�� B\'<c�a��Y6���L,�MY�&m/RA/�'G������tg�I��cQU_{- h�����`�d�PK�:w�����/j U$M�ҋ��r u�P+"!z���8��ˮ�.Y7�Y7�5�|��;�^��	���@`�_s����n`i�>�kt���h�����>g���j��`Uj�P,�1?;�����?��~t��}�K��S�Y�9pT6�t��3�3��
RC�i�U���t��'���up�uo����p���z��z�{6m\�M���=8��n$�ADI	-d�-zH.rD"H�#Zh����NkU>��A�<)��Ւ�.����m�ؘ׆�3�����r6ڰaz�Rj����γx��4�#�H"��ʋ��9�;���rZ��y�%&=�U^��E(�}�z�s߻qх�05��3�?��=���>��Uwg
w��v���wc��a+�y|��G�/����p��;����5\�����գ���g;3�\�!�{�g���LGK� �ݛҲ8Ш)c�����;n�'~���<��c/����m�e������1E�V��斅�F:;d��EU��w|���w�v�o�Li~�����=�����UV�yN�l�m&��� ����R|^�#N�ⒺQ�;9l��{�o��RX��J�<�=��kY���[ �����)-+j��-����=R����p��:�hjN�\�a��	���;%�W���@�X�2� ʹ�M�����b�B+��X���S.鰩)��� ړF��$������G8�@,�B<��(�m6e+�
�̀6ܸ�^�l��cN�NM6���:[r>��q�|�k+A�4�<̔�C��,���������'1u�Z�
�bJ��u�]JԠ�_�K0A8<b�ρ��4IŦ��� tN��Pۏ�;/��o��ս83?#M����4� �~ �����h�MD��6�BWR�������Ё#GO)|J��V�0�����;�f�$�)D�aD�@���
r9���`l|
s��j�9TPP�ᗗ#� ��D�N���B_��l�@��B��9�M���^D�v�?} �m,� ���RU���SDg<��kp�%c�'��癜���ѓ���UBAu*�Ė��~x-�QK�\:����Ĉn��"W(��ֱ��"��7թ�c�@�1Z^fHj6K&����C�O��СCr�ڴy#���da�XX^)��Gq��8���B�J� R�'�cx��V��[Y*adt����^��|��Fw�Wԫ��<}�YLL-�����[ab�;Q��TJ(9i�/:�<D�6*��{�vu7A
�9�zQ(8�dȮ0!3�Ņe��@$�D4�� �Ŏ�<�N��=�Fn4
adc��C�"9Ф �wJ��{{;0��_M=�GGgpjt��_��6�@6��H�����:�qY�+lByƧf12>��SG��O��
�m&)d�N
�������m(%�1���B)c�mn�xІ�� I���@(�����@ 5\�n��6_�%��V�D+R�'��v2�R>��:hy�.8⢋&����:��4*ED��6�Xɮ耎$�BMrقI����SB�b��H��!Fa;*����WS`\*�I�F��8M4�M�i5��xL��Z�P���^^���3Pdˁ?�蔃��l�is�4bkj�b���i�[O�ZꏂZ"��6���5�(:�=б�Q��c�-�(����U�Dr 3'`{�M��Y7?�<iF�En�A��r1ۏ*��'��'���8G�]Kх,jZh�`6�DUxﭐ�$�l��5S�`�DEj�d�{	�kDݘ��d�N1�q�K���V����A��2�b]})Q����0k�hl�"h��B�
��@k��3HM�ԡ=�7 B�R���C�;����9�!I�]��6S�qD���-��b)�\nK�sz���^|�T/İ��q��}
/�rDBu!B���!{$�P@]��I:�;|�֭�e�\��`߫�g�^7�%w�u�W���W1v�B4�`ѬWt�)���鍾�l1y�s��AW�k�k������\��@����h�P��B6�F�RVƃ�j5�K�Sd�[�?��ՇF��L�����R>+�l�y:�L虛��G�qp���y���`f~���2�~���7�[nƎ;t���x��]x�'�������V|�����{�u����W��M�����/�na�~Y/8�_|ť���+�th��:t�j���V��/�_K�]/���}��p��8���S�mY۲3\I/ ֑���.D�V�����,V��Үw�r���^��������EŭV�����̝���K�A�g0�هۈP)���ف���QO@��(��ڜk��f1�u}=x��7�査aN�6��s�����Ș�ރ}��� ���^��"�c��n849{�Zh��p!8ׅu���6�j�9y�p�d���(��^�(�w�p2�*(e�1sf�'��Y-�UuТ�Z�d�.D-�7]�n6�Ąe��ۂ�v�`�d
����n�t��G>,,�ZA��Wu�ׅ�6�2�����jk(�fڷZ��`Z�q�ǈo����^�?�ܖx���p�yQ��>�����a���h���Pk�S��i��t��k���p���4ˇ;/��~;��@��.1�;�Oh²<(���!ҙ(�ꊪ�*���z�"SG$dÒ�;s3���"zc�3��D�66�Ī�x=55��H�@P\T�QT1�аTffVpz|JA(l�I��cB�^r��L��דĪ�P�G$�T��
896�#jtHu!�l���T��rų���6���l��U��X?D˽$��{�Z�PǑc'p��i8��z�fh5�ߺ�D�BY�U��ss3�}ʲ2�G&�G&�hzfN"�������硧�S(ii���q���SiG��c(��oڸ������:<���z\�m(�B�it�-��D��!�t'u�
�&N�k'O!�Oc��\z�6�R��5�+��~�;1�F�BG�_��|��U*g1;7�5�{������N��%	��In�}B�r�U�e8e�b{����+�*ہ)T��a.���vp���c @퇱5$��6�`¶]�8�z;�ۓ@���E�U��-���I���"�! G��΄�p�'�]�^8��T���]crcSS�n�{��O��������k��N��+���*kl�����$��$�c&���Pn�1�\��^G`j��djwH25ե�ᗕ��{���Tu8\)ע���Hؒ��;e�IW`o[�V%���_R�u�/`˸�Q��+ ==	D��T��Gb(�+�����bZ]��V�F_o7l���,�FƐ^)"M"��@�b�QA"ɍ���p)6��"���uY�n=]j��l�3S�a�5�#��0:1�z3�p�[(�'Qn��NsE�� �<��#';l2gHK�A�C��N���ӣpJ"�&}Kj9�5���=H��:#�����c4Y��p@p���ցH��D�2��ao	O�������(j4�#�B8�U)�K�-n�#A�����b�b�J�n����Po����	����w�B	
b����᥎��0uAoC��R!�5ëq��m�D�>�1�5�f�>�p��À�ؚ>����.�� }�@C��\5x}?v�"t6��]H2_��y�PH�<�r�dV��i�w�u��}J?�[Q8�����
�_:([��}>[��D���	ѫ`8�?�%g�Htubpx���.-`rbJv�<W6�J�׃S�cf��ৣ���'D!X�NW�lQ��効�V��'b����@�z�N���I�V��-����A���2wD��y��g��s�E����kW��\j��!��	�oP�/{Z/���ȯd���q�v�u�]���/�r1/����g����L�si<�����/�����\vmX����_��o��r/��2~��sx~��/�-#)mA�l�]�x���LL���//>�,<�v� ��O`hU7f�s���?���4F�g�J����5�ᵃ�꺫���+���	|���199^�6�/�s�M�������@����w=�Ȯ�x"���^��1@�=��L:7�� ��4�Q��p.ں�i���S�֡A��-7�k/FPj��W5��Uiz���p�t�y�0^�(HT�@D�J#%4(�~cIȁ 0[Q�x(kc���;�b*��%$N�-�/�Y��΄����)L�����$��4j�,*�����`��c�Í !d�J��0M99�2�� `����΀|�G�\�[�n���mH#o0�"�a��҉����x��)m�kHkІ�+���`hqI?gn�0�5���z��!T�E̎�c��a��T̆Bn꺿D=���ꢢi(��|bQ��O�O��qI���p�%��;���ITJ���SuhY+R��z����-Zs���BG<���B*Aog�3+����o�`���~��8�ɉ9]S�P��:����S6�������$��4�׬���0<���%�.����Q��|�x8�d<��x�h]���I��a��40=���㣘�YA�gÎ��?�����m0Z�s����<Ş�p ����w�+���:\����UN�����Ǳ���`2��/<[7�G���%�܌151��L�"R��YA&���1m��o=lێD"�r�dj��/,��l"M��^^&�jN�(�Х�\�Ճ}������#�xn�>,,�M��gŤ��&����\p�FD�(�y���9=�m��P/6nP�1_#:�U~���Fg�-�2����7P.�Q(,��wಋv�+�Sl����=���KC&�a9� ����ML��a�L�@��>����(��w f����DZ{61>��vaxu?��b���HA1��&3x��=XX� ޑ@ �A"D_g�09MTOg�P(~�rE�o��pt|�����B�����Hz� ���U�X?<��Ta�8������Q���2����"�P��c���� ��]����2��P"����7'H?K%��yzz;��L"�#����+�B����E��,abr�tQt�x8���.l���ߨ��Pw��0���4������2
�_t>�nR~Mz!����O�o���wu=%��cy14؍�֯AG,���<p 5���l���5z�X�I� J�{M;�Bcc8=6�ӣ9�|1Q�X���U���q�A�=�V���/�@o
����p�u�:{����0��v����<B���nXv\��%��x���1+���)sO��y��U�Ap@r�1��6J`����zV�q�l�QO��WX���UHόc�]H�0lͯ��L����׃˯���l�����Ǧ�P����]t�����scC�_z��J����ڪ*t�/�4<��6�l8B�׮[��
��=%�V*6�h�msho��0��ҩ-*n�}�kƳS��m�k�����=<��wQ���e�B�s�.�:��˩��1O�,�;Չ�n����^tu�ѓ�ç>�7xa�^-���	�H?�.�s7��z�fCC�Qt
�Ӗ<�B F3�G3hK�H�����mވ�D�ęcG�t򰘐m��;m����95a���:U!�����f�H[i���:�y�>�}�|A���cD��h���N��(��@�pW:5�4D���\޻JC,〟YU&��	�LV��A�;�y�V�҇އ�n�ytt�Uo�ʒb��+���_�?~c�SȤK��g2K�ǃx�}w�������w�����/��3�:+��zzq��nĥW^�T��k3���?}�>�Y����>��o�>���3x�ɧ���]�	�d�50Џ믻��p#�~��Q|������Ѫ��;o��/�gh x�_~�·�糯�����M9EFm�m�_�ӫ׈C��z��B5\�e#�鍸�����A�:�c��4[�8~]�����lU
u�I�/��������
Yqm���&X�I�R�'��q�}�\E�Q��a�p �VS#8|`�O*9�^6�J�:�p�0��H��\x9��U ���Ь���->y���gg�j�jh�יB��k�]�U�!�٣�+��]_��->:_R�d�H�R��������k@�a��b�*d#�4�OI޼>D�1��z�"�Lc��a���.��@��s��sC�O*���4�OQ�8LP�@�:ۋW].ʐ�׉SS�
a��!E�J%��P\G;Yc�bM�ذѨ_A_*�ޮ��R��Zu.�0=�����6�Bvc�A�ZՉd����Ï`��#��66mތM[�#��%��l�QA���G.Wҵ�DЛJ�� DwW�	~=n��p�^�/�5�,���3��Β�O[$�zV�i�s��J�$�ѝ�chu�!4ky��)p���S6��O�b|v�D;�މu����An%�l:��S�鑓�
�aӦMHu�D{��`߁�
�"�h��M*�m�|ay	�3jp�r��h�­�	�k��7\�����$�QL�-��16��N��TPY��6m���;���g�]� ���ɓ��oٲ��q4y��F�T����bj6���,�u�	=j�|���o5p�[n�@�h |����0�~��    IDAT�/�1�m��]�����v�=�eo+�To��R��wW!u# 3��|��eF^)�)��Յ4��?���R���9�j��BAds�ɑE<����+Hv&�}�H�����n�@%�Qt��zF��QA �z�62�]/��|Fn(��}1uV��j����X���(�����,�y�%LN.k��1�ϢE.�	�;���&��p0�)SS�Ng���\��t�)SoÇ��w�ƪ�nl�5!�� ����8�B��L���:�9����h�A����1����,�<J�Ä� k?���>�b%�K.��\2,*���˻�b����5C�$�d:@G!�[GW2���å�� ��ػ��;.؆���x�l~�p�ŒZR�e�"�f�b'N�`9M��q�[�G&��J��ZY!_�Y6���ѰGׁ��b�A��A(D.�ǩS�p��&�g��'�z�z��NIbM��h�{�q*c항��@R0�B�E��v���TIϨ(�5��_�ci�8�B^���~���~����
Q��t�� /@п֑�i�Cظyn��-���K����� �R� ���Yg,RǪD�~�{j�E2"B��=h�:Z.]5���L"m��CCk�&�mf1@y�Q7I���g�G[n�l�\�!�8c��z��1�omj�����'W0����sLց;��:SW"��A�Xw������;��@�j���"���g���/��498q�~Fu���f�:"6�=\љ0F� ��>,����Ɵ�}R�A$�r�#���C�(<�"hzV�"3�M���0@jڋ�R�$��� c���F��K���L</���2�y�X ��a����@��5�F.�R�D��>�!6`+{���*h��'��1�3�/aq~I�zL�E�Y�x������_5�IF4
 f��x���؏���c��<B�s��Q��q�.�{�{'�t��!ly0�/�����tx��W��{��M��T��v_�ڷ���ݨ�*B����k�g���hg<1���N�F��T�!��`�.8�)L.7����;�>�c'OU����w�~ӯ|���u�ݸ�����A����������w��#҉�T��h\o�D��M#��6=��%����Ӕ]g�� a[ظ����\}�H�Z�&K��]oT�-UQl�X)���{�V���� wڿ	frc�h�&*:��6ȌZո���q�K�V��b�:m`U���>d�ǰ���171���ÎT��1M��iB�\�(�e(h�)���ᚠ2) AmVX��%�kx�&5C�&ov�Z�S�X�z=�_t9����m��һ�EaG�ߺ�rr����,�l\�rR��룭��pW���vt��k(��J��I���e!��ǃ���s�J�Bn��9����8(�Ȁ$
SQzh�X�r͕x��o��ߍ��Y�
e��ܐ�Ӭ{��� Ű*Y�z ��򠳓� 6�bU�V� }����E�-fP�02��W��w��k�4�uG��Sa{���|j�E�XH��u�ѩ������9|�)(Ys���}_bazR	���tߵM�z�/50zf'Ʀe/���k�>�H�a3��X��QUB�[WW����J�Ь�Q)��҉�?�ۇ�?��<N����F�`͵�V˹�U���/`��&�Ǆ��R�����~�*��J����XZZ���شa���|�X�_ye/N�%��DJ�(�Y$�~w����L!�+v�6�8ufϿx��I{���Q�p��q�CB�?3��S�XZ(b�*�O�1��v��54@���brz��ڏ\�Q��F��F}\݅m[7 ��XY^Μ9���qN<� �ǚ�==�(���$:��L��q��}�Ɗ����Ӡ�Z/�Rq��-B>�a?ГJb��]Q�|V�6�.L�022��Oc9C?z?J6x��-l\Ӈ�ke-k�~_Yѻ�C��W�Z��bS��B��_bp�e���Aф�����"
�!��P(�R��K���{��DO��ִ��6(JeC�dN:��-r�2nE�K�ɢm���>7�46`sDKf�oD�ZUXؼi֭�Ҷ:ҙ򅌆�h"
��]���/�3g���}�狸�������|("��r�̲���C�e�������'���p�5�chh����E_=xL�=�o����O������	\�c#���=ur���f���#Ea%y�&?���Ť"!R�h����'��ɩiL�M�\ɣ�ʡ�/�[�|R�8�BU��"�)�E�@с�1C�9u���r�OΠ�z�mv�4*^s25&�g��7��1��M*��jp�>]+	����֜��J6#W�hЇjf+�'0�
��~�#ز6�}������+�~�idV��.s��$֭��o��\v)�y~>��@�PC(�)�>w�sa�g�!�H��@���h�ׄm�o��1�����8�z@Kj
�����������`me?��ݭ�@�X9�H�m�����#jn�������"x�Mb��4��ɍJ�*CO�ז�MC�~���]w��|׽H��K�����/�'�y���YVv(�)H>��Ss̥#u?v4�@$��&����M~S?���U~`�1�z�P #�bi|4\��9ixd�*P.�,�ݶ(f�A�����4Al����U�6�˩.�b/b�]���+�́��R��(}�

��EͤO��y�P,"_*��g �V@���G��[P�����Eh�+�`���p��oEgwƧ��k��x��gq��	Tk������ �_@8���;/�G~�Wq�e	k��5_��$A�i4J<qf�����O<��^��w��jo���{p���`x(��������#8��ޱM[X�a���}�����d�Y����=w���~�?IŤ��W�|�W���������ݶ�'X�:r2���zx(L1�pqֹA��^A"hc��a\�e8�0�a��s�`bi9�K�cH����gO�ɗNb�D�����!=A���`�⹁������a�ZC�n��N���v �C+�H�豁X�����8��Ә>y(�h���2t?�V>�
�!�� �cnI
7ZH�:M��n#�X4�C(�9&T�ƥ��Q�;J�<A�H�v\��;���F��G��@�1օ^+$G�S������d�Ñ����
WC kFZ\�.E~�_�KX�����(�͡��{�`Y��Jou�9�нsN'GD� D� )�$��#���l�l_L�/\e�G㱲,��� �� @"���sv�9u�ݻs���~� x᪩��*�sv������}�zV9+#Z��iLlbV|��_^�Df�h�L��!���>���QL&d�S�##Z�l9.�P@rT]Lv4$(�t�s���s����素�ÃF����(OR�j,؏�����b��̈́���&{�淊������	�]{��щ'�V�u�����`��n򰺸�,9r�@�Ë�pP:�6����z�T�"��4X\���`g7&��Z�N츪�@2=�gi��B�h�A����oB�8���̺BAB���C�������f�*�tyD�Ƀz�' E���2VW�ఙ�z��)t�}rm#�4~v�m��1LL���K�iJ�R���W����d� ��!��er�KUI�jSg����o���̀�l��+�l���]�s��15D��.�ccu�1�*&�u�#�F����Zh�p��p�XX��?�	
����uF��L�}�v�-��9E�1?���IR��<�X�����K(D�N�`h����]��������|�,�=�����y`�����S�:\z���i�U��r:P�g._��0����>�Gi���k��P��`����x��p��m����&966���~�ku"�$ֶO��Y��o�`7D������X�v��NJQUhg4"�-��g?�g].J��4��h�e[W���I�k� P���*��q68�k�l��J2�=N+N����|
�Yx`�`{g�RF�6�&�N�v�{�1�|���Ο:���1f.���������k�@ww?�����l�c/r���n��uɡ�f��$��+/����l�����)bl�_�D[P�T2���%�g(ݚ:5����l�l���eE�Ti��f��a�s*Q�q,�\��ͭmll�¹�ˍ��~�=3�F��\�,����34���u[���v�Z&��'w���!�p ���(T<9Z	����f^&X���xM�%m�	�Ev�9)���5vky LdSR(�-h�)$v�v�o�����QҩV������K/�X��a��:;��c#x��O����x��W�g��ć�vBg��'2���9��R2Ħ�L8�&z��Uv�+��s�Qz!��g
Ї��^) r��R0�<d��}�����9V%9�<O�ϲ 7%�L#���X�K����;x�E�qӐ�&h|�~N�����9� /6?���෿���lC������?�K1�r:��:��0�A���hP�l��$����g�5�I���`�YI%����g�f�΀6��4���
�f<V���U�$��\��3�b��fWi��PӖ���LdJ$�����{u+�^�M�5`!���_˰6���Ry�z1TU/9�i��P㟆��A��C�X���L�㣄LJ)���<�jU���?�4&�L���}���5i��O���I�R��3N:�&h Ԏ���Q|�����ĄH�9Qk���ǒi1�n�Ń{���؅�jD.y�\� =�~<���מ��Л�3[�V�X�71�s�_��n4���8���K�|��?�k�����s���o7��ɗ����?�ڭ��(Tf�]�H��u!ګI�t9NV�2v��R��a2���8����`w'�P|L[��8.�ɫft!U2��7��- Q2h,ߛ�7�w*?��
�t̌hTQ��$���&:�+b��0PR�e�F�F�t��,L�pyhD"ĉ�-
Y�I���4Ȃ*�UAj$��j�Ɇ��v&�R[, �O�!��W�</�h��"1b2n	(�k(&�ӏ���=�@xP��B�T��)�H4u�͗��A�6�^65v�՘T�z
sJ	���Nv%���%��L���"��S����W6�A� G��M����fA (����ރ�?��6��₣dQЄ��TL��L�zD���*�rJ�l/������P?tu:�SȔ�4�X�<���6�<.�;]�������9��)ܸ5/D!j�9���lww���W���5,�-Jx��@^�#�Zd�R8Z6�Xk�f2��+ֱ�v A<U���)���^#Ӧ%ۂ�O5�.��"7��q��:ۀX$���e�j9��~�~�2eU�%��w�� =�b2G�p�]�|�j�E��89��e��`� �V���#Qܹw_6܉�~��E��t�%	�I&�8If�J�L�P*�@��������`��0��l`?ǭ;+89�.�	���sEBb�G����@&I��*�V7����795?���H$c�A�wv��?����//"S(+]����hkwcx���<��P�j%�����E3o��w����4��0���Ϗã��wq�
��H�1q�F�跛dQ�!&UL�%�W%%<NL��;�B�RC����>��8��9�/걱u���C�JU��lZ�m:�t�^��"G<��_��ߗ5hhh ����j���ű����hWiu��@S+���'R!��&������N����9����pt\�����+�e��:eT�����4��H-�J�!b��@m��1�k��Y1>6"U�F�M}��.�t`]��N�L#��YoC�0�Ņ	,����bԈ1weq��ޖ5���abl�����������Y9�\�rA�O(A��_�>����|�ٽ8���a���d.�G�M���4�,aeeU��S���1;��W�ʄ��*������Ӟ�V�7���������OȞH���A���X�[[8<����f����z����D��W~�6^�v�f�S�����F�b\JCN�Cʸ�:��:/a�J.ЍfN�t�9X-�%<�W�+�Id������/����iS���o���\���_�I�����~�>�s/��Ͽ���O_��7���i>��4�kYpO�rrL��y<O�Z""R���	���:��~IA�W�Jq�z)�lu���[�4<�AS�g�"�����>����J,��ʦ�;���*:D�՜��� 0�`8�i�k�XYY^���G?����Ϣ�o{�������_�5�7:��D��!-� �h�ިe�7��i��}�,L,l8r�\�>	z6��(屵4�'�l`2P��D2�K����af��I�R�@� PCRy-Y��-̫�R-��M��t�&�j"��_�3~=�������&��'�NN0��R�1�p�!�+��()�sk
C+�o�j#�C�"��@��K$J�Hd��j5B�+#�"a/#�5��W�`��½}�))�z#�b���7#��Б�b�	h���dS{hSLx��G��c�A[G��r��zq?�����p�!�/�8�G6�-������>����]��J�����%C,���o~�[Ͽ��ԍ�>8�(�٤Ԇ�TZ0��)j��*�d>v���f7��&לt��Á�����pO7��;�ҕU�N�$�A��#Q1��?Y�K����`dѤ��'�����T��
<2�90ƲZ��#�:jתE1ji��'P8����<�V�ЈG��4��j�c/�Ui5�eq%bMO}�G���KI�l��h��}xģƓ�G�d����¹����j�h�8��j�05Hα!�� ��@k�3<�ޱ3v��3�(����d��u�AT�14��cJ�F������n�C��(����P�R���O� ����pT����mH�Nb���h�
Tf�����*��Z����{��U�s~O������;>a��H��**߇<rꦫ��{O�"D�F
.;�'�(dO����p� bY��-�5&<����^o���@'�{���
͸w�3o�\��ƞ���vt�hkgGڋT2����5�!���s�NWF&A6u$�Av�(Kku���@"Q���A��{2:�6]�S]�]��V=-����6�lʢ��2�R���>��XG�焇&=���F�#k�Q%R���e���S$�$�(��<t��݉�vv<�H��0r���8=Ot��;(]�|6#�k�l��0�8�c^@��LT�>��N��`_#�r��ݟ�V0=����(�Eދ8\Zt���#�D6S���6��pr�@������p{������ڲl�CC�u ���νi1 ��I銱k�n��h'\.;J�*��g�t������EѠ�|�͎S��zm��� <n��i��*T:�Zi��#�N�YfB�F�x�XH��R��6	���/�B�H</z]]��v{jvw�Ba��`����"��mCOwH~w��E����#��02:��+�zT6wP�ac�I���,�,r����"TE6)����,�۷���l��`��Q��Qa��bf3�5���t��>��5�M~�d��6�N��I&��������3$�]�d"��o����%Xh,�����嫗���Ij�ȉ4(�u�K����%�L�3*	J�N��ٳg�ibg�2�;���+~���R���ul��p��<��$�8��$���ù����k�p�ނL��>3����6���ݝ���UٹU	ӝ!Ν��X��N�'2;���Y�]�2)E'h���j��~���C$Ri�	ٟ�����p��)���T�r������9��bwAk$��!i8MU�7ʆZ�/�!���d-���Þ�cVP$�@�zI<�����������م�c$RW��K/�_��7���"����q|�K���="�?~�ۈga��`4X$����a    IDATZRu%O��Pn��Q��:J8���8j�WM�jʑH����R6�D2��Ha F�tZ�ܳ�A~S��½%�ly T��$V��"��r�(A���E�aD35�6
Z]t�bI8ZC�	0�`��k�0�,����	�N���@$����bq�U���	&L�SA�6�C&� ��DԚ��P�Y���1��	�,)�cs�QA�ߏ�P�T�ӷQ`A�#v�\��dm����Ţ�ϫ��2����hu��ڤITR2�֤�U8�k�żZ'������,����g�J5��q��ǂ��@+��F�H��S�������lw��lC:[	0�ETZp��kN�Z���S��d����R���OH镰�L�$��!Ĥ���
0<1%��,iK�u�O����'n4��&�O�B�*3Vb��(抰�m��B��z�Y�x��'>���>���(
�+�򙨖+�z�ڿ��3��׿���e�_��\P2��닏�uk�+��6wP�#�3v@s#V2��]���"�%nL��x���T���{0�����р�P�OM�iѣ·��"������x��s�����i\�q�VQ:���&~-��4��7��n��8�r�qk'��\�Sǈm�"������9S[W.����<���x�L���ӭy ,)��hn�u�`H^GR4�ݤ�E��)!���(��9�(�f0�a�[`��a'eH��I*�|����"���/�
e'`�"Ǆg�H:�CFy��İ�a�YEB`���)�5���ڸ�N�Z�����Ʀ��גG�R�$�p1G�Pݬ�9)h�	Z&�&|��� �8f¹�~ x��Hj��:� ��EV4����Hm�*a򢘾�[TF!����´ A�σޮ :N��w;
5�p��ֶ�sF��P_ �'z�2Tȥ�њ��5D�~�ά1�Sc8uz�p@�������^��^.��c�8{j>���2��0�c���������dCc�����$Y�X��d:�'e�t�f���w	��zvs^�I�����U�+7�qp,ґd�$)�q��b0���!zf�fF�Cr
�@��`6�pt����*:Bm�n��G�tEL�L�e��i,�HO��y�?smKK��j��h���x�h��"��bfn��.!��U��χё.x<6�0�2UA`.-��Q�?���S�1�`��޽��Q������D&W����`J)]��h`(�KF`4jE�ArN._���2L/�f`�3 �,�J��L���]�bY��9=mY=7���M�A��%RB��<��Yx�.��_R��VJ�#�	���Œ;;iܺ;��}�,t�u�������+ގ��Cܽ7��è�n��98Ї��Qx�N�R wqy�t&�N�QL��t�t���A��1_̉��0�83ӫX^�E�b���B�d�c2��́rD6�L���@�y�@'��Tt7�����J"�������l*���9D"��Y������gN��
{K��0��5��x�>�.-����(�2|x��et��Co�#�+�A�޽x���$ςE����8nޙ��ZZ��F��05ԁ�>?��F�U���ܻ7-��C_D� 3B����RЙ�n):�L/U���x��gE��:ꭷ�q��M�F|�ɇ04�#��\��%�[�D�h�XD�Aii�J��;wJ�&v���u|�_~,C��#>	�l6J�xyw��ti���VwW��2��P+_[�Z�0�א+�D�kF��)��w>c-��%�vu�tmue���o៿���X� ���|�._�s�}���wqp�B
�Y�l���S�Bo���$��dDSi�W�.� �� �aX�E��.#��)9���V͎u6���z��>�3��V!�2K�q�{�l���E� @���(s"��A�E��p�Iͽ��P&�=�5M`A��2I_l����8�ư���|�-�X(g6XP�jP*��@�I$�6 ��`��`q�P�^K���-�Qz�'�*�ג{�	��\ ���Ӹ���ى2Ǹ���8��������	��,n5e�M��`�i����R����ؒ+�+��O�����8�&etWh���L�O��xB��F����jB����fa�.i[�U Yij�*MG�
M�5#2���@��e�V��tV,V-\>����_����r��h2���e6�ʔ�Y�������fqbc@�$�F�
]�� ��OP��X���g��(Y�ڍ��6A�'�	9W����T�i7��ۿ�������/KA���Ǚx׾���-��o��� ��Z;�Ŋ~Ŕ�cTUd
d�V�^��B)C��:<��#x��K�d3�^^��j���Sҙ�R�+�ś-l�d��΋����k<���R(��^
�^#�d�"T���\n�t�H қi~�I�'�2�!���͹�[�A�hW$B&]�JFi��PR�S۬f١恁�o���z�H�OP�7V'SW�[d;B4�ԑL�p��/�!�X�4��Aъ�ll�ރ�(U�>�¤w����"쒙"Y����h��3w.>���F�Z�X�?L��ia6��#|d��%��.�*.t,��=Z��ʽ�(�)Y���E�QL��9�]��95i�H&��Y9'����F�K2!�?�U���=�>��Hh4X�݇�@i��YH��Іd� m��X�^�CM2hʫ���sL6�ӁP�z4��*z�lD���'�,�E�6�������e��Ƶiܼ3+��p #��ҥ65������NDR��^'��0>Jf��|=@2������.���[�h�{�G��)�ٸX`R�/��f�%D2��~���P�d�w����F��@g���*S�D����]��E��v�A�d/游7`�vU�GN�t��ЋB�mp8\r�&�5�ctr�<�شR�P�+Ι*���ܘ`����E����""��5%�xj�CC=0[U�s��>~��H�d��Չ�����ˢC����ܝ.4l��|���\.�pѯ]����	��066!�Ζ�"x0����Ⱥ����ȕI8]fE����<fVqf	�Z]�{�B��̞��l^�a�	'�idXUUϊ@XЧ3
�K� r��]����i�`5 �bC�Ca��v�N�ɋT�����N/`� �NAp��&�:�K� �?r"��H�X�	V�����uS����s88<���	Y�߇pWH>�j6!_����@�Nz{�`���ŝ;����u@o�#�m��b�<T�bAК�n��U���NL�<�p���&KeB�A��n��9-�ߢ^-"�K���9�����{[��%������c	<
�BB<���������3�X�9=)��T��x��ٙ<�?���A\�pJhO��7�w��7��/n�ǃ��0Ό�=j��	�o��ʏ�*_Doo/{�C�lg�.��q���r�7,�C��+�>�N_��sx��Y�oޘŽ�w���{/�3�G.]@�f���1��_�q�2+Lv��!T���i�
1�.���e'9#k�HN/C]��5X��M�U�ۚ��|ɖ?i�:[����f���Ke���+id�k{�?��琋��</�?��䑼��W��W"���p��E|�K�
c���s����w$!�	�0\M�M
�L�k�W�+��<��fA��D�R�F�<s��Jm�vLMM��#�J�����D�JQ�!R�������չ��y�[ ���ȕ�3��f�2� ��� ?�p	l���w(�p!vZ�N���asB��`scW.+uJRp�4ACR��f�hVS��w���ցB��t�����j��J���˺��%�N��LBbc3��Q�6?�r�\7��G;��4*��@_��ǭ�����T��]�U���P�U���-�?����De�����)�d��4���˯e�����K����R���� N��f�@>
��4n(K�Ǣ���V���T���4p8e�XFc�����u�:N��H��פ$�&J�,�|T5�vBa�I
/��l����H�Ȕ��� �l�LR�Iz8��k�J��=e�:�n�o�.���J�c����Ư��������Rw��b�����7��,_{�y�{]���&��(n5���U�-%5b"�NUN�	O}�I<���Ж��o�A9����qI��1L�� �	9�ѬϽ4���- Sw�d�ʁ�o޻���Pe�Xe<��n�mFǨ蘺ȉB.���װy�.��LFt$��<[�B��9q�2�a$�O�xt0�-H%�0M��C���]*�N��������!�旂���T6���UI�㡘A4�>c#cx��G�����ӷ���X��E�fG�F6�M~f>WF��z�a��ox��H��X�gp�41ͲA�''q �2C�(�"���LN�J�!��dC�PAls��s(���,#�%ٕ;N	�ΛW���N���(r�
��mN� �T��
�_�4`7��S���4N���A�U&&R�(�����TA+k��\_�|��%�z��L�� ��i��b�WV�NdB@�Y�f�uy��H ��ۉ�x��� ��{s������3��f�`���,�-�n�#�`l��9E�4�fH�	��G�PIL\��5�J>�]��֮�z�Lv�yy=Y�dԩ�5�<<�ΐ�m�È�]m��`���dp�bek;�8j:r��2i)d�����i�&�ɏJ9#�6�ǅr����%�-�
�}��$�=tv͸y9(��D����pphn���.�lbieSR�y�vXM���� l��5����?x��$zp��(�V��S���ū���ݽ(�/�8��gƄNA�0G�7n�����PBΝ9��.��~���+r�����ۉ+F���_�X�~,���}<�_F,���l�:	)Ԉ���@� &З��"��Ҽ2�P�s9�VS�j�Q���y�.���qj���S�mC2U��a�f��{ �Y��� .]��h��tQ(Yѓ�V�;II��\ʀ��{�����8����`g�P�=�ہ���T��ISG��[[�B3��̙s�z�������i�ǡ��`v��窮kɀ��H:�� '��~ago��[�C"]7}u?sc��%��٠�l���c�C�	u�^)I1������ya���L�:����d��M�Ш�y�����{R��V�+;b<$����qLM��u�98���f���E΂��h?���/`G�����%ܹ5/r%^��������ԍ3��N!���:dB�p��ĥsga��q���ebv�l�����u3n�\ǝ���Иff���,�2�
qY�8���*&�K
Z��
i7M=;�kZ���6�@"�h��n� Ǝ��Z���]`LZ�J�z%PN�`�Á?���"}����͟��I�s��~�#��W��u����/���������=Ї�|���˿�2����BuZ�by���� x~� O�#ͽ�Yhi�.�0;!�5M�4������#r�B�a��YeM�F��N��-�>�_S��*�o>��|)�̇�$��v��K���!��R��C�dT�13<Ou7��O�3��sf
{$���z�ܯ�6��d�d�Lɖ^�P�}A��av{$�9���D���-v�~��$��ب��OCW&�4����A>�ģ��s���K89܆����9��yhE�BI&����Y�<�wx��!�@�(s��~>-iZ�R$�BB^5u/�"9:��H�(���g�;$M�P����������	��1N�AS~��o���F��C�8��1�^��J*��K�Fy�������&�>6C��2�,^?�VN��a��E��4����
�"�"4����z�2�yʣ-�v֫y�9�t" �K&},��]+d��e+��~��_����3���(�m'=�{��?XX=����X��F�8"oR��>0� ����� a�|���Ȉ��ۭ&I~4jjx��y|�#���\�E�(��&�����;�$���n�FD��w_^ŋo, Y�f��X��&dU�� ���3j�2N���`�S�v��Q���F|sso����4��� �0٨D����Mi��?L�s{<M�K�UU���=�>���E�n�ı�����,ʮ"Z��,.�dJ�p<\�c'�f����������,��O���7�!�.ȡ���F�1el�4F�1r������+���a�@g�y��YdA ��F]�b6�Iu���)3�f'��g���7��77��Q3M�:SUȁ���EU�������*���4O��,Jy�<����SE�^������X��(%��擲�_U?K:8����l���@CmA������D#2�lI���}�j�e9D������A?B�@�\��zG̿zJOFz0:���D'��������`jb��������#�[��F��~R�/�P�0���������[ZC:W���@(��cϢ@4�5�?u͂��5�(�y�o7	���'(]���v"G��ĳbf&��׭�t�|n���]�EW؀���lH��z~a'��l|���yEOZ�瑌cmuQL�^���\���(�3�)����׶$ �{a�c9�?�B�Ӈ�H������G���プAYv+ҙ<��[��S��x�CS����ɕ�Rb��*677����d���XB�����(��q����lL�u"ɘ]ZÃ�ud�e��.��p��Tؿ$��MF����6_>H��*����+�/���z�[&T&������V"&��3�8}jn�Y��QQ;�X[߀V�Eo_;�zC�.QT���=<$!��`���ccr�)}>�ep����	�Պ��.��#IH�R���*n߾�D�.\��+�jv&��oO���]z+�6r�*$_+͵E���T֕w����N�ayL��(=5'/܌9M�1���:[,�:�x��+�ؼ ��*�X_]���"b�Q�^LL���ٳp{�R|��?�M%CVX؉���i�f����x���x����X^����:v���w���3x�ҨHV���p��}lmDe-u��t�,.=4	�C����L�v�2�7��^�( �`���O��æ�ݻ;X��A�S��n��c��/�r�gw�5�`�;��h�da �<9	1�Ƀ��hC�؀�`�É�h�*P���G��y1����1�3�q����.c2�*'�2T3hd������>�IT2G��_�)֖�ȣ������������?����>�0��̳����s��>����?��B��S�j��J6��3S��eo�c��R����Lz.�.Ŀ���Ȱ���?9�	%�V���s��"�ptY@���߷)�R�a5�c��2�R�����r�u
�J���e6�i}��V�"�IT�F��<���0"� �R�b&�[�Uv�M���{�R�E��ꆯ�%�N��\Q
�|�t�0�+%n�<��V;��(*��l����ӿ�!ԫ9�����ch�g��a�[������5%����L	sQ^������M�wZ	���g��f�Ψ�ୂ�U|��P�,�	AS/e�B��)�%���^ht����b��8.A���9=AX�~�N҈%�Ҩ�tu��ſA)�*0�B!i�nm� �w��HM"�Ĥ��f@���I��{q�Ԥ6Ve����f��j��H~n��U��=&��R9�P�I�rU&�����Y\�k0hn�Ac �*�S�]�ƹ��r��U��|?�§�����7)
�o�Y��/�����O�kz?�����F���
n��u�_T���ne����fW���Z&��߇>�8�LN	<�����Ϡ��@����fG>W���FIk�qx����HU��Y\��q@S����'��+Y� �*լ��f��T����m.b��[Hn/���L�$s�T��W���ެZ ���E`ww[:D���'p��9����pc�,!���)�4q��Ź����C;�H7�F�PW�H�fg��˯�ڵ�8؏HX���=!<�����׭RC��i,x��e�V�
    IDAT��/?���{�(�z�,>�E����8��߫"���$���Q�$����ý������$`vP:�`4j��V�H���M���\4¢�EP�Dm]uZ���+�����x�����E��VJ*�L��¹W�P��Y����P��cj�J��`��@��!�y�U�	��X�afq7n�H�����s�3��4�r�
^��[XXބ�bB�HΜ��㐢�>���Cl�n��qx���^�)�)��� �����S�F�BQk��sB��G]>5��X���!/ɪ�4d��7R�Ҁ��I.Όb�7 ��^�;{��;D"���e��̰L"#����n/���ɗ;NJ�����=�ND�.��v��H�a��?'�I!����ab|c���!W �Lo`~i�2��̂h���A��@6���̴��z���8���8��[�������\8���&�̨�d�u;;{(��2ε8���U��鱾z���M	�
�����Z��>w}���IllGp������k	�=J�t,�h�ePUM��8!(�w�(2��GF�p 8@ǿ�֫VRL�T�<F�:&~R�id��6��+S�����/6��ְ����*��y^��{��)�t�n��$Y��щ���N�`����hC8��Æ�n7�b����XY]����@�c����T6����n߾���=\�|�>�� I7����^dm��C�TCC��$�i�;6A-S��&~�heh2��d.5gƢcẠ&�����-f3�y0Ȥ���߁s�$�����ۍJ�p���R�6���c��B�ZB^�L�����R�̈�do�}����tįE@������I����&�Y���'p�t�\�[���V�ץ�nz$�ht�&���7��w����'��:fs1x\��StM6�ϯaog��cc��+b0�qp��o�ca�Z��	SM��-u�Q�n<��Vs$��̂�F�:~)M�V��]����Jb�.�1��YH�ٜ�X�6K�{�!�vNC�l��_��3HF�eB����wv��~�����3��~���7��ن_��3�·����?�%P7�l�i�.v����yI�g��N:'�ܧ4u�z�[����-��$J�̜�5�(ܣsY&�s-��in�؟��q8��Pm�!�d���M#��Z�V�S�Jp�FU�ԡ���9`�Mˬ��r�3P�}L#k]ܫ���Js�RX��#�q*rBɦ&�5*1���{`��vd+5ĳyjA9T�	����j�p��Rd�1���q�!��-��g?�I��ʋ?��?}ϟ�Ǟ�(6vvv���"�N����}�ȃ$�ѐ4m�����
}�-5-�4�̏�D���(�%� 5�2q���>��<T�at8T�*e��1��a� ��9X~t��$G v�b�a���g����C{���FƑJ�1==��u�*��G.�~�I/������٠�^G�kJ{�;���"�����ҜN�{��z�m��d�oIr7�TM��B��ϔV�
5��͢�ׅ���Ieh������g��?��խ_��໋�������ݭ��;=�'�|���:̨V���Ұ�pYU#�9�Q|�pg~�pVn�4�9�p��0��a8\حF��D�c�����AN�e���/��7��y��z���Ȗ?�5	bEH��o�C��P�1��#����*j�v�ag�6��BS�èeǊc>t���{�8e<&������l.v��~����'�4#.Jϙ-Fx\n�ص���Hw%#ЪE��21f�<`�S?733#ƥ��ff�E���މ��!؝6��A���I�P�.�����������|0y:��1����Ei��e:@������"7���*B��a��$�� }&�GY	U"��]	{Q����"�O�.��X(�_5#���,�^y�Wp��O"�m`/G���f
�lX�Q��C/AS|(T
nx���0Xc1 LA��@��r�:�ev�X݊��[�E��v;18Ѕ��0�:ݢ�7j���ӗ��<��s�w��.����܁�q;�Ql��gN�HA��W`��͕�LUa��eщD�{����\��X<���-,�1�"�+]+;2��	AC�������>դ ��G_W���"�����1)�5��ex]^<�Ky�f�C>���-0��;{G�d�^��qV].ޅJ^̪��	v@�b𤶳��v��P���"�a�|m+���M�s�<h��Po'.�GW���1v6�d���p{p��ȳ�����nJ�����p���:�)�!0h� _RYLY�6���P�9OgF�0�?{���.\<�s�{��T�cg?.~���"�\~NҘ�I�5ʪ˦���&� <�j��-�N7'kʠ�>� f�����:D����4r�����)��N��e	&K��]=�b�v�;^�u�/�.� ��%��kH$Ӣ���mw�����jT�8���
v��Y150��Pn������g����t2���6�l�����N��W�p�k0�\�5�%�\�T�5)l�T�9��@�:J��a24K! �|��`:+R��n��dB����8�b��P��0��ŹUI�&G��+�$uYc`�gE���<�)Յz�p:m�ܟY��7��U��cw[0<�g�����]�F� ���>\�r}.DYܙ���{���ȧS�h��}ｌ�	&��}��[XX� ��HP�*))��b��k+�����cd$$	�����O�bk7)�N%˚�j��Mj*��+F|�IjY�a�D�J�Sv�i�U�3R�R�IxFUo"�Pa1�t�9iU�<NX�)�5k�RY
2��2G;������������瘹uC�O�������cW����}��⏐L��ʣ��������_��9>+F�IR�'@C�C5��$5D�ǉ�'U�k9����I�⤄8L3+
I6W�L"���)��O�D�/������$�S�9��3h�y����0�_�����"%�(@	'�Ve>����J	�J�6�h`�W�
�I��4dH�1@gq@kr ����2b��3C�J�
n�.��6h-d��iDg!�B*[P
"P�;�:����,ʙ$���Fyt!4�����i<��e,.M�o��/��~��r�X[[�����G�[lu�e��>�)�uN�T\H��K�g�ł�I�jQ�Į.��J�V7�ʐ"M��.V���5����E��T̢��uz)8�5�\�:u�h
�h
�LA` lx�ؓ���X$m���� 	f��Jfd�?� �B\#��<JH�}(;eqAA͠����lh�0�X(��.�	���l�T
�<�4��~�$USh��h����f�ň*���A��"�J*V:Q9{z໿���/��_�����������k7�w>����7�{� �ۗ�d��F���Z���K�����
���V%A�ZA-�����1�O����z�|pY�0	b����Bp����*RU7t�L�-ՙ�V�pCfQP��T"�<f&��*���"[�]��Zb(��#V����V�$���F9L�R�a�������)z�=�}�{/�m.$�	�cW:¼��!O���Ȋ��th��e��+����5;x�q�dL�[oq2p$��t<�ӧ�
?z|(�=�f�7�dC�k��O��|_��+��t�- �����ŪB�4Fm��E��9�P�n+tf� ���W��Ƒ��Gvo��`,3�QˋBHRJ�#%sWכE�*��B�
��"�'M�hDI0(�`
���'����{�v����׶��(AaA�ng!�s��	>�W��lI������1:�%�DL���k��D�x�v����b/�:����
v����-��o������?zmmGR��:��ZD(CD�;;�`��rVyD6��J��-����m9�w�����/_�<�
|��N� `S2>j51�����>;e�,~�0iع�a��]����I1]E)�8���Vgg��z�A��A
���=�����B4V)]-N7G�f	¡.��9n�,���`h�W������Ww�eP�Q-��t�ҙq	m�%��N���R������E*[�YܹsK����g'a��Q"ݨ�����]�d�0��ij��p�2v�րD<��_����}<���q�ҘPe��h K�������m.���#%yɨ�KV�E���<D'���@ ��:�{�U=U7���w0�
UȂ@��}�C��@{���>tm^+��,*�(�=����]	yc�\w�ڼvx\1�%3|��?�<N\i�%�& {<nDq��[Hg2���v1C���u��+eb�Rv�I�gC+�L��R��AIc@�N��^:��r�}��Rr\TSC��[�!Upl/�f�|D�m5I ���B�ݝ835��6*U�sK2���L���Hˋ[��
F���)\�8�j1#��a:ID
���#�oB*�{Bpz��;(�7�aznV�GI�.��:0�B�\���o`anW.���+��o3`�(�������Gk���N<r�,F�0�E�P��ۋ�7��BQ�ݭ�15��:��;E���:����L�=���g�S����.^��=��`q��	C�Y��j2j6���PEСt�\U�mJ/�V֜Έ_C���K��\?[�bYc�{i�]t*���D�QD61������l����o�87-�7�Â������<+SȽ�m!F�u�KQ�ͯ=�o~�9F�H^
'g(���`��Ѧ��(�c��E�j#�R9��(W�"/b�D��Liw�#��mv��֩R��\:�t.+ZN�x��l)�E��ei25s�ҳ�6fi��/��v�����Af5�OI:bfK*���~[0,^��I�LR&l,4\�v�O�C[�����R09\�{�(q
]*Jދ�₁���Bz85�:Ӝ\�w����;��T�T M�Fh��orzb6k�g>�g��8L&�������^�gϞ����oݺ���m��FY����3OC�xj5)�ш���b�Tr
Y�����h��	`���*���M�5�o*�÷�h�b��},6;>��O����������q�<�@Y�X�Iם�kz&ut����w �T[�*8M�0U(S6$T+�\d���U�u$�Uk�˂���JQ�/Q�֔?6����ڬf���bq� B�
sQ�]0�R&�,�����K���5+�����]�xz�_��G������_�	����o���?|镟�nW�;�?��.���umE���F-IBF���Auf!�?�ۿ�ݹ�zrq#�VϪ�\������)�>QBE�.3lF�L��&��r*��f��_\ז����5{D��a�1��x�[�)j�U��Єh
Ѣ�����\d�3o�݀�܀��A%�D�z6���6㸹�R'(�+#�ʕ�Ǉ���?rUzG�QI�<8�9����s;]rCw��ho6x���C/1���[���S�&1f~���!��p�^O�H?�#����[�R����;���}F�Ͻ��~� ��:��6h�6a�k�F��HI�	J�y%���*�%ͯ��8^[G��R
Z#�P/*S�,zvKh|e�TbJ�?r@�y7����3��'�q�-�`�9����u\���LǱyp �_\�X0�`�j���jM��En��m���h,�mi�TL�����Sc��d��ູ�����*�����!�`h�v��\��{�g;��6���q���A/R�V7�<��L2'�d�M�����R�<f斱��-�`��W��I� ��"��B�o:]ƭ;��ߏK�/M�j�T�7r�d����b�I�ª�Iijt�~�,<�᰻ϰ���}��Č���@�H����E��$���삄Z1���jW��#��=�2E�X���:��lf=�V:;���a4YqtR���l��\��&�i�c���� 5�Q��:,67�&;���O?��҂L�Μm�ӤG�@a5{pp�5�<l��e��m�X�H�H�r⃠��ܙ�x���ʛ�&Wjh����[�V��`w�E�٨En�1�݁n&?[,Xߎ����eN!y�� `WQi�Q��f�(hQw\H�M��y� x�b�!��);��+{2Y����v��S���;rȠƛ�~��F� ����BowX%�k��=LOO�362���>�,fdry9<��!��bA&���0����H�[�����&re�j����H��>I9on�Lu���:��	�b�����W>����}��.�r�����`t�S�2rt,����Q�K�����	��\N���K��j�?�0���6��pȮ�Ղg�q���D�u}�oϊƟ��6�������ۘ�]��_��3�p8���?ĵ�K8��?)�4ϝ��hlNr�
�Ϭ���M�z1$��g47� ���1:��ޅ����It�t��ˉ��!Y%5���2U��|r+�6E��Z��$1�A�D3���;�U��L��v+(���Jk/��$�whI�Z�M�`�Ȃ�P���|<�Í%�|���p������/cei�*Se�R|���᳟�ut}�\�>���Ǘ���x�/�R��fq��')P/t^/���@�PC���-�ǒ�c%���B))��	�|N�T�ʪ9�?����B��N�]���ڞǱ�����=�$��e��7[��{��؆�뤃��TB*)u͚� 6�ZqU�zS�i��}�tz=�̽g���y%x���9u�4�F"��L�b�HeJ��%Y�Z�g����=3�x�g=���Y{�Y^[�d+Ӗ�I"���9�����+�{�[Mj���>2@�@}�y��>7(À��ް�����"���>�Cw�����]�[K�����0B�n9;qh����I_�t�d
ET�I��H�-▜i�%��Ev�Pg��l:�ٙ=���2�n�~�q|�����������}�oq��x�<��#�+s ��_��=�����j�C��hD[[)��c�&d��JFw�f@��8�D`m===j�ٔ�k�r@�Q��h(�xW��n'������!���ɟ����u8�����0T4�y8]ģݰ���3��@9c �����܋�����&Zn6Q�57 ҽXw��M*�1���S����a/�ͳ�m����Y �T�p:���E�� �����B&����6k����������~����+����W��/��dOO_���1���,�b$����|r����0����~~���~�c���5K%�i�����G0P��{,!���ڍ}f�aӆ��?�ƏN�"ߌ���Q�rY��@���c�ȁ��a�����$������[WP��
4�p{���Tء-+����� P����_"&b����|���7ɼr�._�(�y�:tHɡ\�QXu��u���!�s�^��'Q��H��)���b7���oL����gPT�ŅU���/�^�=]�����V1q��]HW�����8qa�fMG@I�\w�A�J�~��G�.ā��5�F��4�������^��*��*)���+�Pg,D�p7�Bt�C�Tu(�����j���u�����|��M�n�p{{.˥�����:}Лj�Llz�(��^��%	(�(��ɉQ�19:�e
-��L+lf�~E.��IG��e�(�S�X_I!����F,Ew��K���i��XҰB~�މЄ��)���e����X\�Do��hD��U�� ]�� ��
�g���.�Q�
�d��9�����ԋFE�̲5�%1�ׅɽcHp -�Q(��l[Jt����ښ�Kr|)���o<A<bCn���[�<u��|�iS��ͬ?��� ���� =�!�u~vV+eRz��r�@4֭��ͭ��؋�I��5�������p�A���~�h;76����8{���$����=Qwd��\��v�g����t(F�J!�����P��ԥ��    IDAT�".\��F�mO�!��R�p��N��x/��"�P4��߇6]��y�%����>�7�p�z�������n�Q�����@B�:��]��5_���	h=H7����x���0���"�t����,�]����I�=	�\���hWZ�N���������76>���<������`6�W�_�߿o����21�M���\����T^�\���5�?(�{img/^�Z*W�[�R6��BI��Dm
g$}��6$��m������-�ncz�B8~�(zb����`�h0ҳ����˗n ��*(��;����VtI�F�"ޟ�N^E�X��@�^��@O<~Ɔz�.u��.�XB6[U�Z<�+XODT����q����u���.�l"�S��r�V�{Y��ab�OM'�6צq���U�PW'�����㇆p`l6�O�R-�z00H�P���M�=?�KW�Q���%�E�l���:�6�bQ��P�,��~mI'��kͷJ������4���D)���	�R�=���4[o��A��C&���D��k@ju��ۿƭ��$���@����>����S�
f
5��ӧ_�_��gq��s�g�j��?�#[�9@51���ӯ^�F�Y0nx=!8�zx=k�eS(��p;�yD>�D)G�a�M9�0|��/�xw�xH��NjG��V��p�u"C<�M�ep 0�mY�*K��5Qg�N3��;TY��KW��q
Zmpz,�<�����p�-!�K���M�+���Ľ>���I�g�VS�ź�Ʊ�/!O��liR/�_(jʦ�4�-�u�v��g��:�*�Z�
gQ���N:$ϧ�߉�H��;�����u�z��n��FrE� 0�.��]2q��?Ӱ�ׇ[ѣ�F(̾G���:��c�<��ZjB�s���N�YI���ӫ�t��[itw�*M�ߛ!^��G���-
-���/��7�'Aq�Ep��>����S2��I��h@�ٱ�5��"����6�/���rڊ��6��xݰ3 ��b���\����׭j���<lt2�h�������j7�-�?�R�t�+���^D�T�%��-"�8�����~�����#����ۉ��w_�ݓg�}4�ɹ����3��r��j�;����so}�ņ�s( ���ƈ��(A>�����"�nk����X n� ��SV\Tx'I��5���
���� Z��d1�wqXmco]����
[ȯ�!�x($a�Kh�v��n�艛޴�p;=j��V�<ٿ��;��w>�ׅK������Z��cPR�|x#�^���������؁��~�����K�p Nוjx�W�rF�	��8�Ο��WO����Ao�~7: /���E\�v��O��}蛸���Ó7��mC�]B�~�Ssj���"y��j� �c)9ֈ�-�63�,. u�l�lV����a���S\��	���|���6�<�_��]�6P����y�)<��7!g�!�͊�D�r��/�B���ؒrD.)� ��Jt'��g�I�#��g���vV����ml�A@M�{��04@���
A��8��kH��R��\6�Ю�+)Ģ]x�{e��r�ĉ$�u���8}YN�����\w�=6�2�P�L�е���L��Z��m��l�X<���@���R���n����`&�	�(W�*�m!�����u�9m����QD�^=N�5�SM���a#��p<w���,�FI����z�܏ѱnafܪ���q��YT�y����	!J&(Ё��y!���iTh+�h*h�.8{G���A��Ѵv�D�I�KXXY�{�ky��c�^�R�v&�����ߞ��h˥4�JQ��{��&���ifLcn�&�8�#�� ��(��6��/\��&R��&�~����]�`l8:��X ^���ڦ(k�&7mD�88��@"��ݦ��
7�:�E�C�({���#�t�J�����R����좾�'�]wLbl�K�[��qkx����57��sh�t|o�b��ƍ��?����`/|�ׅJM6��bYu��rR�(��V���N�+�8sᒆg��#kD�	��^7�����9���Ǡ�M8�}�( �C�G^v�HP(�����B�s��eKG��h��aC<����7�Z9'�ǥ�^>u��,Bј�Rz{|x��{d{��2�n3�I���&pp�}GН��h�G����~�����8q��R55�>r��4+�ƾ=���f��@6_�����+�p��RQ�ۣ�1<tl{GGD�=w~�n�"����qƵ9d��/�����Q�Y�CWo�¦2�i]{�]�:r[G�]&g"���*"��d�ßلh�����lmwàJL-��͹뺢���E�JE؈�g����~�7V��/�=��\T�
C��N�t5�7?������p�t��E���N�:%k�;����<���142 ���8�?���*�Z8և��q���{��Z���2�����H�,"u{�lA9�x�ۅp,����OC�D4���i�1�v�q��9log:�u�Ă@��l���['|S��5���1PM&��^����SO=���_�<i�D�S���[��d�'��"��I�TZH���hkR�<��3y��I0���d_.MEΖ�\Hsd6C��A��C��f�k�Wݸ�h�_{�웟�G?�~�<_�.�/��g�x��������S�>���
��2��5�Ͱǃ�VRtY�����l�	<��F#бk&�N��i�܀�Ռ������+{ፔ(�|��x�;ގ������(�����_����m��A�҄V��-���]0i��9U=j��J���zE�0Jcv0@���4��yP��
��N0�du�ef�D6��>�'�����A��:�c2���Z>B�(�A�h���L!�\m$���?��w����ѷ�z�����տ:���ݟ��������~_0���^��P�Յ��ho�y�3x�[ߊ��<ʥF{�34�[b~��A���YY@F���"���6��j�M�n46rm|�{W��Ssȷ�+b<��v8I͇�^v!GN���R�b���毢���yX�,*�-�]o:/��^x=Ax��b3�z��F������W��.������ܹӸ>u�}�Eww�^ ���B�7����`�_�V�D�U�hH������իZ�ix�<��x7���pkj���?��Y5j��l�(�V�ڠ���=�$���u�����ZB�ݥ<��(T��:�$�2�:�����gs�wB1����-dgo�4��'h#�iӋP�5�����ɼ4S�[��p��K��Z�jjM����	<��gPt:���%j���Bn�\��\�́&��d�H�Մ�n���X+��;��{F����P��v*-n;�L���\�� �ph�]�t����+��p�ޯ�(!��]kqa�J[[fM0/� 	��:y���XD�����h7Q,1�����&p�=��XH��{����I��N~���r���N�6E�iS̀02���016��_"��o&Ӣ���Cg��^L�	]��ɛB���������v�K���*�\���r~ G�2��E��Kl��Q��\A���P\K�\݆��\�2�d�M�.?��
�a�L���䰐5�p!�����<���P,�g���{]	�~Ձ|���[K8u���Q(�ĩ����kҨ������w߁@4�r��d&���.�Q���D�;(�Â�$/,mjېɖ��e���p/&�a��K�Ϭ��fM�0��6�
��"Q�<�MLGk+WsИ3��sT��)z�|x��1�X�*ĭT�a�����2f����w�ȁq�����VW�nh����`?�;&��k��k׮��;44�=�#���_"E͉��$�g�4X����O���E�C���\�����*����,��x=��l���a���(A�]-E�&��&�Z��RgF�grb}�~���\˫�������sX^I*o��s��6-�����Ǿ�.�v�)!R���s7q��e�*5x��(9ǎ����	Y^�v���D&߀�t"r�ر}���xS��6�?�M���2^�x�iz��Ն�����D?17��6SILݜ�����̰�zƼ��}�=pH|����8��}�^���~PGK��ӧ/�,Lgk�хb]�����o�>L:�H����5�t��u6D�e��GOY�h[�7�͗��\ǎS����ȟ��}�@�Mn��Gi'���^|�����<���/b��%8��/�@_[����!��η�矇?D;�Y�ɟ�	~�������?�>��_���Q��n�Z�����g�.�A��o\9�pH��bn����]j�m��`�5�T,�dO��:�Gy;I����P�?�0ڰv{s��k�JPH�&�,�x�S�L�A�����Q�t�����=�U�E�Y�a��c���G�'#�/_�j��m��!��.4�����t#۰�n��nwJT�PZ�6ɴ���G�ڒ�5tol�2�<j|�D�#틉��D���t�6�Q��7=�$>�������ʑK�ۋK���?���T?X�
�|����@�S��}�����\��w��x4���th2!��\��	��>��-���\��Z{�!��B.'-��������'?�w?�<X�����������7EO�f��zZ�2�M��S:!�d3�yM��h�2�/��75[.[�R᠖�XLS�
 ԕ@��B��_�h�n Q�>ޓJ.�6�Zj��/t,�5P��-3��3�nn\<H���khW����﻿�k��O��{���&��������7������@0��L$�?��֜��pW��g��'��۟|�z�s�_\���&�Gp��a�u��Z;#���z��XX\Ǟ=c���?���(�U�w]�RT��@��.e�����ʋY~�mx�6��<R~oa��e���^����V9P��K*Y�[y
����^*��Z��h?���7�]Ͽ{���t��[��IhP�8��2׋\I���,��~m@�"�jŗ��DpY r��Iѫ�hc`hccc��@ţ	�ܚ����7���¼�
l@�^�������4��w?|/�V*�·N��g�a����MN���E�T�aw����đʲ����ԗ��6���;s0��!����1��ա!���S��2�����������X�������oG+��JjC�aD��
x��o��ͯ��dK��v��.8h2�Hģrja�o�Q�����P�\���RPdY������~L��cRu�v��Ҿ�nT�%%�nl$e�7<8"�(����ؠ�)lm�!vhg"l��r%��D��H ��N�̙��Je	3�,&t����äu�N��6��Riz���CW<��Z�Q,ױ��.�I����p7��5a=�X������ȭGE:B�7 t}'�|�".\�!k־ބ��D����f�3���P.�������˘����Ӌ��=7��d�����w�]G'	�P��D�)�m��1���i-80��ѻ@vO>[�փn_3k8u�2R&�a&~R�W���n���{�����
6w�q��i�����O`�Đ�*��PJ&�
e�������]�����@�V�m|�(�73�xe�Ԏjt!/U�v6]~C�ik � K.2��N/�K��6�{BxӓiPͥ�u��Mk�n-�)C����"%l@��?e�5��|^sn�Ƨփ����k�%�<t��z��c�kۆZӆ��g�깋������탃	Nw;������]���ƫ�a5Y�7�v�RW�E�|)6�y��)�d6`�-D��%&Ո��ha�� &'��u��3��&c ���v3s���Y֦�nN2ܾ�t��<��1���fn��{y��2^=Y��dDp`��;*�Kn�+��}4��s ��7V{z��V��}�(?�����X�d _\�U.���Pw݋����S]o)���kHgKJ&hsםq�~�cy9���^���SBF�x�A<����������n�7��G�f6P�z	��_6������m�� /�x3s˰��p�ʭ'���-V�"�1�P:5�u~)�6μ�fKN
z�b~��B��M���|�]<�/��H�^��IAk)����P��:�_��G��U�ş�ٟ��?�#!|��ǯ~���~��k�26�r���	/~�%Tm����vp�J����KX-��$����P�g���D���l�#��H�v�{��rH��n����0uc��9�&QS�|n
����b�/�лH����(<�����٨�I�^���>�F��^n��dm���k�1���b���
���|�י�K�%iA6�M5��;B�I�蔛S����Ԩ��a(�5�<S��|k��crRx�r`A9�GhC��c� �w�-�Z��~�3�5�I�H%�3���T��D��h�X$�I{�.^�$@����PD�����M��O���_��t#�B�p���{��f�.�S�}7������m�|b�.��vL/��_�&~��SXZ�D�}˭?�	k��Zٸ0��h�`��M�=.�!�w�V��#
�V����:+D�����9Q�h=����8�N�ϫr�l���%��u�y�#���C5��)�7�46�Q¤3W�p�K�{z��[{��|��~94�|}�������ϗ�_���s���Ð�A�B9��c-�ް�>� ~��?�W�^����/�;2��{�|�7�����O����>�����������E���� ��5|���8yqC���=�i�t 
}5�ٍs�,N�9�=��(��}��먬ހ��Gu�▬_[�찹�j@�~��U
"����{�������O`gg?��06>���Gt6n�|N8-��3������Ŀ+��^�^ �TQ���lY8%����!�����ҩ4���q��9|���b.J���O�'�A�$�Q�\���N�s�x	k�.�{���օ7��N�p�!:T�+�9��:��!x�v�N/`��Z+K@qG�͢����5�֘�M9-[9�Q�-� �/�u$OOA3t$!oN�̎�!ҷ�����|V<�ō5����+\RČ�`�1a �ܸ!��(�#�1;-��=T���
��F�������<D1�~P��`h�mn(l�l�ȑ���R��O�6�� J��g�nd�FjQ�Z͎<�|���l�K�*z���g|X�f~n�+�2�pr �������^bA�1ͻ�&�⽠�'���~kb}3%�W�}]���&%&�!pq뎭�,�;;�Ts(FcHm�p��nͮ�VnH((B_�ī�A��)�u:k���@*����T2'�aҭ�m��j������8��<�yn��ҷf�1?�l�e{�q�Gd2���B�L{6kIܘ_B�L�W<����k�qdr?x�.���L�.gs�t�2�o,���w�}�N� A��I�W߬��'��沐)��āz����&�N�B�ڔ�;�	��ٴ�������19`;i���6Y�\�Ku�����D̃g�z�J��D�k�SXg@��2�9���`=�߅��9����q
�(kv7�����Ü��H8,������Lm�_J������_D>W���E7�٤\u�q��~�\7D�:{�f���D�X�p'���*�k��.��	�i8���9!{F�!��L'ക��9��r�)s�BJG�L�J�\I��멌�ݑ�c8zpng�4;f���p���^���������q��*^���r��e�h��`�������`����N.�l.�ͭ"V6Iwh#��"�����0��1�B��������qk�$l�`dϸ�����P��\�0���f��=��]xӳ�Kߔ��P�83�����dJ�,�v}ttPg����> [�Sy|�;�E:O�"�' ԕT<T��N���_�!|�#�7���t��U�P+6�-_�9[u���H_�:?�.�P    IDAT�~�#�76ej�ڴQ�U���ˢ;�#�<�g��D��_��N��7��c�>�}�=��Σ��R$ˀ��|�+���� W�����"9�y�lΫ%X�"��n����@,��XK�Bf֐��?�-1�E��?��t)}�v�?��+�|���!|���[&g��iOO=�1L�&ȗLn��3N�&߽ 7�?{�(b���a��^�{�|�ZI&����5,�na5U��V�%�[z��E`s�d+J��~���-�<�e��U)�Z,�U��Pŀl���{�8��'PoYE%���k�{�������@?��cʃz�嗱���A������ ����+!��\٫���3�"��C�B�����ζ�����{ �9�ŵ9d��s�m����0�N�����{	�T����Q��M�������~.��Z�K�� ��'~_�v�rڌ����M� '��~��sΨ�`��1����w%��Q�9˞�Xg����v����&��,�쌈��hol���S�e��q��l�A���;4�����ǟ8���Oz�+�Ք��~��O?��?z�ܕ\ސ�VZ�@�~0�]����COЋ���>�� *@տ�J���o}��x�0�������A_���p��p��x��''�w| --Q������' �/n��������(��
6�Ä�-�_�QQ�Z*b�L
��%dWn������7����{M7�+�B@�@�Y�K=D_c�x��o��� nޜ�ɓ/��s�G�r�of�r��-��CDkWX���O���k�1�#��ѿ�_��X?_�~�J��J�"�J�TË/��s�"_��f���O��h�9'�����?��|��QĆ���l"_k��l�ؐ�J�9�"����F��s+ظ1���2��-�*+��V��N�!g�#t�Φ�H%1��i�q���y�f�4}7���A�P w��a<���camղ��w�]hR��N�b���t jp�3��۩5;?!��Y�YX+�l�x��/�W �Qiuh����9)��=�Ji�AW�0���G��N�99����۝ύ��#6�M��ɳ�|n���ķ��Owcmø�8HW�n�m/y�y�$���T�X��m�����T�O�K_�RB|n;"A����GW��Z`}3�`�I�Do�n�w�PfwL��{���A�E8O�9mE�����N��n�l��8��*s�k7@,va�hFG�b�U�-�a3�#q&��:��#�\,�P��!���,R�Z��PKK�fn{�\ݱ &�C�p/�^���u����tQ�؃���`�ǏZHn$�2��	:���ΡTm!Shcfvs�B�v��T���f�%����5��g���/��yy�7Pi	���7܏��4f "^���6ֶ0���,��x��.�w�9a�B\���Ϲ\�$��cBї�VD%��E_O����ו�5�6s+��O�U��'t�Ir��8zd{����iy���
N�� ���I��W������U����ԁ�Y�W�Dw��Z\`�/�Ѿ(|�|�:~���z�&��e�ݩՑک��Ԝt&L�C���@r �-be}S�}���XDMb�X���4�M-cn!�'�:T-��t�1����H\I$�@�ʤ94P(���,c3��Q.�16ڇ����� ����k?��|Y����<^�~�����H%�8�A{fA�Ñ�{��wb�/�v��3l�%��L)l%71�w ��A$����b6]h�C+vB[mz������������^�~q P#$Ӹ�N�"U��tQa��6\6x)O��U�A�e���V��$%�D�}��5����б����8{�6Rk�;m:S�{�q����'h�������X�)#W���ۣz�-@){��������E^x������ɟ�~=;pW�y=礪�]N�/�!�������'����z�!b�������8�������	�	�\gϞũ������-���	��|�'q �=����VV��h8B���f�qaj	s�i���Pk�`�D��Ѧp��[u9�1혯+���ʨ�*�*��l�tg�Mܜ��$�M1�N���`�z�(=[,D"���BKE��V�Q�0ŭ��	g�Z��Β�yRd:[�g����3̲�\)/�^_o�1���q7�(^�p8�^h��TAn��K�����{�g���<nL�Ȍc+�G����P H@0uY�fLf�AӃ]g8�ln8@���;$X"�إW�5��Q��>?�pm�Dj+J}���Ѱ��.�(X�"���V:g�t� (�Nֈ慓�W'��t36Ԭ�Ԩ��@��Z~�v߱����������_����n���/|�o-��c��d`��/��Zi�Ǉ�Y�#��ޣ��wcs��p���#n��Μ�o����X�����z�.����<��#����p����i� �ZХd_��Y���*��n8�	�0��B����b� 	&ZLgm���+�H�L���r+l��m��2��Ku2vs��f1?�ч�Ǒ�	8�L����'���k�q��K����x"/&Zh��vP\���*��(�]z������HS_���T��y�'�I5���I��H��f��r�h<y�Q\�>����{�ɦ�q���p� �==�)�-�_�G���M�M<��}�"�/#S��4W��K�G��`$�&���/>��W7�5;���2��-�m�Z���&���6=��QR�)�����2�0q]�F���rb0�	�Pg�ឧÓ�y;	��꒸�D�����kȤ���7 �NY�����e&]r�jԘ�Lv���:$���*�3��5�mU��&Փ��27Pe�!��i�h�}�+�+B����f����B�m��h��fɤ7�Yc�E�^C�0(L�"B���{��w2��K*�����s�"b��˴a�
�;�؝�)>�a]�f�J����I�Z*k������N�|m��R�����l^x�bQ���N_k�ܓ2���%�{/+�O�t�X[W"�%���VY��@~���ִUQH�eC$D�}��Hܶ(`��@��NrD�����?��3���>��w#�P.`c}���L^V�]]a�yd��p���mm�=	��.�U���!��"��bqy�TҸ�9��QP��]~��zw S�C��C�`[ݴʅJ�z.w����c���u%_�b�v�k�_e-`C��_"��`o�6W<p�g�`�;@ʗ������"������ � ��RS�76��-�<������{�g�^0ɕ����^�����L��L�zG�ʍ�|� m:�d�!1���u�h%���WNS�X���k����-T+�a�h��F�	:_z�R��05���W��;�G|~��B0��V����Ts���(�������XZނ�lؙ��B$�ơ�Q%io%ױ���p,��#����2�V2��Ӯbh0��;�����Ŭ���V)�-V��GW'�~+�*��(�׷e��͕�pǢA��q��^nx膢���d��P*d�z�?��&7Wlcfq	/�zk�����YM^$nI��A�U+L���^@�䡓�{�瘎F��t�0��(�שp��D��[W�\Y@3�S" ���ZNju{meh}#[IwЍ�l�>��;�	���[�/�L��KI̯�1�̠��A�%�	�c�!�Q�P,���~7Z]
S������.T[����%`ǆSvʤ���X[��O^:���$R[e%�a�888�'�x��{16ҫ��g7��O��������kS=�ΒU�-��t����)���b1��w�_Amd@\���W�^���6R��V N?7~��qC@�n�^4�#��X.)GÀ�&Ԋ��ͧ��x���W ��B�\@�L�h�AQ4s�8��>F�s�r�KL屔�:�Xw	n�� ݔ���q���S_@=j$y��O���h��۲�m�ͽ�����{�s�����uN.��,����$���A�Dp�l	���8f��+�~��-cC�m���͊��#~?n�M�Bj?�՘���b+�G���9�"���S�РYs����F)���Ђ_�
Y;�?6Nf`� ��ِ���/��6-�
ET2��C���o|�O�_���O_��W���5Xo׻��g�K�#U	:)<��S+�=$�E�O��L|:���O�~���r�ȇ>�'yS�oaui�Lbt0{�U�D;�h;�Yv���/�<~zzt���2�l@-�%�DN����*��א���Vf	�m�MXm���̖��' G#>� ��x�s����8vҫ�3>"����D��M]�׾�Uy�9���;1�a��������ߟ(FMr'��}�eH�c�U*�c����N�}}��Ў�bjH-��7�
�a�����(,�c
���pvs6���/?�o�'�5B�s�m;�ng�HWj���E[�5�ǡu'����J��mV�к��Zf6aw��p�Ԩ��Lb&m�F˳zYu�8u0�e��v��@ECA0m4�.�=���7��?�fЇ��E�km]gڟq+�3D�h1���A�P� �P���
��z5i 5�4�D�,"W�7u�(oVԼl'R�;ऋQ3��L�r�0vkL�&�����!�=!!��@���^�;L��u��7�PI��������Xx�/�ntDO���x������Y`��	#� [6knԊt/�y^t<�Ӽfk�B��b��Yr��,,�m-x�Ɖ�F��dRAd3h�/�b��1;E]����I)����
lV���j�x ���j�!���7:�4��*��pR�h)�k���.^�L��h��9��rsXmT�`F�hT((��I������R~��	$m�jHe��U���o��g�a"����^�,��?@���il`�3gǕ'[$Ռs�]�t�^�5�M��t	�2��|��۸uh��q�Н�I���8^�
��
E,.�J�GKaZ?�U�@!���t���9��g��0R�:����׭!����R	3���d��8�#��46����wŨS�� ��z��f�)�}4�qYmD��7.�N4h l�j��d���^9berUl�1���7gQ�T0�Ӆ�xD�!��EC�̌�G5�)�Rm`}-�3� �� ��{�G����@G3�!��X\Z���w�aye7o-K�K�[6<3Ba�R��"��J�&��Z_�6`��c�#�S��joI�ᯧ�U����	�Æ�ϩ�� 7w1�D�1Zs��/���o~�P���,.ߘ���m��L5i��wM�(Չ7��-{�1)�ry3����x=�X���T����DnZ�
An��X�v	s���/NnS�dicy�Y�Y��J7`sS�܂3��k��12:��DP�(u�z=���w�+���:���u�`�I�mV��0��`�w��z6��!��DTr�piyl��E�k�PN�Oבc��^>qFt=f�x`�!2}��A|���3oz� �qF�ŕ-����>�������@( F`��Rt�����YR������?D_����n��秮azn�\[��nf,9�ږ)j�Q���&��5��� ��9�4�S�M�#Kpi��S�)q��B�ZJ��'�8c*ěgX�[���5
�,��JTB�͎���Iu�؋s3���@q�<P���6z@1wx��}���P:�W��������69�8q��/`C�n#������G�7�u{F��j�ag�Hg
�����c�����6C�J%̜7�c��GgY�X����v���r���I&��E��Yd��h�+^v�5��$UAz�I{�7��a�w�������+���/|��G-����W��_M�ι��������~�W�w��n�o�^�ỳʜ%�;�x���]^v��t��o��G�_������~O=�4nL�b��6NNb�;[���@��U��߹���ZD��M�V�+���_n���e��ن�U����M�G+�4v�ZR��@&I�;r��FF�����h?y�>L�F��#[C��BA�|��������:no�i���C18:�r�,J׊���6��BO�KBTL�4��|�on`ff���G#r�����Ӳ�V�b>؁W�| �+'\4�,.n�o?�u|�K�Az�Gl��߈�G�V��T���ݍ��|`U
�k�E䆺6���D���$��MԶn��(���3���ǀ�z����(p�Yxz:I	�ߓNmrR���łU�6`�r�q��O�M�{���Kj���*$�ݮ��:t8���jX�x�4J~
�ZfJo�a�:a��zE���T�wRW):֦�n8���w 
�$&b��v��Y*�B�<Gn�ZlX��_ϯ1V��Y� �˦IJT�,�\%����n�D���i�P��q�s�p�<�mt�J��˫À�{�R�B��1"͖�x�~"k~Q��BA��D�ZE��EU���ϯ?�AhDZ,�lɝwj-��dLׇ��||�E찷̪���(7Eh�ժ6JmiF*rKQ��2�U�&Y|�����d3p���U�X�א����9�M蹩7�`��磍6�U�Ɖɢ
b���B�I+MRY�;F�BX[Ru2.#v}f�C3�Q�F6\^xv�5�+n	��:A�tk7��V��&��IT,Qd���EUj�$(G#���k[���g2�|�����E�g���68�"��=B���m�'��"ڤ�x��0Pò�X*#S�+���ݯx�����g���>_r�0����lH���)��C� 72lH����E_ODw���9%�,�+�ftd�bA�ӵ�4�r�g�Ъ6v��w:���qە	����i�8ئ6�)�{�G��`����{G0������Ï�+N��˳�zm�2�E]�=��0�߭3�i��'��z��L+�:�-c'K�Y~L�|��1u�T���,lm�ò�q��9=�Px�.�B��ظ�?���+k�q��y�n�����%��ѥ��m�I�@��n�#�Ƥ��>t�a:b��|�)&	�`��
8�5�x��Ν�;��Ӏ��7�1�m��`  ����S��q�ȱ�8txJ�4�\:���)T
ED���=�,\�\]X����W/WЮVp�1��a�`�LsE�^���U�M}n���qQg]f�m8���VB<]�fn-�qS�N
A$����}�}����0عn++I���~���3��,SK��r�Y��J��ݥA���
��Ό%�ު#�#�7�`�S�p��"6�*h�T9����J�(�kT`�Ƴ��@@���&6��"\kw[�K��x��1�e.�Z� z7��|F��`4�Dw���*�T8�*W�j-Ke�:f[��,tB֜���'f�o��tHst�	x1\Qr+�\���_˚Đ9�6�����i��H�����nMϨO(�j:�<W�uB�.�N�S[{��U�F[���Z���?\.c-4k��94���n4}n�A�xF�W��@A�E�#Чs#���B՝�(��A��5���P�v�&)I��<�t�&��I�|��W�#���/e�'.�|�o����|�g<L��p���8����jՄ�G���n�B�mo;_�7���?�c����C��qu���i$p�V�*��:���\������������R#���:Ƥ`6z��rp�ۤB��]Ϣ�8�����,�4PM�Ɣe��J��zʂ/�������h&XN�+@"���ذ�9ZԘ��B�V��3����-{������w��p�\&��Ԗ�2�A��.ٌ���t��/vv~���oZ�q���׃�?���, B�Y(,�q�^G,�%���SW���w��]�71�����0z�>4=>��
�9ikW����r�hK(JS"���ml/o������;��rp8���e�UF��`%6Z�]�+1�D��v�In��ņ���@�oN�    IDATR�u\�����O����U��V�^��X�a�6C��΀ m��5:v��\c���47h�b
��vJ�m��,�?iPoٴyb�Cx��q͆��(A6�w]�,�a�,0��D:X4i5� �&'jU����f��@���RY�H�O��]h6�,~-	vW��E�r�,Sϻ�&�M��	�H�`�%�+�6�w�:Xi�tآUi�	.�W�|�=����A�)Ho6��v������q��z�Ɔ���_�o3)Sl}y��_�kb��af�6��č2�hK4�b�(zj� ��ф4p���U� ��\�;N�����ψ~�lN��+�h�b[K���7��9�0>��$��g6E�I�5��y�8-�I�$����8#��jD���2[Z���9��1��ְ#_����`�*]��6�k~��j�"��y����J���߯AA�.^�z�r�FQ�:��k[B~���/��CJ�.��&�6��6\�rx�@/ݐ�@��L�(��,j`0��Kg�B'�f�Ϻ�h��,"n��+W�re�}�AN�0W��2G���I�i�Yu�ٲc��F	M[	� i	�*^W�[��H��ȃ�r��kܠJ٬��^ZT�]B\�Ɔ�����i�}f��*e��Dġ�TEh�=�FW�p@�n�]���3�Ц6H���a�͵����ŜU*EZϖ06�/KUr���5_*cyeM��`0�B����-QR}�(jM��tt9"4BJ�?��[t|k�Ɓ��4�Kb�=B"S?w������^�J��x �w!����ԙ�@>/�e��h���.p�X��y��Y��|	tE��±{���� f����+/!���&�{	������p�GaE�J_�Vr�Cɀў�����u�^-��M	�%�,�I{G�x���n��G�lD�NRR"qm����(t�����E+8��4Eܿ���xX�#�(u��yQ����e���Е� !�;�@w"����d��>o��eYX.�Q��r���2.^���z嚅Z�^�BżhUT���0�̨)����;�x��kYq��ɦwMzM��Z	�JNR>I����ހɭ��p�Qk��=_(�J��f�<9 Q3�k�� YI��@�10YC�� �`.Z咝`��8|�Yb�	�n�
#t!�Q+���>,����ի�5=��	5n�&ưg�z�����2����|�-��Ѩ�����9�,�bs#���pL�'�I!�K�������I!��+}K��\�Z�rkM+�LN4qY�����@�{���I}g�䃽2|���r���C���'?�§?�˲!���_��/��_ͯ�?�?8lѕ���۱/�zȡ�+���cx��C��B�[Z���*��l�~z�,��?�S��?��O��c���)�5;t�]A��"4;�O�����VK�KgVQi�����s%�̓�֌D�y�y��'GGyե)l/]E)���@cۼ`z�8���n���HK����(�M��݇���#�:�m�%똎�sy�ng��J [�cemU4��|@Hav+�l6��%c,���(F��L�YJ�_1��٣Mە���r8�������G��*d%�Nb;��\� �Q(����:C�pq���?­���6Z�.Dz&1|�.��F���A�I'��u;�,n�ӹ��i�Ë+(������vnNg��[;�&�R�J����+�5��e'�������@@��r:�4�_��Yi��v��7�Q��ߍ�n$���(��Η�����w�9;�������p��i�,6�l�L,<z����T��9lwH�����P�<'0��;�|��L�RV�����F�5n*�>��#��a�T"ϝ�ݳ�Z�mZP� 0a)v��4��#����y����s��i
���KFg��aT������)%�2���69��Lm�W��;3��C���c܍Z���^��\�:\(�gl�+Q��ܶ���v��0�9D�% o�X��ckɖ�{.r�98)U8r�^�wD�uNK�q	��y�F�+or0�t""����Cz�^��8n$v7�&
Ղ]�L9�^8�GVj@sD"9ᯅ������n�L�5�	>����Qd�U}�X�h�D�Q���jǃ�8z�i����i�E����Aت1���F����6�L(U�h�׀8�k�v�DU"tD��.�Lf������!��T�����i.h��-�L���b#O��ZGp'���B��wJ�rMJ����RQXg#��;ͦ�N�\A����I^�C�W|>�D��"l�ꨁH?��冻懣�N�[�
�<l�<��d��MA���5]A�Z�;��p�PPXS�i	@"�c|���G�+17�(s�9:�>�cQXn�l�BNg�*��|n���Fw�����~:ƴ�(3���.�W�	n�8�r ��tP�YRs��W�oz� }/��~ؤ����`��j0�`&]�Z�Ӌ��d,�Mo�g��)�&����]�E�݆|����u!l51w�4��x	(� Q["���$���fsh�"táMu�X��½���K?Ņ�'P�fD��6���#�w=�f�>���ܼ�����(�6`k�4��}��v�zI!�����t2t
6T:��1Cg�H�����a�<�[Z����7�E���+�r��tI"@H�>��~�Em���VC������E�s��7���t?��X��;�v=����CQ�\\�Y���%$Se�Y\���H�0�A:�`eB�����hvx��~����ؖ�٨���F����'�}n����;�2;Y��e=[Dwӛ�ً%Rx���
[噳���-�V-,ҬS�8MQ3@ ����%7�d��`�N��|�]G"��A��:�[:@s�z%+�w�O�晠IoL`h�^�&f�N0��?��giӀ?lU��Nnca~Y���7�07=��[2�������`�Chv��̷H;�@��%�������ZC��� ���L�xS�����Td�m�8��̽g���y%xnΡo�΍ht@H0���D���9G�ؖgj�ry\�k��;ikf]����lY�i�G�hF�#� � rjt�����9�m��;��V�j6�����{��9�	�2j�d��[<�k_���<rl�b�f��>��)C��3��|�������ڱp$*����J+�K��ܔP�gob������qݾ}x�ݷ���/`[G7|�!̬n�����j���o���	�?�r���{���+��c�&jؽ�՚�8�X�l��ϝ��-����2H,dNX$�+�� ό���ud�Ϣ�:�Rq�n��q#*���6�p����O�����"8�o��~�����X�����1]H��{�SW���+.u<�5=�龲��.4�e'��Uc��Ӈ���h����i\�tQZ��;��*t��9�Ri�~�x�z�߉���}�ML�N"S̊c�k�^<�������W��o�E��ĥ�KX�,!�1�����ߵ�k�(�ߪx=�q�[����@HՈ�>�l`sa��e���&,����$,��UψSh�R>��J��`���=6���@r��rya�WW�}x�{�|�����X�o��&��(7�&Y�֌�X4��Z	"")A#_K�9Ц�0�Bn��)�6Qxn׽�W��xb1H�2qyh�M1�l�m�m�cG�Ĥ$��
U��;�∖�S����l,�b�V5�r�)��x(�v���f��87>6tq�:+�*pX���0�rG�|E;�����؜J��J�H�66�!�ֆ�x�bE�8���Q�16.��5ΐlp�FWA6�U���S�*Ő&�Z��ɻ�5�V��4���I&�B�⪐k�l��+��C���cA1_����k
����Lq�]�ʰ"���9��ōfQZe��|�|��4�D�����M�fe��{b���#�J��)p����4��9-�$�<� �r���Q4Ά�19��,���GĶA��F�<p�^,,�h�(��E��P���C�p$9�ֺq�b�J��/
�Y#D�X��.D�����x��a�q*Ģ��$w�礞�^m��5o�ې�GGV���kMp��L"nP��\]iz�~�F��Ԙ[�=��$o�M�"�(UI[(	$��E$��[�X�z�� m�-��)C�fe6b>�*����bC��Z��dl.7Cԣ ܸR��v
U�VXS�h�\B8ȵP�0�^�l���2���,=�� ʍ�l8e].	�6�pX�
	��z�t:��FgG��0&���_M����F�*�IM��z��*~;<ހ��,n�a���L��Y9l��ɹ��do�Ci-���rq�ܱZ��,,	>8��ٴԄ�G�V̜=�so��3z=.(t?�>b�WDL+�ȷTaWnM��7�~3��u�&/<�4N���N'�.�4Y�D
��N�v��=p�V�	�ؒ�@1{���ӂ�� ��|��SSF͍&t|f��Z�j���	(�<Mg����z�݃ٹ%����H&�؈�P*Uu-���L�m�N�āa��t
����X,Bw��=B>�@�R�Bf5J�bIgd0���:gE�w���cf~//bc#�l�*Z9�Y�jY�4e;j �9w��Z�
�d����9H@��ԞM�Z��C[ďѱ��M��Lk/��������6�cjf���&&�g�ɒ�Xo9/2T�L&��56�_��W��̳�˅�R��^>WMRB)Z6��,���d�hbN=��.�kX{�ո�]+�j��3�GGċ{'p���@��V�F�<#���J�+�{���4i���ڒ6��E� 9�U�\�1?������.NN���,6�>fw�B4��5�Ȭ5����.2ش1��P���&u>�4=�0Sy�8�u:�4KU4
%4s��ݟ��G����؎_��౧������m��.�>ah`���~j�A7vl���?�i\� ^{���駰w|_x�a�2�?�'J��׿����;o��b�����h�Ӎ݆�HHT�L��?�\݊�XO<}�^��;HF�#��t�����薽#/r%������PM���؄�����������(���r��d������=������0����)�C{[H���U<��c�x��P
���߽{�8��I~�f��"�Fy��v�ѩS����7h�Z����ܜFY�J�H�=X^\ҟ|�i��Y�؆��#����ϡ���fkǹ�s�xm.?zv�7ڇ�L�rN��(�mDG�L���9MՍU$f�Q�������4ʅu�����N:y�:R0�@���� V�[�9S�*���jy�ڔ<�q�I�R`��q��q�s�F���R|C��b��Vr&y���G�j?��`>����2%Z_�yP�}(��ߋ�<�iڬ=�Rc`UE�9}3����|K�*.x�Q��Q#�d�#�K��X2%+�d<�P�]E.�k��#�ފ�'%��� ��(?���H7�V�P�r���$��`'���M�/�/h8���P�,c�A�
��������"�����..5,&�r,
�],�(Tr*VH'	�]��������7V"�~�ȖST�%Q�Xܚ ��k��e�3�!ڣal��s�r�^w�R�v�܊��ʏ�ut��p"`�0��x�k��B&a�<l�d�H[3�,nYl��Lyp��X����'w�º��i��r̨J����4�+���2A��fW3�恮1�=mҌ�#���&��e@�y0R��p��_�$�^Ŗ����;b)�9a*j��� IcT�G�:*��������}U���>:�.cqע�m!�,@DH��;'U�ㄏ=\�YdQ�BC�|D��1H!jň�I�W�u�b���L��G�6��!ѕ��"e�k(i�K�]3�i�v��&ʜ*I�c��a��M6�'��ze�*h�L/���<5�p`�)bn:������E��k䔏�:<n�����FE͏�eqM��L�d�T@�φ�)%:�Ҩ� �����P�Q�c����rW+����*��Zʩ�IX5CN�x��vƿs�m�'K�?Y�3�ȼFi>���M�5i�e=�D��|�k�� ![!;0O��o �"BL>o�RpmQ[W�3&�9-���V|��|t�8���ہﾃ>�}d67�a*2D�!h�p��sp�)L^��ܵY�������V�P�~�aY��
�0��6F'��5�ϫYf3�t``��^�8�1��䏰��p9bX^K�g8�n	Lh��XkѬ�4��0atw�~��;5eތ�h�N�	���(�����/:���v1����_~�s ܨVL#+�H�V�l�9yf�X�*T�B�n��xր��b	��٬��#=x�+�G�p?�]<��{NڜA����;�هB[8��W��g�W8}�*��"�U� �L�āM{�&�����>�(B�6����x���155�}?m�Y�S�S�Ŧ������%���OE�]*��z�&NSz�E�pG����n��b`[7�C�,گL���27 � \��|�l��.?4����0&$�
�r��ӀK4G�Rm`ys�O|�+�K�03�kKkȗ������4�嵧s^!��l�j����,V+�1�MUz�޴�u隩�^>Ӆ
�X��{�>��_������� ��_{w�{?|��g׎qt��p��G�o�^��ʋ���{FC^��㋟�4��F���8�����7�,��'ψ}`�u��^8wQ��ޞ.�`Y��8uS�A��ՎLŊ�xO��$�?�
�g��͢��1���<9sx�ؚ��瑘:�Bl(��RO�Z��Ƅb�<�~X\�C���r�p٫���αA�㺃�ePF�T`#��?�����{߾}�.���Q�0y�gϞ��Ғ6鲜Nr:8����هP$��9���BcFFw�KNf�����8�<*y�����:�l�( J:5����$�;�P��p��<Ws�em�y ��A,r,Zm��Λ
v�-Ah�T���������֮^�a��c(���(�`�V����I�N�
2eS@>#|���������ٝ~��!X�D.j�:�8x�m���kB���4�2��q��P�8�_q��%^&��mQQ�lE/b��aB6.�Z����@�\�B^�;-ȉ����e�����.�A0d2�R1���H�_�#����Z�����s��P@��)�M<�$���\G�W�q	a�&LC���\)���(�Vvr���Q�d���G�qw�4��2��rLlv;e1�@&�6�܊HE����t7	n~|�`����;
`Ea���׉h��ɏ`X["�A6[�0�V��T��dS E�B��2�]�-�)`�i�>4ԃ�C��<u�����²��t�ry|:89Q�iLd<���9���œ���Z2͇����%rdj	�~�"B��ovg
)��zո��2z�I&N�Bj��l��~��tR�i�(�g�JjK��x��d1O�}u{�f�r�L�8�Y�h�D�`Y#��7�����D~m�3��SP�,�=�'���|���r���}��$]�UQNjV��)Sj�F��@�&=�6�6�(�I�r��r	e$��|�E"�L/ͫ�&���8Q�V�kgS��+*��Y(�n�F�E��Ċ��'��n�G�l�PG�()��hI��բM��.I�cXe�4�ݪe�`���,��`qu����Ph�#oQ
8=�c�K�X3m
["A,�f��:pϒ�d�p�4P�Z-K�
sY�f	�BM:t�Ot��{p�|��j.�)�-^Sԓ�%��J:8�!��HnO�G�Zw�iq��&����7#6�N���h�� �쁎m6��Q��x�Q��g>���o�A&z�oi8wO��TP#a�#��y�KY9�:�����{�B|}����~|J����û�`��7����s���g�ѬҶ�
G�.�WgЇ�#B��y�%�ϑ>E��k��A��AM�y��Fw!�މ�'N����rP8��Q��-/��o�I#2��A��A���ۇ�t�*d���l�U�X�    IDAT,5�SIsY��qO/�n*����ݳg.L�?|��^QC�Y�;��6W�o��������E��tr$2�j�Yd3Y�bG6We
��G���������܋/�{�{�1�
ػ��x�_GOw7.����w��#S&0T�3�i4����sa���*��������܅�x��������@'-<��8Q��?�گ90�A��MN�\�v�ȦXg0�)���'?��v+U��1����h,"�H!�+ɱ*���⒞��f�U'p
PB1o���'댎�vtwv�>�-2�]���
ɡ<_a.K+�q|t�2^z�L.��Ɲ�3u_
��<��ې{"�	�E5�;^k�EF��}�M4I�e�U�j�\/T���*����'��_��_�������ɹ�O��;�wl>u�}���?��x��p����}{��/<"�������\�����pߐ
�t����qJ:?��`&��١|#.���݁<�N�+I੿��~����G�D!R�����EE�i~�MAze��KȬ]E#?T��5
,M���5���0Fv����\�Z��طs�=]ؽs\�"�T��Sb�������D7��k�҉[���]�ũ -@ҿdB0�1���9=�>,^*�I��^�F,�D*�l&���^l�1�H(,i �r���Kk���.b��t'O]��F�C{P,�p��<fW2��#��G�;f7��R��-´F�҃P��F��k����֮^�3����C���r�!OI��F��Jcg�D��k�<�������"���ARH=� ^;:;��ϗ���q��[q�C��tc��2ż���t 6�QW�[��G�A������I3�_����J�߬!�K�Ҩ�A��u{��ak&~|;�f���4�GV�b��,Z%�S�K�|~�#�}8r�������b��E�%S�EK��Έ���"�U�c�����/T����K�&��� o��Q�&G�>�[�0d��������/�Qk�����/d5! M��hY���Ul�'��gu�8���3�J"g<dt�K���s[����v(�F�6�D��ȥ8jO�w�`\�(R����j<H�"�k�
�	`t;��{�t]����A�)�dpi1�^mp�_����+�Ӌ\�����@���ϠɊ�'oW��ƝJ(m�y�$�E1$�Ă��IS�RAN<�2���̉(����O�2-~*�<�#ѩ�1�/�Q��[bv>�*VC�QB��E�YR o:q��gC��
� ���
�f��3C�D�nO@��5�ԏ�X��DץF����ynMH��u�ف�5lN�b�����'B�*d�K�E>;�p���� �+R�v ����W�;(�e��3�7��-� �,������?߈�M!J���V�9���C��]j���;YgM��}S�,�8�<`%k2	�
�.���S2��e���k~��
�z!'_�#���6�M&��״��ϡJ�"��e�؝��������Ӏ[�Ϫ�J��u��m,b�I�]ᤌ,�Rh�`�B4fY wcN@T�4��܈�4q/�d��1?S�S�2	�a��J��5t<��-���q3!�Ur���\���:��]���i5V	�h���7�+_�2�G�ceisS׌�����`P^韛�V�XMbuae
�9ղ4�'��iG4�Go7�Z�o��*56n�[q6FL�us�hw�ޏ��D8Ԏ��/����'��A���f3(Pצ�+r�yQ���³��d>{����nVq*����%#��4�NƑJ%Dg�n���B��nGov�:���cx��	���8w���ܚi�7�#Q�Y��X�S���y>�_�9I���;A	j[��������O�{������.�	LMNcdhXxc���o~�w��Եu��w�/��:��!�������r����'���o��o⡇��:yu
�?�~��O�����
H�B`� ���F�N��STA����,��vR1����dp��~�s�����(�~����9	�I���
X]����<�ԸٜbeLO^C.�F�M<����z��M�������3'���]���AWO�r-BA꼀ٕ>8}Sk�<����F����=�C�S�ZD��7�B�N_@��|��L����=i����tG���R�l�r��?��~��?�2!��k�|���bjv���X?�����n�.������go�_Ѕ���?|���/邞8u���p��>i�.M"y�b�.i~f�͘
ː?�p8d6-�Uvَl���������<�M��L9���%Z�o6^Z�XRIc}�
+�Ȯ^E37g��FAM��Lv�6!o��{btl�l4S�l��w���;��o�W\/>�D|��?�>�~�i9r���g���@�N4F�YP��v,/t� >�<��������6�ql�cr:��6��]����)T2�ʢ�)�k��:X�����ꡠ�lza�ki�<LA,���E�/g�
�cp�u�l��z6�a�	��L��kޤ��Ө�+Ed7W����%���E!��F~h�d���EQ=�q[$R xh�3��J2��A���B�@;F�Ɛ�䱞�a�����A3��Z*�D~��F�Ƶ�F�vډѓ�v�䐷�:���3�����eiV�� ����ۺ����!�R��,,�����A��J;.��K��3E��*����6��8�Ѻ����!䜼X��!ξ\T�e�P��_[���S�[\� nK��Q*�lDT�ܒ�R� 赡+�C{ă��z���\F��$eڠ��:��2Ւ��j�&���D"��K
H�k����ʱ�#z!z�(R�J��kBkX8��k"g��p5�ť�������t�(��FG�'9ldrB~��r��uF�ķe��煿���� �pHD�5:���nHd��)���"���O��1t�X.�������p3�5���?Z�Y����iW��"W�b!/jC������!C����˽"
a-�@&[��a�r������	6�>$_ȠXN����}�ެp$otQ�r���;Ȥ[����I����fF��1��^"]����_HgQ(WP����>u{���c��|��(�OL����{�L����7�SK4ɕ�+Y�=FwG��K^N�H�Z^[��i+����PD:������A~���ɥƇ���%�'b�f��i*[HG1�����.� :�P<�&K���<�j$)$�)��h{��f��͍c|�m`J����uN��K���@�m����#]��߱�bR-'	nPc�Y�����!�T6�������+�GZO�����u��l��� 0�e,�I�C��sM���j�WT^G8���w��+�Q��������%ңx�
�
t��Q�����}A7f�|����$cJyeQbͦ&7�~N�(R���^_�^���~|���d�i�4�;��L���.�����<��	BU�O�P�q�[�-FI�ΥSp;���B��C&|�*�6��"J� ?�5dN�R���\^ �e��rhp�g�H�Rǵ��h�$,�ޑ�$�ͥ[�1����?f�  �M�����at��#�Ƶ�9,���G=���"ړ�����${6�f�e�S(��|J�ti�hSD��H�L��p�O�������c7�ǵ�%<�����[��ge�Ix�.|��_���܇d&�������g^@�lR6y/y��Z���Ƿ��-џ	�||�,^y�U���I���!Q�j�E1��f>Ӗ�֩�����(��pYq�-7��i�ph�4� �-Q��q��5����X�'�c�Oj�������Sѥ��#HG��O�*0�!
?oq�@�T(�؎q�ݿ;�G1�}7=��H
�&2�r�������ƻ'O����*���)A$�:����"��.��!��� h: �%�a���<m5�\�r�M���7������4��[������x�}w�k��#_��.V�3x�W1�4-�W.��!\���0~��q��g�"ab|��
��4�n��vb���,gg�C�ɀ�Ć�M��/�t��?x��dӨ�o��0�	#Í}6��6�f5����HΞGi�*P\j	Xjy�)�O�������oCãh��l��Ã���q��>Y�Tk<�{�<�ԓB�����q�]w��r��L�yZ��`'֊���%x�.���s�qmzR8�|@��6D;��nS�J��M���s��?�LGL���F����f��N���2���t�D�wD�!{0�z��J!�P9�a�H���ZB9�Bfi��e��)s� ��̎n�93wD���;��&�ո��Ł��<���&yJ���m�3��I�!8��{Py�J�t��DZA�؈N

9�F���ل�m�.l�}�7��r���:��c�PƷ�IQ.V�2ʦ���M[�g�i�B"ml��>أP��p�U6��ӂ�`9m�|��� ���0��뛅7��d�f��"�T�%�`��� �a\��dS9�������ͥƆ�fY�Y��{hy5l��5��5T��Mߘ3�H��Gg09��J���M�dl
��ӕ��kC���'�O�^�PF�֜��t���̦7�#�l��I̮��H���TJD��L�Ѩ�f,��EoWD�!����D@[�߬�ǑLet��E�n��ZL6��B����+W�v�W§�����o��(I��l5��2Fj��,w�:R�M���ub�	l��Ŋ�I.�D�L�Ħ�T�XX�D*A]	���>ن�!|�
�.���>��x��w�4V}�r�jV���h�&-����?�=+_�N�k
@K�p ۶��V�������d���̆�� ����O��F-��L�j����סtꚖ��tqJ![D�J0�=���c�{��}�=���'�X���
��һ��bc0���k3��}w8iqj�Nx� ����Ζ�g��n�Y�ժ��c��ƛ�S#��<z�;�w�n=��Gs/����{����̼x�ܛ��z!�O�A����l�+���bp��a �/�����fF��&�MR�H�2Ϲv�G�4��X4�V�<�R9�Ξ(���������z�-M��`T�ܴ#���3��nNh�c`#�h��2O0t'�$�VV+�2�v��RCZ��9�{�,�9h�*r(<1�iB!_��Q�ytx�� 6so=�4���}�36&+q^�D2�D6�d6�*�*�>�)P[��rA`���6�|�Ql@��]o�3��8wu
3KKX؈�V���р�#������C�y�pl���t3A��I��Y �ꑠ�t͖iVԿp
K=�^���5�Ɛ���v���i�F��JǴ֕�S΋ۿE��}3��Zg�W�1t�2璦.������{õF�	;R�A~�ڢ�ɜ�֪py��E&��TI{�CN�YDk�4��|�_���o(/cfn�����*�ں	P�'���ǿ��7�������?E1�9�]��S'��Rf��z�ȗƃ~J�6A�w�y�s3s�H��2i�T�&�7 ��WL��s����ͦ6��Xp�7���,����FM\S��YXF�a���><s�t�\�1
	���2���C�熇��\�xj)81cC���VJ�y�r4'ڦ�ɍ��g\�<��<v��s����=�Z�:p��)���W��VKe03;�B�, ����֜.x��#�<�q6�e6V�����ojʨ�!�q�S�����/��П�����>��o��o���g��GF����t(�7�w��ӅJx�������*�m���B*я�����~�$q��BXN/�V�כx��8~bu{|�m�e�jl���Dpt?�y(�*!�6��+��9�@2�٪�!P����^Hm�������(�"!;��f|���X�,�f]H���s�=��>������4&&&4�f�QM���-v{%���mzn��˺�]]�'cXY_�Ȕ{:G�p�@P�%rω�p��7��#��Ҧ288���D����`��q��5|t�
�WR��ic�7ڏ`�v$�Q��X3#�V�޲�d�B�b�BRL�\�A��5X�)4�����b185�iN�H$u ���䴽D���FOW�l8��
��v�>p7�-Q19�B�[�{E}�p#e��5u�-����{j���}����>�Hw� ��Awԋ�C���+��Z�"�-a~)�W�ˣA��,K��;(Yt�Q���(>�E:�0������Jj�Q(�j��3�.�Y��� �F(�/��o}�S����J����w�)lK�+{�q�]�HfrL"�����@&WF"�G�^C��!dVtE����b�k��]ũ��X������
H�F�o$��`o�Ý��A�i���|�|	M�hAghl y躉�Y��X	g�\��ʚ���GA����VB$�Ǝ�^�w" �C>�ս�F;��z�L�d��g��^N�X8�����|i����?��܊��.�_#Yyfۍ��P�-�9�`��D��a�d���&
٤���Fp�!�F����H}r;��;���^~���N�ås��������`�a�M6m���ׂ�;�q`�x<f9_��D�d�p=�~��3/#�䨼��GE�Â��^��9��n6i���07��ɹ⩢\`(����-{Bf9��o��㶠��c��6�
�����S��]A*�Ք��%����mlC1GCj��'݌NlQ8h�KD� R��6S�]XD2�E�\����<�gx<a8��36ׄ��l�1��eP�
R��D/�]�14 zD(�W�5*��Y��C���FK+�XYO�Mf�����$�q��}�/� �)94.YF�Λ�OQ�5NY����e�beQ�������|6�tbU�]�!��vhm��#�@,�����
N��67Ә�O�nʙ�nC�#���0��U�;\��H[ u������6~ �f�����D|#�x��	�^9�\�9���1s�}\y�5L����n�ݪI6i~�L
�l�TR�����_�LOg3X[_Q���m��;OR-�b1,s�V.#U(�zA?�R�,�h�lX<���s�!���|�hXI���CrVZv�O29��a��d+hR|}6N���T���DZi2,�9�k�rp�=Ғ9)���a�l[��n�8Q+�Sc,�Z�@|M| 辣` ��
U�.�*�Ղ�2֔�J��Ki�<��ሦ\l��q�I0cea��/�{���g����Y�W�.�?z	��>��T�k8v�]������ݓ?��x�mĖ��ޒWȓ�UCg>q��
n�e�ۍ�W'��K/���?D2������ݑ�sch�N�䖳�F,<W�����1�}׭8�{����*�����S�29����l�B��4��y��64 '3�iD�>�N5��s�!$�"����y.HA*$R�	B+���@)�Mt����#�3�7��#;�F��O/�puj���6�y�$66�� ��{� :-�I��X�4�0�٢����i��
��j�ݲ���ˏ��W��.��x��o�l��?y����{ꩿ�H�n���{�����3Vݖh�F~t�ld�s]��������[!��r���d�YoW=�n��F�wwh�Ǯ�/�Y�����vc9��x�)m����0���ǩ��R�\�*���&O����j�D�[[6Ov�OBW�d92ف������S�ނ�n�Ai���XX��w��x���dz��w�U�A,�����'���O�D�@�˫��������qÍ������5iH��%��[�ƴe/W�0���l:/����\ n�D$�"���F�̔��'05��d��� ވ��Ӌ�<��@����nm��m�R@|v��/ �H �/��iЫ��Y:J(��x	K�k���Q�Tatkp�`��T��ay�W�6�?v3n|��v�o,k�D��.N �#��+q���VS#b���5VXj�V~J�L=x��    IDAT�F��w3��۷��ÚJ6W���&>:}����PR:soW}�m��Vz��S#"9tC*PH��G��!��HA>+�H$���(z�"���J��$l����ά��W��F��`t �_�.YvG�Rmnv����}��R�Kk%֨��!�	�(�v�B�RF$l��۱o|ȰKn$��Ss�:����8<
���:��`�H/�yL!�*ԑ*�P��R�F�d�B��0������z:����X�eష)h���:Ρ�+�B{���ٳ�cC�����@KM�ኳYX�X�4�a>X���X/L�8&��t{�0T�����@G�V �PFw����r��T.��D��C�سk� ��8�l�i#ɉ�>��sPx�����9��8�Ņ�%+\� �mm*��0d{�c����ؽc m>�4\+jd�m��M-�)��3i4�^:13����U	�����$�iS3��8"a��	�J���L�o O��ƟA�#8�#V��V5iE:�~�����3�@��`f:���U�?)��v�F�p��>�8�O7�O��Y>�jdN���&��<��`Qǐ%��XR�/��x
��r>/n5-�5�i|��7�(��Po��`h[��(�g�W�젡�7ܗ��*|�嚳/`~i�+XZ�T�G�
�E;1gi&%��K��kĐ�n9��Nѯ�����J�J[�g�PBwg;Ƿ+�gD���94j��HY�4��D"�SggpmjIϬ����.�&uH4o���27��CC��E��\���K��8��E��XX��ZC�ŒbG��+oæɵ�RG�^2����k�Us��G>���w���e
j�i7J�)!���:����c��5))���xO�|۬�n�O��Ӵ;QmZ�-�����x��/;K��R�f��d��kѸ�W|g��[�5����8<;H'�Q*"�J��d���4�V�h$�tg�,+y�9�M���ێbd��T�#���Im�r�K�E 5ԣ��-�q�tH�B�̜�w4&��A���@+��M\���ȰQH�Ӊ|�"[�k���j��><��~���w�8^}�E�,^S&Ӿ[n��o��]p�������3�1�����ؽ�����~��Oj��6�n���
�>�Ʒ������`׮	�it�y���x��gq��G�	r?���P�-j]��l�Z��%QV�"���=�Cw��3$�bz�2~��ϰ����D��6�f�`�-J��UÃ}��hG���c��4��}N�؄s�xܤ�D�,����2����5McSϠ2Z�WJ�*8Ь������#8v�n��&t�w���V��;�ěo��ǧ�#�Y@����.�'�Ȗh��S�)T&���V5�b�!(�P/2���Z.Q���CO|�k��{�0�={|��<��o���G��ݏ���	���i�w���(vn�X�ş~�?����������A3��51�ߋ�����92iT��Iڐj�t/�6�E��W����+�e�p��DQ"�A�#��EH]N�uؚ%�g������PZ�)X[��������w����E	{�g�0��p��
?�b9^][]�_��_��?�7܀щZhD/���ܴrH������\����uو�sy-�cw܆D"&A������ |� �$V�64rB^)#c0�+����w�����`6D�PE�f�z<���1��k���P����=E�T5q���C+>
��k��^~��z��i�^<�f.Ҳ��9i�æ�Qc�Ƒ)�kt�u�z$ʥ�o�"�as�e'��)�����>�����'�w�0�N{LS��C�T��tYxj}���Y��ㆀ"⭆���n���e���ƀf	�Q/���ػk}�a��t�������~��6s��11��j c����/4��b�@��`�d���{�w����r��ZelO�B7Z��6��������d3�u�㧯�ęS���Ѱ�P�1v���)�-E�tc�� �AjS�8ـ��}'N����3H$J�l��Q
��Ò�}�Cp٭Hnn�5��e||qsk99>P�M���G_��va�H���ЧLق\�<����Q.�v;�sZ4ዴG��Ӆx���/Lbzq��^O �ZI�ug�O���n�Y�yϗ���X�4��V��4E��-q���M��/#_$u�g��V�ֺ��*0�)�b�t����F���ń2	l��>W���ct�;Ǉ1� jri!�Sk�Â{�qY3�sU�ry+��ep��$�;}���xPj9u8�N����6�v!����M�:)N�F!�Z�l�jHgJp��X�e��M�.�I�ka ґC�p`�6Ж�B[���U\���ܥYĒ9��t}I��s��$���h�����.tw���vY�3Q) W'1=��X"gP�FE�{�{��T��kDd�f=�I��L+�$�I��l�t�"�a���&.L�c�\�<iv�Dձ���@*�S5:�2zB�݁p���955���Q�E1?��l����.��t)�$м��Ç�Ƶ�x�a��>�N՘� ¥�*�D���ЄL�`�N��I�att�aJ�I�&�[�
�����Of#��8�H�H�{�#��h ��_�l�t�6��g�+U7S���������P\\k_�(��,�
K@�Q�gi�ubQM���2p���^3TR��J�F��"�3�q��~�Kc����U�=��,R#t�z��m��p{�p��B*�x��6T���p���{�����pz<���aw��0��'���&gP-����!�4�{&{��譄u�ʤ�㚑��p�a���E[5+&O�{
��h�(~��X���h&��S�MD��O���c�qY��A����R*�%l�0-}5�$p�`���"�u7'�l�9(X[p�����IlX�M�F�&;��ٜX����o��/����ѱm ��ˏ��{�mX]^��?��_~��\���������ؽ�:||v��c��
%�r�P-ep�Λ��~�[23y�����s/ ��A.��#���w߁�>�����_6�;���+�aan	�no@���VNIrw4�rԡŨÊ�^����r="!��^>��^y	�\�Zl�`��rJ#hJ��]�j��v{m/���Ōhsl��v���E�7?�.sm"6��e5����q7ds\�xs�K��d���ie���cc��֣x��{18ԧ{W)Wq��4~���|~���{qqvk�J<�9K���aU(�?� :�!��^d3PD-�,���#���/~���7������Ϟ�����}����W�d���m���hқ�)m�[���k����N��#��Sx�ݏ�+��d���v&箧��{�>�3!G�r!��ϭDN����D�T����z��\/�v�+%xC]�s�g�K/�fM�Mh�W�:�QF[���&���;���fa�V�ޛrB��S����(�"Q!)��z�!�꣏`�D?Ƭ[c���E<���p��8�cccz�Ñ6���B�Q������4V�V����10Ǒ�ƑKtte�JՒ��N�%7��Ga����qj���,������Do���B()D����z�?�V�(�� W����텷�ug@(�l
��FQ)tV�4ds�>u�˗Dfkҝ'�&�yX�UY�jR`"bM���&��-JST���vо�#%Z��uȢ�g(�#�݅��%�+��Ϲ��r�lu�|���CdGX5v��B"ԫƇ�E��u$�k�{��� �a'F��`�?��ύ,Gtu�&���!6��% ���!.��h?z;B���So
�[�L*񒖥�T�Ix��Ƶ���0 o܁�?4��G� [���UP��x�ͬ����G*�"�Z/��ӈl8�k�����0K�O'g���{�13G����7�6&_���Lal{'n8�}��XY�ǵ'���¹�eX�~x�4d�����n�th'z�L�m��!Q��z�ҵY,��JL�ඔ16L�_��E\~:�Tq��%\���B�h�_��{�w�F{�&{���Z�l������xV����������>���G#���e��5#ԓ���P9�8Vx�L�cWWqfmT�9%Y�ڻ#C�URB�-MN��X_M����=��49�/�-��c~ur/��B�-�V�MC ��´U;�n�PW��t8ԫp#�*$���ėד)Q�(<�%��_X�f<m&d�M8,�56�lp��	rk�9+.M-�����k�+�v��v�4�����ng���D�M��\�.����"R�Q3dA�oí7�8�F/~�.;5PK�"[�m*�?�((en�[��RU��{������Z�R"�|Á�ë��o�.p��j!���;���M���AjKC	��#g^Aӊx,��)�? DЌ�-�>i�D�X�gV0��,7�T����t^BgM~XŴ>d5-�*�SOѩ&LAm5
*�*E�cJ�����{|HS=�������F�P*�~�m2O	!�c��c��KǦ S�����:>��<N���b͊�h��}5�-���6��s�ggcE��dO�ik+�ݼz!�
ڴ�L`�L��MpH'�c� W=�@��^��Oމ��X���O��>���q�l&H�����ɄY��VЙK�k�(g,�Bܿ)l�yO1/')�Ѯ^0��.f�s�Hl&Q�0ܐŴI�%��i1�?�u�
ɲY6�Ee�h<%�zS�|�W>34�P^J�r����q�������c�F.�B�V�Ή�x�K�áC{����JZ'�4Y�p��y\h��dS�ߣfQ�ԑ�pT_����&d����z�K<��r��{���d��B�"3������B����������~%K�kul�Vq�����+���E��8>:sO��\��E�aA&�Dqs	7�q3~�w�7�=n|�O��<����<v�V|�_�ѣGE�d�P�T�����^{/��
&�Έ>�F�v��c�0;�	 �s�����e0�s���_�m�݄pЇb1���Y����p���&�j�᠘������t�͸��!��e�4wH�TLkO�A���%s�(СKnc��h <l�N����%`-������$E,�%���B���,�_zq���������h����8��9����p��Q��և�����ƳJ@�E}x	�UE�$�,��r�X[�B7��}�u�����_�����=��O�|���Ñ8m^��<x@7��X�;�M�i-�p"M.a:��G�#�U�x��H�uv���qQ6\�|N�Z���ф�v�+6̮�pq����0�T��e܈�Vʚ�J��C�h�	C��4����O�t�}�Jq�k%��[����Z��Z-�!G����Q�-7��|�8�oHE����"N�8�^xN��c�;�s�N5lJ�l�8!�����
f&�Z��2򥢊�={v���:$g�g�P1����#��
[���g�N�������?�O~�Sr����Y,.��w�v�����S����P&��B��D��m}۱�-�n���P$mF�ldD��T�k��͹��a�d`A�z�z�&��+�!h�qn5�b�_n�ː]"W��[�<Z��_�;��\�ɻq����s4��NЖ7��Z"�H����\&��	�_��-��64	C�P�"�����D�ߊm�m�F[ȧ܇r݂��,�=y���XM�n���H/ڃN�}��M�nD�K�,����d��K"Y������e3�Z;wta��6���4w�C��[aq�p����݅
��v��i�]u�m�¡�D}N�H%�6��T�����ӓ�6�F�	�/
��#j�b9�����0&F1����/�,`�8��E\�Y�U��ZNc�7��vb�0���2�+%||�2.O��}�(@�50�ƞ����D�y SK����EL��>�n���A�C]*<{:��jdl��Μ�ćg.a#���δh��E����#j�g������q�D���p���C���D9��5)h�
*��6�,�l�v���C����&���@�l��b���+W�����w�Б=�t���{��P�Z099���\F*SVC@ABY8��M��5��b|��z���VI\�_��\�8n�*B3��fڅ�'�9��	��$K�f�K�پ�h9�(�[��K��q�!C�2\�\u,&�Z�#�\Cw���T�L�7Ӛ�n��m�|y��_���z	��vp�����@9�1s�Gڅ��9�l�kO�t�U���@ c�#r��R<�)W�C62y\]Xŕ�8���!��^�*XkE�R	x��!���~�\ �N+\���	*������D���!���� ��CƉ&�zqiW��b3����u5V�7Y��A����� 5:�ְ�R0�# u	p�N*uX&Fq�7 r#����ր�E6�.����^Ęp���nk�6����G��z�iO6���+�x��)L/���py�$F�tܰ�/��i����\���40R��Ǹ�!��V��I�H7_)�M
n%O-���ߍ��=���9��̏��s���y[��g�� ��`@\b>{DO��r��Y岀W�F!��|6�6�>:	z5����,Ъ%�R/�4H{#�LH�m�ݜQ���Ĝ��ݫ9(W��Ӟ�׍Șnk:GZ�:�Ɏ�Z�rV��{�������;;T/�I�i!�<��:���L5f�p�]U��lv��	�d-�{h2�g��n��{\N���و�bҮc�<���S�������.����U3ڒ�KgI��f&��=�US���x�ױ��!�B:�D-��[�����B����}�1��'/jB>�k����q��T,�q(�.�̹Kx��8w�.^��x�����H洄�i1,����i$�_!�A��|�ˏ����}�]X[_3�p��ill����T��@(���vD�AXmu,,N!����c��ppG��P͚�zIS}�at76��PE�&i���`�ت3ج9j�A=�6�*
t"�,c~j�.�`��`j���.|�/ad�:=��$��k����Y\�gqm9�,�-�S�G45�s�0Жu,oM�Z�dlJ�X��;?��_����3!�/?zu�w��w�b�����VڇRDC�x;�I +㚉q�ᨌ�]�gYo��q�Ѓ.#L>r`���j(�s�j���N�Z'b9���\�)��B	�k�*�����F��  ������7�yS��
k� pPhS/
�`V�6�f�'�?��w����MGvb��CӐK���_���,��:��?t��-/�"�LH��Chb�NY�}|�,��`sEj5��#
L���f���!�$wF��H$�<=5��s�-������L���{`e#���]X�����?��;H��>�|���9���<;��"�H �c�IJ�MY�(_(�\>��u:��UG˒,+�)@�H�"@d�.����;�;a'�鞞����^=�_����a�n� 
؝�y�����󼇛wV`ּ0L�P#��"�;��dVR���+�Q�\����f�H�z��F1���*�[0U�f��b�[I�ݼ	��Р,��N��J*� 0�g���)�C�A#s-em���pW'�{�#8��=Ƞ�d!����/��P~��B��i+�s�5��V��!�F�SIj~)!�T�&z$�Fw" ��,�!NT��Сv9����团��L�5������D�d��Z���xd��V���A�e�B�߯\�,d�*'F	�R�=~�:6����^���"1�L�޻���^~{�
��� e�Ξ��^x-M8e�gF�ܜ[��o�����狡EJM��hYA�Kc�	A��=	���s{n��w�-5e�CbѪ�J^��+��!q!ShaymG��{��ٜ������	!%!�jS�B,B��h���F3���L:�=uGF����(�'�lP��vk��< �+�ܬ(x�**��Ŏ�X�A�A�n۳'��R�Zܶ��Si�����B�i���!@}��Q��MhZ���3s�61���=)��DF'�?�@�@��"=�p��m,,m����DD�Gy93R�s�
��`\D���=\����ʺ���^�l����N    IDATr�&(������z��PE#a�'Q�L���0�݁���1�m]2I�{������,4gPҝ)�bC@��~j��Q���F�`e�8��I�����|?$�ݶ����qx�W6�!pb���&�޸����n7\>���J�<;Ƈ�1؝�$S_CA��M�MV̯�ཛ3X�Nð���`%���Q�O�m���9<|nva!|&�]�˻�ާ�����llmK(���)R���^����yn�6����L�i�6,��Z3Poh*����M��,�)���ix���bah%�N�hZ��G<�?z\|m�\�REV��l����=�|2�p7��"=�qdd G�d�æ��00ugo�{�LwH6��-����h�ddn�H�S�����MY�X#ߛ�d����3A�Ԏ[Z�xQ�3��`؅W^�.���K��Z�)?�a>S��p+G?9V�aQ��w���SM��gsBK�9'�2-%آ�� ��[2��q���k�����HCc2��I��ө6 �H�̗�;6��0�����BTR�ڐ�Y�FB���G3����BCj�����U,��
YP�˪�p���o�iV�r>���Ri�,���8���(�~�)��Z�f9�*w8�)d�I��SO=�s�=�|��?� $@ۿ���w�����/9=|��	�ܔA��Y�+�P�����_ċ����޺�b����]�%�Q�%������ob���צ����xw=}���{�E:��SSwp��$�_���V�ԾJ27�{_68�A���A�+�7�Etw&�_��}�i��vb{wo��.\|�k�F����{D=Q�汻��b)�by݃��8Ѱ�Q3j�W�܀��/j�%�''�WaGe0G�/�v.k>��X�Q�̍� I,n8,<$��������Y���cur�H_��/㉇Ǚ��d������y?z�*V��`�r�Q��f7/�[�`��hi�b�uc0�6��=�ؙo}�>��������Է��'��N��~X��ɫ2��%	�13ʞ9 �n	�	��j�`���e�-W�F� ~�,N?���F$ٍ�2��UL8�v$�-\���k��X�i!_!�ϩ�����MREi���$���Xs�^�,߼ �v`5W��D׬�
��B�nҐ�S��`�hX��C����FgGX��}����w|>/�XB�P*���ƺ`�fE0���S(U ��zG�%��2�7�N!_ؗ�_
-�	�ݽ�G���B�ݹ3+��#G�bhd�l	޽��~	�x?W��օ뢍͕Z�io�]pz�����v!Snʕv�Lf���&�Ey"����A�����+	V��T�P[�^*@��>dn�qM��J�e���i������ώ�ge�����Ob����7*�!8h��CMnh14��dX&M\���$)1�bԣ�D�I?i4ʈ���
"�#t ���7��v�%�-���������qt��<x�Ps�����b��.M� Wb�V�ȔH��9��$�E�_)����Ã���X7:Cj���k�9�]���;b-��c�8s�F:�p[��4j�<k��1���W.\��N-�.W@%�����ZC�d�zU&��p #���ܘ���֞�j�mb!�	'���ja�S�h;�)�����I>?ߡx�%���DV�"J��m$����D��BhH'7������NF�k� �9n��eܘ����$C���PN�iz?�e�R=0a������Vp�2�Q^"�P�>3B�jgS�����K�5��Ãy� �\f�����g�rC8��_@��hFGz���Ogj��]���Y�lg`�xa����r�G|85ԍ��L���]Kg05����%є���CqTt����V8�.���|�y~���dCcHC�pߙ����d��2�r����%L�,�ڴ�3�C�8�b!��8>>�#����� 
UG:]D�d`y-��y~ߺ�mBA�4�}Q�&B|�`3�"S���%+�M{������dkz.'�^7���u�#�����]��W09���7��큍�lR�i�?t�?$�u�D����[ť+���lN� ���)yR���N����S��<'8���G| Ys������b3
)0�8RҪ��Y��p��B��et��%	�
y�x�C��A�L��`��L�;����`'��&C��E�)��Hx\V���{9N5�|��M��8�[3�R\p �).�9BIbc"�^�Xפ8⹠�僠��:'DVǢ�awj2J�/��~i6�zj�7��8����-���O��^�ì�染|�V�S��!��-�S��u�[-�9S�;��<(��<��X���s����"���_v6̗>�!2f+�C,�U� م6�p����r`���f��SPޣ�2xa�5�jv6M-1A3h���@��2nT���N��� f�����䦆����u^+N~{�#�ض���� �pz=�կ}�����8����>����ׂ���������SO=����D8����v~ ��d�W��O߼(�Ê^�����=<����O���8{��5L-T��4�<Ei�$�$�����.,#�)!�-����nq��D% � �4CjD5�]_��/����"a���ο��W.!��/�[�}�
~��'pϽg15}��:l����1/Z6V��f�I�����,�$1����HX%)6K����J����y�ܵ|�mĆ��t�i�tւH8�#���!��1yu/��m�\�F<އ��c���?��O��ܜYǿ��ą�wP��K`!�M�[n()�f*HZ݄f�B�A&Y{�����ڗ>�����7�}ϟ���g��N�Od�2�EG�Q�hs����ҬR��i΢��j��YYG�ێ�|���I<��Gp��149��D� J^B�T�L��«o�bi�����#]��N3���7�"R���ݨf�Z�#�q�w�B�[�f�����6���*��$��Y��D�1��a1��c�>6���ݝ	�:{�Luө^y�!�>}ZP�4g�ӫV��C&Z:^z�ٌ0�x��ú�7y9��b���^�>!Jx�P+�K�f�O�`/���1x|�u���9�ý�H1=���d	K�{��J6?|�.t�l����h��m'o�,W���ds4���d�q���6Ѣ���4갘��B4�z]�9x���㝡.��:�BT���M�XX���N��g��ч�C�(c3�+��T9��@�~�!hO{���	X[S.�<r�e
�6R���tC�0���m���+�C,�Dg<(�}6*Â��.�S�Ǎ�ہ�ׂ�#�8{b>��9��ؔM�Zƅ�o��dl�����
X�����"3��8v�_���nT��(�`}{ْ.�Q��Q������pld�/���\4�p�������b7� !��w��+X�"n�R���>		P��|U�g�0Y�r�`��%��hHi�N�^�.�@N���K�K����9p[�����u���5l����̪|�fGHz����^i��"p���&t�6�x��ܼ���/�ԲБ�Fy�.�8��T��l���0��۫`��qH@��<;ju 
�6\J>������G_W{����֨Ѹ�>ɂ�:޿>�듋��2!��]��p��r33�hY�����iI���q:d�mE�Ǉ���BN&��Z��4n�-ana�|�>w-�U&�:�9�*|�I����l�O��S�3>܋X�+^)�xߚ���o"[n���@
�jA���9��D�Y�6�܄�]���N�JyJE�;F���"~'4)����jX��b~uW�2�*�~����u�iZ5$b89>,�W���_`s��w�M�Ɲ�Jy�a	ecրQ�!���N�V�O�.�!R���O`�X�?���R���!��*��:��ctd@��_|CW�7d+E*��6�(�����������[2�Pmv����1TzUbk�tG��G%�$_*A'��j��掐^�6����ϑ����1�˰(2�?r�)�<6�X�'w[�,,'qkzI�/*�&,4	�� M�j�*�6�1�0c��iؘp8�b�P�{��۴9)�ـ�:��Z��^��Ҁ��í�o#��H׸l}��a!H���;�F��1�$��g1�L�L��?���q��-?���D��0�7ᦀ93t�S�(�児�	�V��? �T5�K�6���%����6ى������46-2L��A��U�����Y?�k4U�6e(ԄĂ����ϱ%nh��`cv �:HNgax��Q�7��h�x�j�?�ǉ���ï�_����������o��E"%q#�C�GG,����82�޾Nh�d4[XZ^���i,�m ������r|�G�K��Y�t��YgX&� U���`ye�_������X�E>_�Q��.���r%�R��&\��^�����"��������5��%_��7_õ�kHg�������qA�ӬMi�������	V�j��@��D����$9���ﬨ	Hlk�����p%���Aؠ��<�4��!>P!�h���h�������5�J����*^|�U\9]�>�̳�§?����Ȕ�����y���/�f�C7ȷ�ׅR�.@604�Qd�[�����V��j6Y�����7����~�d�χ��_��������dw{��� ��Ύ�VFݠdH�҅�D+�Pl*}�*l5ͅz���� ������P_�t�,��B4�Z�unΧ��˓Xܨ�藆�+O���G�)"�<�x	֕O�i���6�ckaFy(���b��e<�g&P"B!���q��3,h=�����.z�;�=����J2��h��_ 	��^��E�ϩ*u١PL>RȺeC������r�ǉp������u���W�
Nq�i�$���`8�����lզ�+�XXNc7U<��ȁ�{��7��\Y�jE���&������^7��i9/�z1���J�h���F0�5^�A�
�;u�������*L�k��͠j��^4��!x���ч��n����Z�<*�z��!eZ�0����� x�v}���� eRn������v������ݬPYV6�3����C8<څJ{�j�"�'r��x{o\�o��`\
h��H8��$�er�,N�Za�
�EC���̤%� ](c��Rs��H�MՑ�>���1ĊX2�+]N\�u?~�

JJ�{9e*� �V����⡠�I%���"��24��ί�ki���d���\�����!��x�n;:�L��!���s"����t����-��,�gi��$��nm��O��,a|�[<DE����4WS�K�z��9X~x�4�I��t�����h�=s Z�v��X�Mc���?k$y65Ѭ�P����0�B�Z�լ�h�rn�Vq��&n�����fg�Q�F���A�@�!![�lW&�1=���ހ�OskN��#�����Ah��v�����0�����5�%ɥ�J��N,?��<8�e�KzIS�3�3'��bn ����F;%���?�f��q��-���p�Ip�K���x�':�θ6^k5���sxo�li~��S�y��ѡ>��t����hՉ�4���ǝ�u�,mI��DŤ*�_�eb'�U����=����F������XO�`���|���h8}�����iB6���ܸ��+��(75�Ba)�9��/>�R7���������J����l�o���.%���3%��&��LuE���e�!��""9��MhJC`55P/�e^ۉ�~���vI�Spm./�R\�:���s���h��d^��"�$M����Ȥ�;�x���q�p7�hg ���.~�d*���2�2a����ቲUYN��ٍEC�g%��9[8�IK�R�f	N��
�P�Y��o�(�d[�s9�A1�t3'����64��"mg(��j�Y��L�4>Ϛ�^��L��Sn��b���p�/���;`�@�Zp&�>����{f�ʟ��˵�|Gm�����|�"2Ez��ז&�BW����)�#e&�o�O�������H��5�7�����puϵ���I]t��{df(Xa6K_��W��/�/����?�3��V�@h�כU�E8T�c�>�s�ߋ@�/D��.S~s��Oa;E�_]�Ň��d��)0��m��2�ze/��-�g��AVf�,$/�vYx�ڣ��ܰ�sXѐASz� ����~gO
���{p��5$�)������`����D��"q#�B]+��(A��(�K�<=�bN�|��m�o��������;Ndk-Ec��{�`>3A3�φJ�*Y���\z=a�!x1h�b~j?|�'�~y!g ���g��O~�@'�����?{&����e����bC��Ca�`n�`���XB=�����_��|�D��G�?�������/��'�?�ć�K���Dj�h�!�
����uW|fI+e�"V�Q�T�@����c5��H�d&@[�-x(��&�[2��|/�6���:�.�,�n�qe��6���0��f1r].`s�:�'/�YJ�(�`�e�*%	�0x_X5��a�s��=]��E��+ԡ�8�O~�Y�vv��Bo���ޒ�bnL���"�!)��"�vv�L�J��p���yD6ņ���D<�!ʐ<^X8108�Pz|\��m�*i�g�37�L��@�S�AK�i\�\��V[I�j����� ���C�XE���fE8�b�\����I�!6&��"�B��u�6`��톀�/]$
��SIJ�r�|ß���uR�]�1�U��H��g��a'�%F��^<�ܓ;w�z{;���pXE���A���h���F��0RU�}���߄�"U9	ꎋlȦь�4����Ltg6��-�����='��3���E���ֽ��~��e�#px�"��"'�⁠Q��~C��><.�.�<#<±�<�wuB�H,�@Ѝ�ׄ��C�(b>�z�h�L���vy�޼+XY�9��C*�Js̓,ld�+R�X5!qp�}��gA"�]�)01�Y������~1?"�A/�A����vj�=��յ	�"��LluZ��܇V�bXn���a7[��A$&Q�7�� ��M���h�*�ߡ��!/DfV(U�$�� ��nH��b�q�+Zd�-l�,�?����b�#�
�������L}z}A��r�$�mu���ۘ[�E�cj�9ģ>�+�I��U�9 Zӫצ0y{�Z]&�I���gp�7�V>+=��Ŧ	�J.H&�@�W��. �) S(K�S����	M3�M�.���� ���f�k��X/���R5^��[���u۩�K�}ܐr���G9���S�^,������ǵ�u��4▆���٨��p�Ό�'�E�XDS7!�ӱ���;��X�L���u�,Zl&�2e��uvM�����0��{��fӐJWq��m1䕫fج^as�D�؃'���`u(�-�N�bק�p��*��� l�vP�M|$:n��f���:q���z�173��Y	��;�2�㦐D)�b�^�ʪ!��Ŭ	�efaؐ�ܪ)�Ǌ3GFq����L���	-�6i޿9���hN��Jnm�e�6h�5d����1>֏��A�;�(�,-n �oH��Do�����Υ b��$�$�4uZ�*�@�~pN��B���j�I�;'�,Λ(s0�
�4t�=X�����h��pY��ᆋA�-��K�7@����L�Y���4�ag�k����Kx��?�$Ų�:7c�M��O],W$�@V�1;��l��)bӬ��k|ǕY�@Fx0�� %��{B�J��m���-�L�	I��y�(���f��>U ��/T ��P�H�N��*�u�&`���E�	��ZJb�3� ��[�2f�f���>e�5�����K_��+���o}��d�bvXPmV�)������/����7~���Mt)�d[�TdyQ����}�v��2�����?~?�����+���R5�3��    IDAT��סY�0Z�I�S����'��k��4���1��g�ů���dj`��ܸ9���5��U�|nDQ�A�������@��C��|��=hXjh��(1���$�\V�����M�ڰ��)�x���->�J�G��1��������l ��0À��.������ayn?��˸v�*����������z�'/ /����'�3��I���D��vC@.=��>������_���|�X׺*d�~�����������9��O|���~�ӈ+p�$ �CUjJe{��]� �D\�'fs?�Fڹ9���[�(ds�y���q��'XUÊ�BW��A0�Mfcia��.q�7Y�rE�&j�!z8���8l�^�.l�\���;0W����s)r)�xP�l���(k2� ��tX����������c���w���V�p�u��6177'�Ξn�a)VcM�]��ueE����:]V�vv�;�"����OG� ��4P���dm'��YGW���l�YZč�Y즋�[�.���<3LX��K��4](ևS�L��A��$��zE6n7	!�sw٬��
(���Z]FugMi�qh���.e���(���̦�/�2x-h�����%�P�ŉL��<�1x�8��<�3i�Tr��U7�Kj���	�P5��o'�<��u���62�2n��a$"�:,��i4�ڭ������n��\7��;���.�Bn��N�1Q�Pj���x�'�`u�����?�*js�*4��^�rp#����h��.�.#�˵��:�5��:z�!�F���»_K���\��e0�"!NMa��sapͩ��I��|fɈ禌+Y1�x�RS6�^U	b�"*춋T�#�E<ꃋ�%�Zykܺ����cs;�+�/��������*#�40���P�Lj�5��^����i�;�<-x�״���R�U��֎�Y���8E��r�E'���.&)��s��􇐌�٤��Hn�O�P)��aaXڑ�N�%p���2�rzBXZ�Ǜ��ܗ 7��Z17N@Og>J_4�4�l޿6���T�u%;^����Ν�HĦt�Ōxjf�����v�6�@!�B�RG�Z��KJ��vӨ45�H{���*�t���X�%� �j�^�j�6S9L�Y��ZR���vNo��(`���=t����{��n'K��WEx�!%�J[g���h7�H�`X%���lV�9��<!8]�x�0,�Zv[K<(�c=�i@j
��l7n�a�β��l��86��S�݋��@�Z��E)[[�2��Zč�U�f1(�̔4G��;5�����v���0�>/V�WE�L��&yf�L0]��6~�l�H�t;��n�	Kd���w�3��q���85�@���9�mn���l�1���;K�QvdqJ�?D�̀@��6Q�g�T��#�0�ad2,�]�Ѳ ��㑆@B�^�2��Ɇ����[m��A,+Cq����&��9(	{Kd*����
�������6s���L���C�;ͅP4&hO������b�ڔ�����5��	;�fWk*��r"�����1����I�H�:n�W��~�܉LGɞ�p�B� G@L�jcȉ=,�?�W�>+d�k#BEn	��.Y8&�;���l��jC������C~�2x�(mj�YA.�TK�Y�pe�B"�Wάhp��M&���92LM�!���v6��F-�_����_��H��y�}|��~��t:?���A?���'ŵ��1�ׅo��_Cg�l;+���O�UT5��UQ&P�Q,a���$1����x��Rh��:�����
���fBI�D�%6�a��8rr��?����CG��p����q�*�FvB&e�4��$���KHv���;G(⇍�o�/�@��@�M?�lL N2 $��5
�H��猍@[r ���_��a���Z�(���攻��
�Ll:�l\5����.�\<���t��7~c#g�ÿy�������6��Ț�$3nø!�ĩ�l�AOX��Zn���s~�_���|����GC�O��7�������=1��ǟ�֬��������REBk8m$ݡ�-�II�jECg�[�J�R��K����#?,y9!�u^��s't^2yS��x��7�МQ1gP7kjT�Iި�f4�K礁�?1����ܾ#�������\J�uihdke\5��v;�:6܅�}�	;:��ߏJ�$]8��<�I�����y�֐��p��Л�]����)��e�n���Tj�lZ&����gN�������7�4�-�N���:*5R_�x��ܺ����$��5*��F�l�+%�A�AI��j���B\i�&,]g������{)l��#���Fr�Bh�5˩7Sa��69�~�"TSf�H#�S���Y7�ϏR�%?4 �u�s�������V!�L�(/g�ȕ$�H,jL2��j�D�e@�x�L�Ĵi6�ed4a�Z�AN�]�B��C|���=�H �]��U\�3���e��?;ћ��#��`g~��^����#��W��{7���O�
��Ϧ�U�ܸ�M��gC��%�,�@��{���`h�S��z�*��]R�u��p��R��v	�(�_��fo�w[y�\AXܤǰ0�a��o�JY����eij�����.A)�P+W�;����\�38�	��@��BW4��nI[����4��� I)��1�������Y���n�����C}���4���V�^��:�YJ�8q�����9f0IV��u�{y�v�ʤ)1Ι�qM^V��լɆ�t��Bv?�A���Ō%�d�a�Y����'�`�3��,h��uY]�,.,m����[�_ޕp=��?���(��A�u R�
Na��H����%]�����pb��!'�Zz�x<ChB��F:�wid�ƺ�i��:r�
�u���%�0���I��;e[��J����#���[9�������3�_ޔ�:I�m6$���?�8�Z�LCY��\��]��~�N�s�io)s�">��<z?�A��)�h̝�����l�����I2p5vj��	p����p��0F����ƱR60=���������pt0��>r�!�RV�M���}��2���l$\>�|�Y,�LVE�>�\A�T�m��M��� ��Saj(2�x��)=�.�g3ٻ͖'��6٩�ef[��If*�ڪ��5����C8�C�VF��-L�]����Hf��G:��A�L�Y�r�I=IR2٦Ο�|[��+�;��v�3�0���'��lr�˂�}���)�v~B�kû�N�h�U�!O��R�Ӭ�e5�h�SX�|���pR*ܤ�W�qcG�>�"90dQNz����Ҋ�w���>2�=��x���af	�`�[I�<�L4%7E�s�|6�_/	V��5~-2�����J6���+��k��
$K�N�g�Oj�P8_���ޮ� d�R�����������8a28�	rذ��%�nz��/��9��簋�:��*C��;d���%2?n�[��x����g�q��_�,���G�{���o��d�$���-��빧��>��݆��*�zG���s�y���"�p������F�(\zB4�T��3�D��^�O^~+�ۨ�L0D���%����H�݁Y��	pB��p��8��+_B�`B~�ć޽;+�a��5����Eܞ�B���/�Dw���p Vs58��ň����Lm\�`��l��.��| �����=�<#WlĈ�&��M�����hK��ŭ��O�e���#��i����0{{���0�N᧯^�K/_��t!]�:���l�d�҆f(@��n����{R/�T�y���|�+��w>�s�|����� �wh���SJ�ު��2��{p��i!P�r���������йζA����rZ$Q���x'���n�� ��� #���jMRtÁJӁ[s)����XX/@s�`u2����W]��q�*�حnx�N9��]�޾���@n��,��<X<`��E�Oi�������O���Cp;]��rr)pE��6�ړ������*\�1!S'^4^/Y��3r�[��l�H8(	�^�f��9���^�@9�p��,	�-TY�p�Ey,2�M�pub��u\�\��rJ�@��P �@G�THV�
2�,�������h�hH\�ɭm,�/ ��s.-�a���e<)B\���R@>Ѫs� ����ץ(�Nf?�%V<v��J��o�s����g@�^C�\�iN6_��@r&���͉2u��K��ߤ6�%���Y%X��?7l�4��&���.1fE�NxVa.;�v	���qg}sk���c1a�+��xHB��6���\0<�5`v1��߿��}I&< ��^r8mQh^{��p�������	ٌ|��\똼5#�mfb��ѡ.xm��0��&>>W�?x��+xj�h�l�[Z��h4JJ�f#��;�r��0����-%�c�5 I��9Q�l��&7�Q�ëݱN��J�kXT���&R5̨�[��X��ce#�t�
�n�����;SN���{���ݪ�}<p)��	�㦮Z��1�N�';V�w�<���/N`vi&+͖��I9�{nG�&ʺȑ��Rf�` �B�6H�rH!�qScn"�`t0���[��	�ש�5�by=�K����DV7�^?�VMd:D�����ʳĳ`s{�gW1��ښ���Ɔ�8��ȹ@2���^�2}.	y��H���*C�J͌��K�<1�L�,��:"-$��]Q/�z�"�
�MB"�aniM�X�˗ȗ����Q�=yB�++��M2,�8y{[�2�U�$уBS���<����XDg΂��37��1��)�Z3#����4�,~�$����&���H.��g�e.�cei�]��b�G $�'F�����$�XL�fn�o�K7��.ð��p�9�_����E�.u�ي�$Ц!
�y�/�|�Ď	�*j�hR����5b���`Qa����j�̼��܋A��K��Êýx��a٪2`�dwcaso�w�۰���yê!hQ��h3ͺ.K֊$��[�J-%�`��NL������ިF�@rr��+uO�Wá���*e5���Qk���-��J�<Wex�M�Zl߽�����c]ȥ�������HK8T�`QvK�x(�R��0�.��ϊ�R�X�9�n8�Ԫ,�lajzK˛����3�p3&]���ߓ�>���A��'�ɼ��P�V�	�����&��S�ln|�P��g U��Noo'��Hb)�-+��
Bѱil�O��3��Ѱ_h:3wnA�+�(�i�iW�L~�X)��C�9U��FP�(�7N��p��Ty>Rw����7~�x��GP�+x����O�}��z�y�|�ӟ�P"?��en[J��=��������S�ܥ_�d�Ѿn���J~���ە��ʦ�*���z����/���E��(�U:\���aS�ϧU㠉��z�x����y�˥���h��]�����zVB9Ý^��ek��(�$�<r�T$�_�Ī�i���,�=Rj��j��Ć��8L)kBVD
�������t.ލ�R����1Kj�>w>����v�/��>_��fU<�w�����@���IS���&{���x(�oq�M_[��f�'���o|����G��N�_��o�З���ċo^����v�iG�F�G���'?���n\x�<����He��%�GUΈA���8Wo-$�<��S�;��;�3848��'OH.��K2<��y��ݘ�I�7�qw�(&E��Z���z��V]&B|H$�Ns��`ѧ�\ˉ��MAy{�Z��t�l�x��?��`?N�:���.��:�~3�=pV�F�r�Y���ؽn����ЦT[�����c~~^�8��h)/�A:��ΞN|��:r~~�tZ��9�9u�`T�i�%��@�z3/*��Z)˺:����o�o�{�Տ��	8=��@�gu�_��&�3� u��h��x�F�B�hTudRIl��cc����lC��L��t��U���5m_:N���*��fv?�g>�9�C���hU�Ɇ�Ŝ:�����02���Vs�Q�N��U��4`mc��,�`c���������<ڭ��g�y8B�T��>�7�0���L�E��]��K�7ꃏ	�v���Yd� Y�*Ȅ���*�ޠ�l�Ĭ�-�M�\�<Hh u��l����فD",���s�e�W�&�q#�V�=�ΰ-��kEŽ�9�!x�wqmz�D?ܑ�$��Y/�U/�D�cL��ᥬV�r���=yl��J��(����B�`3��HL�:'3u��ή0z�b��IJ9��6����uT����GnU����v�3�kN�y8;�Π���q�\�AB��/�!�+lؙ2��^�ko]���&b��~U+"ܭ
��@8�B,��3�ٜH(��n?[���Y��b��A$�}G�	�ӄ�ǆH��ǁR���5�,cq#�������*�D�+�x�9-J�*��7qsj^�k]a���D���a����i�E1��_� ������4�C=��6&����*5�u�Zv\�<���I��VYE3��͐���k����;,R����/�
�2��I����Ӆ=� �!'*�*�
i*��y	�Z���v��˯���0�uil��$�^RW��!������]�Y�B�Bt�]?Y�)���<���]����0�����
K�/�X[���;7Q�p��z,83އN�ok�Y/�t�jXp���yi٪	�PL��rQp�񈡙��ĝ�������&�"rS�T(Ѥ���OE/���dg�AT]��8��u:0�ޓm����I��b 걡+h
WG� \!?�6���[q{~6�a�A��SV(�϶��  ��)9��ͳ�dsf�����*�x��Ta$�9�I�N�vC �kN��4͞I�,�ITAY�Hsۛ8���0���<�#ý�A[Y_���;�[\�~jO6�����R��*:>?���8�C#��E�z�
bP���e���-�2��o�/_|	�;��=�V���j�M�
#&���42����5.���8�� �:{�L����I�,�9��D�թ�αC�������H$��[^Z���VW6E
�-$?�H0�H8�B1���9	�c�֡���Y)�����ո�f�J*#�v&�����W�4��=��3�`:aK��H������{T|�צ��;/��_G���'�{
�|�i�9|>*���g�JY��i��޻���^�3����P�1<��C8v�d�L��	u���=]]���)�M����_��w��]��f�0ds��Qc=��� ����8S��Y��"���G��x%�/W����U�	:��$"'����4�+U���s�*���K< �?@L���@<��"��r��~�so��I�w	���^*�#�-Qa]�sE��,�+*�<?\6�����3���^@���݉卼dҰq�ei�(�2��B������F5�Va������o~勿�s�����ߟ��7.����v�;�07��jY�tE��g���z�����)��Wߕ��x� �-ME4��v�M���|����ƕ[��~'�������r%/锜s}N-|�i���4^zc�|q��>9�T��$W7��9��R�p��I FӨ�P�Y���$�'QJ.�lƺ3q�*R�@$�ϝ�Qj�qy�N�R�����/1�?���^�D���Yt��?/^D4�u/�gawθ�|�>���lll���,ҩ]���s���Ԅ�k�jM./o��,��8�E6�Y����-���7h��Q7�219|�� ��M�gh�2d�*�/�C��L�(�p:��Bg�J�)��R.�b2����M�`C�mU�c��C��	}�*_�����r�dC�9tAV�b#��qs�?��M�T�:��]�8�E�*�N��RGo5a�Dj���a	�Z	n�E�a���_�Ύ���{Bza�W*_�%    IDAT���Agȏ��wE�Z�JCL�4�ڱ�,���S�r�.\�(�ހ��(S�AC�(���y]v����N)V;bL_�粓����*�7�.�u)Rϝ:$�׊&xԑ@i�߹t7�6 G�jdZ���!��:�#N;+%5Mcs�ل��Ï�i�� ���
B�ir`!%vɶ熂27�n���Ɖ�#��G�7'��ݸs��!r6��L�'�дj�ԣ&l��0�S�2rE�f��Ҿh�]^���\�/�nbu#r�ܾ��_�l5j���튊.���|Ge�ca�d�L^�׻�+2}��x����슊|����s[��A	���4��Z��F-��$
�l���7���8�l�\��1;���yR9���=R�r+46�'[*���By��>V���/א���V��ǡ�^����R����'���n�^�N�ݰ˴Z��u v�������C���8���dSJҶv�E[��8F��$h�RR�J��ť5,��#�.���aw�d��kb�w������}29�3��)b��nͭ#_��`Ѹۜ�� 5)�(�1���&]1��bl��D����6�_�))��$�C�s��B�����R�]����Y4L^x"�T��Le�&"d%:�I1��ud�T 6@ɿ���FN:=dz�@��􆜑~�N6�� X�^m�yX�A�fT�ڑ{�4P/&��׍��!��Y���.c~ynoW@����B@a�5��LX�F�ŋ4<�9�m��=3dA&�b�A��LnUک��w�R�{�)�L�ą�K���"�cC�2��!8��g>��c�53��i�lobqe���"{"0����bA��7���phh��F{e��
n~��^Xq��\��߹�?y�y�n�Wʫd
M;� ��g�yp?Jդ��|�j��|N�1���!c``H����|��ߗ^n���ڐ�rp����O<�s�����͛�����vm�r�*jٰ����K�ڡC�8<>���~��.�����g�g�<��\��D���%��7�/���x�|�(fj������������Ҩ^�1���2�M�F$�7~����
�ɛX"Z�[9�2�X��ҕ��7���q��5ģQ=�U �x�i<��3�m�����		H|����G�BggB-�L�m�~�o}��v�$�D$���%���V�ۖ4u��ǃ���?���)yL��L�cm{v���0�a�7̎�BL7Mr#	��́`\�����`>n������h
IN�=��#F�9T�Q�7�js��za愜!l��Y'���f�m�`j0�ʅh ��H7n�|�G����%HRd�`�p�%�Y(��f�%e�¯��3��V9�Fa����|�W���sG~N6_�_�����7���LtۼQ9DMF�V^;>t�>���08؅�S�W��oq��|�"ݨ�*5.�����=�q����bki'ũcGEW���*�Op�&�U����񛷥!����a@�T���n�8iN�a�_X�aC�+�,��˲�L�݁�ߖ�B�E� �l ��z��̧$�~bjv���W����HD���"r�Q�O�P>�h<�9�z뭷�+�p��1�1)�Z�����b���$��,�t��#,���!�����Ԭ3JJŁA�����W/����2L� { �O�CG� s�r>�M���9���Ϥ� ��/�;���s�B	V�,����h30�ԊS��B�g�!u��喀���@3a��q|���Bl�i���tJ��5M�<`|�
Ѐ�0�L��.2���s!�tI0�L�`@pl�t�b^23�x0��-� �T�:Rْ��^�^�V:/SB�ӎ�xP��� �Z]hAV	@2��,��&qej�H�4��t5D+Z���ZY�W~�݉8�:B�����2�����˫k��	�T�-���NFWN= �wM���Z�ݘ�z� g0�7 [6����4��7[�d� S+�W�y8re�I ���Tq���I
"&��Ѧ9��d[�n���&yj���ǩ#C����4Y�X����w��ʉ��H~��!�Fw�)�����5�WӸy{	{���6�z��BmڄN�
ŪhWC������#���H�#vH�mC���Ε�%��d3��U��.ac')����^�&���l��ڀ��eʹ�����X��V��G��Ƃ6�G� ��drH����*�n�I(U�ER�!��D<�p�%�"��
{XX[�l�n��
��{0���'�q*==G��v�*�T���aG���a7�������iwV��ۘ�����4�qy_x��x�w����L�cquS(C�`�b4��*e�|1�vF�8qd�	7jzS�|����W1qkْ�'(����S�/���6�l3:��I�p@���ĭ\�:+�)nr(�:{x��B�G�'~&�x��MḼ����}Jo�@'�=B�%~l D�HiY�S�>l(3���Rn�֥���j���g�yh6C��1����P�_X�̣��tI�ު�{1>�-~S3�`�'��|�!�'�,0���%\{ɱI�R �ۍw��ҲcC��� y�%�r%�-	��ɭh[�d��!	Aj �麨V�m7<���
Z<O�ux@�����tx�x�0���Z��T6���M�R)ih��vwS��:lv���0Cx�6��A�[4�tVJ��˧aW�L����"R�y��r��m��-i��!
b=^�4"���=��U�"M��(c�����>n߾-�gJ���pX��!�o(�=r��s��˫�X\\��Դ4��NJؚ�)��Pȇ��.><����������<��{�m .:@ {'ER�DK�E�r/��L���dw���nf����8���;��[�eYV�,Q"%�^  :n��}���}A���svN���s$�p�}���-��y��vX`7١��pSL0;?_�i�dL��+�������7�~W��7`�V��G�����Ï�'[��O��ӿ�-ܡf�{�}ػgBV��[-��p��udstv�J�/���ׇ��� o=&�N��
}���}�Q|��F�X��?�#�:u�l�<���򻧧.�n`zj����׏be%&o6�,r9��-��e��m��i��F���C}���M,bauE5�p[ �v?�6=�.J�|�,�;��H��k`m3 )�BZ�wUC�s�-[!O3����,�~=�O|�g�9Ai�ZC �~kT1�J��6�����t&�5UE���49��n]��į~�:~��W�J�3�dC���b��h�|6M�m����HlZkjم�=���?~�?��4��߾��S�����1y�Q�s}>K-aܷ�s�<�^{�M|�;���|�H&jک5`p����������~����s6���&�5���7��8S1��d/�}�s�Ai/%p{-M���J�S��\�$/�_�bh����ZDtf��	d�3h�@9	�$X���áC���|	]==�11����0�yi����b��=]�p�.��U!WL,�9y���y155%]lww'��x1[PU����Q;�.n����s�㴡�+�Gy����.�<)� �po&�ǵ�Q�����׏!��
Ҫ��Q)�hݸw���3�_��l�����-�kfJ�D6�p?^�����(��H-."9>���^T3�H�@��φ��G϶�8��� ۨ#Ỷ�I��S�)�����M�C�N������*Bojo�5腓i�Z�z��cX^\A���^l�t�;F{[H�<��"������i��q��L[wn����V�,��a�Z@d�b<�������a���_Kcq���R�bV������<��-2�"W;�Jcbj�3�P�^椫���f�������,��z�z�M�^;v篍Cos�����Jæ�|�xJ8������DkGX
N��n-����ނ�x�D�
�M�l��g����Ј$��j�&�"�[�w� |N�0����-�8s�&�^�M!C�����{��ju��g��㖧a:�����b�eR1�l4���<,�۬y�k�x�'y���p�oB/���I��RL�2�����[��5pct
�#O��tώ�c��m�f�L�������x��(�r0X�r���I�w����k�b�`0��U,��|�&Ƨ��0Za��Q.S�O��v`��GTj�\NL�,H،�8��=-�}pڬ���M�j<%Ġ��e�*Iu����[��Z^��͛z���$�8,Hkaj��s�$���H�Ӂd*�D*#Zv�ށD:�م%��m�B����z>�~���CR����|P�֐���y����n=\���J�2�JE&a��g��o �6c�`�4-f��Ê\��I�<7*�)��#��-�طm@<�l�Y��p��(�O,��s��)Nۍ&!gq+���]��pBh��t�;��>��f���b���`$�,�k��:�Ӏ��?�`q�
Ҍ�x,�|.#�dܹe=6u�Í���Z�pȧc�Z�R,�R�([1�t99����2%yl
��,��Fn��D�c�(�F���j��%�-Z;�)������X�M�5}�I�,�F�r	c^��F��N�_���=X�ւ--FT
bɄȧ
�<���P�Z"���d!�Mxlu��/	�s;rngRi,/3���fRɜH�n����4������d��sa��p��G� �BIDJ���g-�4���/�r��lK4��ccks$���N�v�i"�4��H�����3>�FGg�=������R�8qM�2@�G�@t�r3T�E΢���wpuxL|K��/�����4�a��}�� ^~��q��q�݇��}Z�^�J���:�.N�:�T6�C��'>�	X���p?���8��i>0ȕ�_��gg��≧~���/"K�\*�������>�Q�ݻO6�\Z\�:��|����ѷś�&q�gJ2)��u�����&7�fG�]��k����
0"�O"_�Cg�#�ꅯ�������EE�ae���ѐ���PD8�ܮ���
G�v����m�O������_�"�%Y�!���D0�Z��p���sF�aҌ�f��*�J�K�����E�Ջ�ז�Ϳ�1�9>���a�:œ��q؀����GC@�BSqv�������?����c*����#?{���=���u�Uy�M��Ղu|��b��~��<����^��J�P�ٝ��u����ۺ��_���	<p�0vm�3�d��ë\Y*&�kfܜ��wƤ!�ٚd
���v��'��5<GU�5|�Q߀�mA=�Dry���K�d�P˭BWM�VL�a�?0��|�#صg�|���E�R��&/��;�������h,,yp�!��#/�B!'�,���H�adl�O���p�ho	!����K��;�J�;(*h�I� \��/���^9�d�"aXd[�$s�Ύ��~ ����JW�'h���,��\���4 ��x\q��q�����ͣp��!P8��͠��E�ʉ���ZC�A�j0zT3�j�V'�fv땊�4x���چ;z ��J����Cƴ�=�E�()����5�c8��ʍY�~Z���=܄����fIN�ԋ���."��\	�ဠd�[C�,�т�Dg/�alv��Uѣ�I��|C_���,�8M��S2�p����x��SH��"��p{|� p�N�k:�c�Ⱥ�[eZ�I���@�R���<Fǧ�L��4_)��q0��n����֩$[`�;E �ڱa;qQh;n_`--��Q�Zuz���F���b�*+��]���b��B��=l�Y�v�����8��-Y�mN�,�JaWGW؋ݛ�	����CF\����W�P��Z{%'�
�:��	 �w���h�"�R��ѳ8��E���~)[+-$��!PS���qMC�1ӄ��I��l��A�`�&-)Spq$ި�.�S��sW0��"[��c�z��� f6�`ԕE;y+�S��DΆ���tf��m��k�&��QR{O����(`bN�[�s�����B�lTQ,�t�s�iԨ�%�dC�a�:d��8բ��K�'q��$*��fu��D�Q.ee�?��C��=Z�������0|^�55�0���l� ��T19����8T�j�BAҐ�U�-:��$f���F~��H����*�]�"�M4�W�fT�\S+(�3p��R���Aw[lf�ה�4pad�{�ȇ�M~��l�iž���p�f�|1�d'�]å�3�г`q�$^�Ɯ�����DL�4����R�+��o���"|t�{��FD�-�C{�ґ�ԗ+��9]n!M�j&���.�q��5AS2����m�qh�D��^4���d��K��<2��X���n1�k����y�3K��g6颁�ba�����q&r��H_�{q-�MJ5	!7���vC �Q�$`�_X����Y���jT�4)p�k�M]Ctj-N#��*�v�Ж
��4���@���L�I�a���Kp��9�s�� �ER�fff�P��4���JB�?Y�(p�E_��)��Y�!�����!�)!U�0�k�QRDZT���x&�>�2h��2A8%#Ԃ!_V�:�[6d�"Zd0r�����ٍ��	\��B9�P؏�&�8��jÎM[���'�"��ԋqu�$.���XVp��8���'0<6-�,R�L./�n�)e��|�cl�0��W�����w�×��%����,��;'q��)���L>�<� ��/�f�/��:~��pmxTR�+�4j_����/}Aҋ���8��),��I>T�V�?Є��G��c��@�<��Kx��/���R�H5����g?�q�޻�ro}W�_@�% Ԡb%/hӺZ��[sT�=D0��0)�zL2P�ץ�A�mk�}�!�<$�g�h���
�Oz���`�zQ���[�%c��.H��'h�[�� y�Nk��6`C m)�F�B�0	i��?�3\V7�:C롯7���zO>�<�f4�^�6 tˠ�y�Tl&��G�IÎ
eh�|䑃O~哏�ׇ����&��_}���_<�]��Qm.�4Peq��J.����A|�Gv걺��o~�^��J(�A�0���G���!����qkr�uw�C:��h}5 �Ɋ�yj
�Y�����E.5�1+d�J�/u�l�	������H��=�9��ƠdW`��_G�)�-5�������؍��Rٸ�y�twvb��mp9�+jF�N��%��� �̈�v�4�*z��������Sr��ChmcrlW/^���}�܍�N�h�u��
ΜƯ�y�.�`%��7�O����h�k����0�ܘD<Q�8����/)=��U#֪q�4�x�R'��NQ�X�buz
j,!��$���,�i�&I�]�ZC �f>��i��7�D�Id�I�
�����{�!0�(4(2 ��;�r�/r�\hI�$�[�Va�D�@Dhg$�f�K~֚�.r�sK�|�V����;�zDjR�2���?we�t&/���,�t�=���qKک����!�C���W���A8ҁ��.�47�,��,�TY2�Ը�"��4�F�L���ctlF�����*�V=�A6�wJ�H�47D�����]Ǜ�OI��?�"�vJ��^�5�u�����P�W�p��A`��|^A��ex8������hAs��ф��e��Ob|��h�C֞�d�uu�����z�N
y"dPl�0����%)�t�:�z[�0�ĺ� 4�JCjE:���%}�jz;\L��4 �4�Ya��`!%�D�O&��JI|=\�:mF��6�����D�ߡ5A:�� jUZP(*�[����2V�I�9�=N��c}o����*���u������	�.fDUoԐˮ �d��wlA_���g#G~<Q��xWe*    IDAT�1��C5R�g�{��JN��a/tL"�qWH/��U.�����عm=�������[Ņk��y�@Q�6�mF�i�U���)��x0m۽FIF2������!��0	#{jv�G��Ӣ7{��9P&����zE6TNka�Mr�m@k��tK+)�Z����i���03��G�d.���*�^-���B{3ַEZ�vpU�G��������NH�:'�0����Chi��f�ߌL��c�.�&*UPaq��Pe�� !�N��Uy]��qᔸ"���6�߸�DT<_,"٨����َu��h�8�����A��BCW��!sV�l�Nn-6���S2�6!|���}[���C5��D�T���WnJC��q�i���b�I�+,>����"d�k��Kb��k���E~�,d9��3FH6U-���?�D�5,�y~ަ��t�C �7����7ZCE�����Z�F٥q��'0��X�y&ݯ�� �"��
�DA_ �]�v�}�F����{�5���sB���l�P_��w�bQ��Ή��Ɓ�ΈD.���Uԩ�2X��$���96/,f�bCj����|��->;j�,��P�yfp[Dꐃዒՠ�9��I�L��,��3�u�y\�aj��� �L!�� �N������8���	{�m�̎�l3�㵣V/��=�;v����	��f@B��3'�l���42�"&f����g/��T7����d������p�TH¢/�s�>�ǎ�'��g�*~�ۗj�����\��#�8��q���jlI��x�A|����v7~��/��s�����H�wQ��?����"ҙ~�̳xᥗQ̕Qa<�Zm���o�<��cطo�3���8v��z�)\�~]���C�җ����ӈ��i\��+�����%�I
ҕ o��]��Z��m����cA���|���|n3����6w��$ UkXgh?M��4���"a�}R�x������L�:7Ԣs�4��f�Ѐޠ��;u�L-F6��Q5!艠-4��o�x_�ۧ��Z�����mpka�N�	Tl�Mk�BI$�qv��|�˟����`�������g/����b�r��Z�/�ػk#���p��5�NNb�ƍ��G���N1t��c�t�:����+7G�/a`h ����ap#����`��}��g�v�N[L��UF�HZ�#�Zpu|o���|�
�3�1i4635���"��������� �"��3dE)�Qͬ �(�Js��4}:Tdr��F�� �{�^�{�]���2� a�r!��9U�f���!�!��\��x"!�/�f��a5;$`��9�/�N��]�����AM�¢d��y �}�.�v�DL�ȉ��O����\3�������"U�!�փ����c�֊�kD���/�#�����b4����\��O��n��y��e �jEi�����^�f����<b��$C�ܖ)�y״�lD�G�h1/��C�q��5�$#�՚�����!N4��h)��\M�I�#'g���:t�i�i��~���4�����Wp��9	�9x�4�L\)��'�-`|fc31����z�se���lj7���a��n!�XL��K,x�]��KWoHb���Co��!�:�bx��Ve���U��&F�����E*[����b��*J۷`��-"u��,�a���\�"�Q������U.�H!"]!�Oc�P�mְ݀]R�W���@u��p��u)�ns�y&��V�Hwu��f�Z ���gf1<>��ŘH`8���rh�qp���v�`�!��a|~��I�F��pꭖ�n®�}��l��a���hr�	���x��5dJX�~�1Q��TX3@j3M)�!�R��$2,�lx���pXL��]p��p8��;��@a4�Ɇb�&!X��X��9⮗��ƞ����T��崊�ct:�g�ca� ��J���upϡ����S�g@,���r�n�`5�ȶ�����=vA�R��τR5��UjZ��1LJ.��Adm�7���)[���U�<���(���80��:�~5�%�5�>��>(�o���E�V���� ��&��AscI�r&_��+7$8+���I��ʷ�%y�6`S�m�Eo�咦�^YI���IA�V������6���̔Y��MǱ��w�؂���I��ɩ�cs�x��i\�X���l3�&�4�X�;7���X-:�N��|GO��|4W��S&oܼ�P���BslNB���[׉��v��dB�*�ͫ�#hf��^��l��Gw((Ġb1��Mj�M09<Hd�ȗ��'��62)�ybt��~;܁��I��T1 S�E���lL��-nz���>]��A�T�\ �e)`Y��%	����L�e&�� �����4]�1A�� 0�hc�[iX�8��ɴTy��<�vH'�R�bת��U��%��8�+�(��V+hr��� ���P�U��U.+�)j0Ԍ�W�#;6�����w�!�][7bۆ��{��Ƥ�#���J*��3Ө[�*:,��"��ٹ�ヽ!�*RrZB<O����Bgw���&F.c��)Xem�@ο�+)1Ƭ�P��q���?@� �"�ŎhYA�4�jYd��o�c1�7܌��կ�����N�=��q��qXFX�FDZ[p`�l܈�p,F���VG�vZ�K�!(ab~���O�։p�[�o�'��Ãl:���q�%��
����h4jx��w��K�,6lَޞ.��/b��M�,. �\�R�`߁�x��'�7Z�~�_?��旅t����~᳟Ɨ��EdK��?��G�B1W��&�k"��?�ٵ����{�l����ַ����>�u��ԧ>�{����,��$�Vnaai�rV���R�lV�V�5nc-@;��AR��4�T/pj��'�qY�Q˯�h� ƭ���
�+<vE� �5����	�F���V�p~��� ;B(�k�P/9��֞��F�3ə+��/�^_D��aC�^DgJ��7�׎^E]���n:JY��}54dpɟӠ�I8�Zɠ�Z(?�ȝO|����i����=?��K�.���;ڠ3Q�a�G>����^x�E��������'?�!�`/Z���ҨR\���b�<p�A��<��[J�޻���A�|:�6ԉ�\;��	M��=��^C��7ɴ�:\-�Pk�v��r�@,�rX8r:̂�4	ư��Pz`V
(�o��^D��(�'�������V��䰣���'����< n'�<y�������s���%��7F���o���������dZK�t9PQ�_Y�j4*ɪ��I�7-�+��6˴cqi�8��GO���<�Ul�f��r}�7a��]0:}2垚[AMg����x�2������z���D=��Y���t�Eo� �����WQ_^�W4�Q�7�ZK-��V^+eN����pǃ�kA��|��vX2@�����^C`P(��x�Z����b}_����f�*����8m&d�u������;W��5B
�ɹ���
��H���������`]7C�X�8��������|i9�D*'>���>t47��)�^'I��	���)�K+1�����*�5�LmN���"1:v�vo���"ԤG2Z@*_�U����C:����-X�e�4!����1c��,и���bu��a�23՚�����m^���mp� c�S����)�y��E�Z��4��`w�{?���b)VXM�02=��sX�qC�09�z�-^��>�u�A�Ͱl�������x��e)�ހ&"��v��b�B�i>�xa�/�f,&+��<�p8A��%Xmӄr1+�xCt&!pXm��r�O�xk�;��앇�;�Ã��,�=}���"�@�R1�u�~�s����ü�T����E\�:��x	f�z�*?��P6�����1/F�ə\�2�|�*�D�ɈJ6.�����:)��Aob���R4�Sg��}n�d�N�u�b�f(�����m"_	5��T*ȧ��&㰚M�[����^c�K"s��
����*�!�5�Px�p��4Ў=�7 �Z���8C�N_��|f[ v�_��F�u]�J�ز�6n�ց>D�v�wч�̅������Dav4���Z,*������;�wkg;�cL�>q�"�o��h��hq��=W�m�#�ZA1EK��{�> �n'��: ����gp��E���8CD�֡!l������*t�����(���\�[����y)�MF��"�~�s���`uaJ��ͭ��8u���b8Y��Ch��Pt&1�k��<�k��K�d3�hkFGG�Hʦf�1��(?#	a�ru��5l<D&����FdN����L��X�	�H|Z%2���L)�j��i,��]Eq�t�$,,Y+#[*#Wִ�e	��&�,$��ߍ�®��11|��铰�뎽h���%�&O�nu����|"��K������f��!`Cύ<e��|����;=}w�q@R�o^>��ѳ�-��9�YBU�m%�פ��P�A�]�2���A�T+� R�%n#�ʊ��#�������׾���N�`\���7�b~iZ��`�	�6n���m���C0�f	��JPaz�J�B�|����_��Is��&yR�N�[�����g?�>���1���N�;?�1b94�u���Oe�YI �����I|���η��т_<�~��066!�S�z�M:|����t
?��S8v�42)n��y<P+���{������n����w�7XZY�y?��.8�F��sP@	p�RK�E��W�H'�/���s�cEMGJd	����0�V=2�l�6d=p�3��/@	1�^�2����NiYK�L(h
H�U��D��h�1���B �$�&��+���F����vj6�1#��m�{԰���@�v�y���o�?��Q��F�-n(�f��R\��󆀞�j��b�C���W>s��`��������ٳ߿5��>��ٍ��G��o}�{x�wG��7a]O'؉��v�]b�
�]�B4jF4�Ə�4�9<���~`PX�&���PL�:��5�x���l`i�a-�Q�Uu�CR���$�I�bQ{�B�VT>�Jv�~7)4U�D�ƲL>fǯa��48E�(]:-�ڵ��>���$^|�E����b���C����;q�}���r���w���c���hk�ȃ����N~��5�D&!���6��^U��eF~:�%��F����M�FT��W4�xL1ٰ�ni
��{s�
U6��S
;���YX3��͔ɪ��f��>��L)�P�I}��*&�_��J}u�m���������5�5�4�1��C"4U��`���)�P�\�W���#�ݚɕ�T�e*�'ΰ ���k� %=m���h�8����DF�	|4���|%��"t���(&oŐf�Q�꤀tX�����+yD�.��@OW���4C����f�X^��������!�^>N��ʠ&J{FL�.bv�dRLNXln(��T��`p���mEW�I&K�XU�i�M�g/������J\�P���mX^]�j�����ZqTfHW]��79��>�4[f�*䟽���uc ���r:)h��LV+�'�q��,�&� �44���؉�f�a�+We�2<qK���:i
F�x����D[�~]�lt�Q�)��ur���|� �!MB��q
�BF[k�D6���R�eBKEW$ѵ�w֨I�*`��d�\���u�&N��}]a�t�ć���Q�\�>���/ciyU���K�4Љ��6��9 ��b��J���Gp��)6.��X�
��ހ={���-�T��	�~�,n-Ť�qح(���j�����l��9T� Y$����qsbN<DLj�ё��)�tj-�.l۰m��}��[/�`ZK��a��X�I3p��5)���&�%��bF-3D�Q��m��C��l��e�89=��g�bx���^�/*�JI4�j�&��}۶��퀩Q��b�pĺ����$�<yc��pxCp9=(�pJ�����]��a��^@i1bnq	箌��M��8`��&ic��𺥡�R��g>ý�����/�Z^cD�}�4%�v�����҂��6��0�k��`&S���FFnAU9Qf�Kdz����l®��2��p��9,��Wf���3�_M��jt�{͆@t�hC�V3q��nۺ���XX.��눧3b�%���z}�\�7�L�g���[�n�I�X����U :i���<�}Fm�I�^��U�Of'`(&�_�A%����_SAe�R^K/�P��P�eii���z�A�ޱs��x�g?F!þ�[1��'^'N���l��ï3=���xK�,R�:bI,F�"1������u���j�"��-�v n���J���j���) [=_��t�X��T咖��T`3}'D^+
J'�5�RY��+�c����������8x�a�s\�.T��x�	c���Է	�P|,z��q�3LA.G<��P�B�82����BEo��D���r4)�j�����9���gç>�0��{�wx�����/��(
�<X�4*TJIɤ������׿.r�g�{�z�\^-���b��~���g���
�����ɳ�V5�����<���A1C����0>�ǰw�.��N��g�����G>�A���b~qzSu�;TmT�Χ1���X2&$���6؝v��E��::�[�)(�2��j���\ߒ�I?$��!n��<n-V��>�u�\�uŢ?��%��������e�p�()�uɦbc-�m��-׃�~ �׌�y�4�ZF���ܰ�c���e3:}���~���Ë�,fkB]1�nk��9��D�?��v6�J���<�o>��PC�w����|anu����{6��C�`��ܚYē?��h�9�t{����۷`]{��:e��v�5�?XU�I���1<x�Cضu�pQ��`�K>+5d��ks�!X�ՠ��a�:u7%Al�uB��g��d���2�J�Rf]^���R@l~��W��.��]� )GE�T�]�cϞ=B�x��$��\t⩜.��hq{���u�N�!1Hi���$y]��@�E��N�8�1B�J,�/cnn���+&'���bs�l���E��#��%ŀ��n�"�Pu4ff��$��h����5w�L��{h)���ee�V(1��m�IB����Go��{��=Բ�!�2�ְ��/ɐ���M��G�����.�)mp�n�{�~8#���!�M�5 5���I
0�>6�M���"��bY�֐ݭa�\vX�u	�bAϭob�ix}q@z%>�(dnW&gWK�`i��ϔp1�O�e�6��ٌ����8�6���xH���� ����|M�� ؈�3�Pd��^*��j"��xV�D�$q�Թ�l�`<���͂��0ښC��&ʔ�}��h�e�L�P)���у`ЇD*��6�� )�8="�J$�x��Y̯�`q�œCJ��QX��]X�.�� c�\O�:4����9:� &R2���5$�}��r�IܜZ���tV���s[H�#����6��+ ���Na�p���Q���E�F�A�Y*�e$hi������RR���
�D�y��/ѳ� ���-�j4���B:�g�l5x�z�v��܊`�.Iz�|n,G�8u�<.^�������9�����d�(���N]����8Q����ۣ���[�s{��ADS�_��q��0N_��L6'�M.�n���v�א5����?���(����RQD�H]�A�K�]zl�Fo�E�T4�qJ���9���<�=���	Asz0�d�V4��%Swkt���sK?z;�0�j(W��Z���ØY��h��$[_��2�>'z{:�*�
�N��Z^WA50�����c|.��P���,��ɨp6�w����r��F�����1�F�y���f�S��l�>�Ⱥ:Z����})YE&+�&�p��,�R�0��0�$lV4�U�i�SS��N&]�R7�j��V��	���bN��a'�o�BogMO�    IDAT^���;3�ɳ�F�.�`sd����1���I��E4�Y�fw�ڍ;��,���g%��Ave��IksJ��	���Lf1s�*�����Ќהn��]�Ezy��֝A���ʆ�ii�m�CI/ˆ@�ĥ!��V�tȗK"������
Ƶ9ģx���عu��c���?�č�������P��ܪh��0lr~�	dj
��ӋQ��.�LS��JU2b�	������!R�R����h������x��`�J�<U�ehztI�e(b�($*��
�7�\��مE\�>��7obfyV���o���=�L����I��|
��G��F�=��{�b��6!�x�>��6�I��t[U���$�T��k����������P.�٠��X,�dH-e���/��s�����Ͽ�_��e��>TUn�̣�cM���R�j�|��}���7����o^�/��-n����:]��bƟ��?ŧ�����Q�Rr����jE���U��R������%�r%���v`���h�'���/��ʧP��Q���$e0�{����(P�>Z�P�U$R1ijl�׈[��Y���b\�[E��L���!n'S�}2l%Q�>�/ZBa|>4�(�M��.M��O(���YN�iݠ�&�l��ƾ�fH���I���1���ч6�l��iބN��x� 0@Ͽ�����b�~8/*Uf��$��V6�A����ɮPL/��<����|����!������^;��R��im���߉?z� ���<I%7nB�7�j��Jӎ	�`]m\�:� ��TK�k ����ś��^@�ߌ����u� �jU��t�� [�����P���,�i��d���u�!�;�S5���s)Y�3��^��j-z�L�l�P�%��8���"�2��60z�HD��Er�A�/�Jo��,Hx�6������Q&�5񿩩Z(/:Ѭ��!��)�Q<�6�ml�;�����DĘ>#�:�� ӻ�j�#�!I���D:DD5�<,]M��<�Vƒ��N����5�$�Tu�0p�c� �Lcuq˳3Pb�����=ɐȿ�yQ4�(���ZL�x�^��0,!?��"
|����	W�Eqa���u_%c�r$�Æ�`���$=�M�niɅ�I�A60�(�ilt�*5A%.ǳ�ƙ[A4�󟞅���D*0rMHҒZ��iA$��;� <|X ��F�rr�@d�r��A�3��R�WO&QS���r�0l+[�����k�l@0�/M�N�	�z�%Ԍ�}��xQ�J�d
�L��P3����/_-������N_�]��o�uK�,~��H�1�\̠Z�	6���3kk( 2lJ��x��,�y��ӆ�21�����k��ZH
z�� ��+���f��X�H���"Lz��]*5������y�$ƍ�C�O��N*�ľ�Y��M��S���#DݴA�5 r��|��8	.�BB���{HJ��i�,�>���U��H�	f(dK�%������[���GxƵj5��\�*pk9!Z�T���'dM�#���C۱cKj����`P+n-�p��y�--�������a]W�'QU�V��[���k��R���l.��E��Ȇ؀��m �����ކ&za8��iF;�a�bY����8{i�*?#l6�ݥ�)9��ө�����&�$��js��\�1%�3����y�tvE�u�F��#�J#����M
�?�b�0<�h�o�U"�^A5�Ǒ�݅pЍL*
�ہ\���XR��<�LF|MAēix��D�m�zir�٤\#6��r���1<6��ފ*osru(q� ��mSI&�f�ր�I冉�%����[	���+�<��:,ܾ���׌;lG��%N��������\z�K08Q��~!��3�����bۮ=b�>w�*���ّ���Ĕ_��rI�-�)�v��v���L����L�g�4
ZF����<W�i��]��e�+�rl��`���Rl���[j��%i*���W���G?��~�#X�ہDto��"�&G1�ӎ};v�mwh0R|֊s�&r9�zT���f���-XZZB<��;�����Q/d���Bkg��
f�'P+���ej��i��,>9n�%qV�Zh7.y�t�a�a��P�V%�����q��y�����k��v<�ÌD&�w�ǋ��K���������@���*�)u�^HG�f$	1ٛ�.��~�s����g0���j!�Ɖ��A)WB��F{Њ����>��$Y}�~���`%]F:_B)S亁^�%�ri!�������o���^����J��%X�ZC���>��D���Sx��S�-����l�Zn�j(Y/�6U��F�ۿG}����,`�V �d~K47�rh�A��_��-GC� �:[`u�-�a��V�e��I����C7!Hմk�9<����Fx]n�<�B���d^_M.�N�ȅ�����-�����JA� 2J�(i���5�����3�:�o��KJ��d�S,p���ڀ��8sz
��o~��9nH]�����2����\������)�T<r��'��˟������	��_ki���211a�_�|���\�+�����������E��:�0)��ڧgՊ<����,<�v#�mb|���sϭ �)J�#����QJt�#F;
������Y�؜�5ê����W��!�Z �/���"2L����RD����C)��B�h�ULܸ����~��F��
�v�)M"�_�� ��&T�L��ɦ�]/C�Jfh89a�ՁwmK����f��)�,<��D����U�X��8'/�2`s�� Y�PK�F�$gs�#���QB�Dg �_#���g��bQ*o͸,���Z~�WT��]�!1?���P/��/�h7��bN�9!�x|�sڱ��>�8|t^V�y�(Z�Ь2��S(��9�G,�J�	Wn4☌2��V V���Do���.�	�r���Ax�L'ҹ��a�$
�\��|T��Ē� ޔN�@6�U�ߨ��PUbwb����2�߄;����˚(�5��FCb��%�r��{�S�t�(M��bL�Œ":h��O��bѕe�l�@������D�"2�d2!��j��	=.�
) 
��"I	3���8VSYxB��9���,j�4�J��o�6lܲ~�z��I1��بq���6 N���f���㝓�MW`uQl5�?C����[7u�����rb�BY'\��7����㚱�4�
=E�Z�߻��FLT�tr��;Ԕj1�Zc���?�QWE��V���L�Ђ�T��7�u�*yX�5�6c���t����\B�^-<b���!/>��&�l5c5U�)���Fg���aF �'��$3o�Ѝ�C=���(f�rM�+
�FfW��e%���5,�7&���N��.�,6�5����^��$Bs%N�4�>�m�䷷��a��\m�c�Faܗ�����3W02qWL6��e�	2_/�WnpQ�JQ�����M5I]��5���fB*����"��q����E�3��|]F����쉷�Fbvi	7'g1��F"���h�n�eb�*�"\��ܻC��s(Vs��aѦ�Hk��y��3E��_k����$9�����p{�҄S
6���� �)��O��P�$�D�I�yC�ٮQM`Ҷ7"a�GP���8��p����l�I~W�4���=3����y�/ŰMJ�¿�v�%�v��.��TJ�
��0�{|��%"=}(2[�������4;m�d�5b�ךh�9�`�πSv��T��VihR	���
�sN%�&wC-�jb�Z�*�	�2iJE)�\�	�%��0&��c��G���=�t�.�}�t;6mD{W�l|Q�s�f�g�P�4P��*7͕��(2��q��2��|���(�cHD���BC��Q�'`pjC5�s �5ɉ���&���=�Ao�����yx��//���x�7�֩S�_��lݳv��F'Ν�ӿ�)斦io��m[�~6�5A���	ה'����1��09��:�����\��bt�������w�����?�>���(��x���/~��Ÿ��T��ެrKdD��D�Vl���ݍ@�	ӷ�$D���ⳌF������'����|�&�s/��e���X�h�\�(�m?��@>�Dk[�~��8|x�x(r��N��,��0�0+y:��Z8��fu� �u�IN�R0*P�*��5�$N6�Ź����/)bZuI���M������s�.��nc7k�ɬ���i��ÊJwI���^K�1���R��[�p�G;�!�����W���h����y._Z��~���dP�[G�O�wX�C��635�ej9�jf���G=�������93��_�|�?��6�eWS��)���|���.��N�u�u�C�s1���|�zK�*�����UBH��X]����4�͓�;���0�6nl>��_���(�v�^��'A"ٵA��P �<��R�����e3��<״�\�il�*v��<���0#[���U��E!]kxJ���hw��-:��pK�$`N��C�U�.��0��L��e�bܲ�Hf1Ia�Ɓ�����X)��r=� ]*A1���B��FX�!��4�5P,�u0��|�đ�� ِ�@�iDr!+b>��n�Ĉc����$�,����4��*���ↀ�71d�/��g�φ�Jɐń��ޅ=��i�b&�^C $��V���b!(��rzY����Y'r�֨�<������j�C=��w�Jpv�8�"��X��ϔ�A(zon|$���̆I�Z�m@I#�k�UT�s��u;	�7����b�B��,v�3��Z�t���vx�MBhᦢTQ�!��Y@2�	�V^L6OW�,Mt$��=(��qM�׮i`�VN+��ɔ!�6d�y�W�XM�̂��D�TC�\��K?
ѳ�_�aP�b�f7�i�f��ȯ�P�����N�[��Đ�OI���L�(����s�(v�m>(Fʣ�0�*�$��,����ÏP�)��U��a�RҖr�2�6����E˼#b��υ�x$����IC�Y�A�\�]^H?��tF�����4W("�a��}�!�9]r�i%z�&�z�)Ud��m�ӋE\�9���UD�UPI��}L�IMp��)2�a˺v���1��V���CMBӌ(I�jȔ�[/�ՁZ̀��e\�8�h��M���ԙ�K]8e2�����w���;vnD�$3�.J-U�(��z�_�1��O]����b���y&[s"����M�ZEKЍM�:���e�	��Ny��$��%�%4�Y�Y�~���f�H�v�{|�U+��gg163�h����U�F�	�LE-f`�)0�d}W�q]�n��eF6�o%>&	�
@O$-�������@ZH�D\66ަ����L�5_�V�l�x�ː�c�͙�+�u]�Ǆ���\U�Ar��g8�����|���9BFڴ~\V�H�L̝ ��`�b4���[��mIx-�l�GO'|^R�*�p�0='6X�>�pQjDj��x����$��g�������ֆS�]��������`H97Bl�J��L�l�2J�u��(�����(�,6��L�T��0>�����AoG��".�9�z6�ݛ7���]�F*'���|V�9��G�PC����̒��׌6$�E��)�<voۀ�����쪮E���ԩ;�A $$� ��c�ql���66����k����d2"#I		P��[�թr�:9�{ǘkW|����]���Vuu�9{��֜c�p��T�do:��L�7R��  YZK��s��:mrCR��	#]x_�F����W�P��q��Q|���߹�C�����Ძ�]�ܨ��G��}�,�.bp�[��(a��[020�T$)��R���	���L4�Ӌ%|��w�އ�֡aA�j��N�ky�@o��W��/��R���W��o��K9�;�k�e'�gֹ�vMZ4�htw��.��߇��U�K��V�Z�/��f�|�-b#0����A1ϳ�붮5�)!'�y�!�3�+y\|�y��׼����%k�Ad�8>��O�@�����|�`(�3��Zڷo�2�={w��R�!�,PC����|�h�k&#�4d���@\��sH��Q;	���i�` $Bܐ%k"N@�l5z�2���7�&�V@�C���Ջ�R(��U2�f;�p�����;r!�?1�~�N>��Mt�M�7��@83��!�3����6/�w�'��G/������_?!���]�~�����Gސؒ�"$����p�۱{� :��Ɗ��G�&�	4C���A2-_��]����J+�yZ�����S~�/�EPjt�&1�P�7��}r
ɞ��$m������~�Pov���刔�cفM��(���?�Qi�PЋ��E�S�@O=�8ٽ8���p��C��~S���LB�� �(~�|0."��Av�1-�@4�y�6c�	7���\|������rŒ�C��ڦD�@��Cr�c;v!38�XW/���
�z�>G�I�|.�Z��B������Ի���*�T�&PxJ�f܋3s��� �"��&oB`\�_�X���KطC��a�.~=�+^Rp�����3_xZ�����PD�)
p��(�@�/{_@c<b�ۓX��5D��þ�"d���16ҏ/:W���0��E��3_�0���Z�nD�wEQ�������Э%� �`)k�JǑJ�{�A�\A�X��ڊ�;�;w�ęg�EWO��C6LDeNOLcjfAM�m~�RB�B���""VXy��7����ү����,�2�^,,�`e��we4k>��O�B'B�vn
z��kiR�j��4�{I��א�Ǳg����+ǂN<�T�uK�əe��A���Bj����c�0���4�ڹ�[��k]�+UL�,�#��T����E��,#�a�#��R*U���1�C�T��/��@)���D�n�� �0kN*���fӏj���"eӞG�^P�pO<�g_v9�{���RXJQ>kR��#�Vs�c���CǰRn(��k��'�PX\�Р�����Ͻ�
��1�[������P�D�H�v�@Z��ࡇ������
�z��P�h>��uk�;5��5�K/>]]�9�i�K�y��u���_���;4�H��F��Me��sE��Q��h[Fp�Y;d����T_�5�$�����%,��o�v$�|��l�j5DB$#)q��V��8��i�+���_�!�U�p��SA����0�ҡ\͕�:�̈́CZ��>�حTY�
�W�@��o�|��P����#���c*�c�^�q��4���=�9��x�Iu��}����s�#��Ѻ��"��G"TÖ�.��<$��K�twi��5�c%�Q��Z>��:`���'w����C��+��� U�Z�>M�Ho��uDg1;l¸g�[feK~<�9�����BH�yDku�=˚�H�`ڬ�Y�}r�]Ai�:�UĚe4
9��(�ٔ+�D|�r��
j۲m���|\��8c׈�~����,��½{q����Vf0}zB��&�g�&g�Pj�����q��Ќ�����0�}p�1\r�^\t�ػm��RFR�.Q*[�U4�g������3�v�h_�Ã�d�4����!����R3>9�o��'���~��-;��{\��g�P� _.�!�Ɲ_A����X?��8��@?{�0�?�L<�&�������/�F ��sE|�_���=�N�[9 ̋a�º���T��	�+_�䖗�}_�򝘚]V�&���I�b)T�uQ��8��u��tR��k�V�!�I;�w�^�ܹ[F�'籸X��bAZ:4�p�N�>j���c~a
O{����7�{�؂���X�. � �m�����iT�M�Lt�sV(�4�Ʈ�����-��uPiW�,���,=R���F�D؇0�L�f��ŹC�e"20�$iOʏյ5MX�|p�%l���lX�(L��"
p*��It%NФ?h*E���$x�=;    IDAT3�:5}�m8c�%x��)|�cw��x�e�hE����KVWc��ۄ�݄ ?_��W<�S�����s���X����~+���G�����n���ߘK%�{����W4�>&F(��(��hIK	������������ف[^�<�{~q�/�����Ϻ�[��{?y����|�Zl�s_�NLUˌ�IX��dKH��8�<��8�M#ZCݪ��*XTJ`j��5ڶM���V)���X$��t�v���ǱCG����y��˔/S�k�1܋�5zM�P�F3D�h������0�m��1Ca4��+1W�z�b�lX��G�=<��;���G����_�-���Ew����4��lz���r�j�,�Q��ksGB�N�	M:G�T���;uX^�	������Dym�]��#:�O<Z�����'P(�m.�'��|ޛ��b���y6�}�-���EI�^��^&�1��)W�FSv����D�D���(�������P��<����B%X�s�P��Hui]S�G����7����U,D�8Z�JKs�aAkF
��l��[���^��E��7���k)���_b����M1�+�h��S��曜h�tO��bll�#C���R�>M�����F .���CKU����)_�	^(��,�x������a�B��n��-�H&�[>77���YM\����
63���#h���,���<Ъ�ZE�<�yJ��29N����&u2�H\�;�� =����k��`����Xo�m��5��e,��\$�޹>[�?{PIǺ�������r+�4HD����e����޴@���ݦo��jk��C/�@4��?Lڮ����^ɪ@ٳ}W\r���%"Sh�Ȥ�Zi��bl���p��Je�ϸ4.��^���,��Ry�誔�N ��;���~��!���!�23Wŝ��f旐���i3\�����&`A?�&y�J����at���*рhr�!��I��5��I���g�S�B�M���)<��I	@��(ڝ r�
�nd�4�j�����zi�����k��3w����`d$f،��fgW�i�Po!ݝԳ��k(C"�����I84�t�H4� ��~��X�9��Ŵp�=Q�ׯ}�ɵw�ʖycM�B����I1�*�|t�;��b�����E�0g��dJK\���}��KE���q�}HT�'Q���	��
��h��'�v6�4-��g��T��:�''\+z��y��r�����D 5'Qq#���⌄�܏4����!���0/*���nz��x��W#��QX�S���O�/���lIw����J.���0`z���v�tE;vG&'Q#���Ș����d#�]8o�V�F����mx�}�q?�&Q+��E��P��|����ए{��9�ǰ`FcPߐH��\��%|���G�x�.���3�?�J	��xt����]_���i�{�Yؾ��#���8��$Z�G�F
F���7��?�Ǟ�­�~r�~b��,l�)�6�KS�>�����<�9W������{���;����U*t�4ې}R#E���HS���t
�v�/hw*���)܍�s���hu���W��k����J�!N�S���i<��k�xF�����a,���i��)bfi�(C�"	s��ҠK�R���k۶1�¼�YMF�4I��3ò�H�V���[�xJFV��c2q"�fneiYuid�D��>�,v~��E�0s�se��:�?��Ʊ:�V��݈`2!%֝�~2͛�>JR��X�}��8s��x��Sx߿'OP���K9�$��R����_�Sɦ���k��W��E���W��^}v��o�l��ߺ!���̻�?x��C��/��#8��~�L̠;��8��,!ߪ��fD�NA���l5+���n�
��W��[��_��6�+.��#;Qo0��iߐg�F��C#���d���>L�5�ي@4m�nr���ۑ@�OT����ʃ��,u87[Y��jS�j�R��A�� &���o�0:FW(e�8r� �<���(4�U�FQ|7n DU��|�8�Q.zң���+VE{a��!E��0gdr�;@���!l=��lA ����
�W�*��Lҟ���ܺe���Wy&��V���g�!�5�k`�į��8���	��-D�����)̟:���,|�\�\u~7K*�]�����j�f��ˣ�G�Qv�D�̵�<M.H^��(��q����Y/|��S��(�\H�����vGw��R��L��ZMt+�Ѷ�vݎ���Ƚ�겙 ���������MFu�
��	?x}i�G��l��_�͠�
xE(@$B�9�$�;��<�nb�#�(�C#�~�a��Ƈ�M��!*�ü���9΂���������'�Tʇ�l�؏ɩY�3�Ʋ!3��o}��b���Z��J���,{5>W~Dšg���KMEV.�S�`���#�8�3JNKI�~J5��$"A��t���p���ȗ+B�#Q�s*���^�{kٳo��z��oBn�zIk�~�΢T�+�s��Y
�/d�G�ߓ��F}��z�euH���+zݬ�ff0;��r<���V�

>l�]�i��B�{4J��v��
��Q H�b�Q'����c�g���&��lie�E�tsb8�z��Sۉ>1M�<�$���F14Ч"�rww7��'~�q�i�b����	�[]7ڮF¦C��)ãx��!�am�aRM�kei�R	
񍖢�,z|���p�z�\�s�X\^��V(��Xh�k���B*�h�L��P?
���%z�Uc�������4]]=�Jw�ȣ��t8"��(p��
���abzQ���$��қ��� ��xM������6��g��5h��Zm�f��c#����Y�v�����RQ�O:+��\�4`���P*��G������R�%ŏ�;�?W󦡙�Ϛ�4����:s6�ux���+�I_��_�]v���޹����h�_~ťi,O�DquA�2�P@��+X0�"�F��7�`2f?�Zu�?��?���q�jUlK��5�F-�&2M�� V;>�ZXi�pbf�,OJ��tm�]�v]�r��q��b�N�@���yg�Ǝ�ў�����V�ҍ��>��/�������N̓IT�ŒXk�q|y��?����ĹO&���wa��]�����������/k�u���c��]�P����;���QW��Ъ����Gw �=�pt�sY��c_�w~� *����C	�VZ���Ǟm��m������Kw�_�&��
:C(�%r���M��e҈��₾IﬖVѕ��}��%/�'��w��>��[XY��i	m�n�)�r�kK�I{�v����<��k�淾[��bbn�jZ����;���)��@�+�`��y�����M�R��NQ��q���_�d�P��ɰw�s���5�@"F�v�� z�z�5�=tmqqݎ��#����	Hq�6z&��s-�eC@#�H(3���6Z	II�F��H �X0	3�d�Q��\��<�~�K89YD�у�?�N����݅*����r��l�y��_�ꗿ��������[5����}���u߁Coݱ��ƛ��+݋;>N<y�==��"h���*83�P ���jL���K�v�=�R��w_������]�-��ܳ/���Ս�X'��V��$����ů��+>5�D�.�
-�NZV�I�Q�������B2�Kk�RUa:��'�A$�X�Z߷V�h�50<Ѝ�L7��Nڏ���xh 
0k9��(|$7���l���7���)��nK�3(8.� 7�t�]=�����g"��'�A���J��2�1�	�É����{���R�u�z��F��դ�!��+t
l��$���Cvy	s'N"w�4���Q,�����M��E�¦�h��G�+RGQ���@�=��`�a�m�\z�5������&��a���6<Є����tX���+�y]]� 	�|�M��tB�:���X!��
G�|}� �F�R���g�]�r�,ʴ�؄IX�`9���0$��M��ZԄ����j�/�YD�y�xp�@�3V��I�D�גMU�]r2�I�#�?S5~�(f�14<f(!�$�U�5�]�&N��cG���y%NxH��R��U���p2��>lj��Tij�|�Yҟ���
+"��s���W.&V�(�^k( _��A���gh�v#^�G^'�v�mt!7p�Ŝ�|*�%�tk���x>ּ�j��T���o��m���<��6�H��֝Cq�����D��AD�)M�x��Y�r���V�̄�h�(4SR����J&tٴ�n��Q��~�����~2��b�IoBE����d����N�V*�eu+*�\�8)�h���A��Ҋ�P�:P;@��E��+�Q�$����6�G��g�V4[L�>����L:�]�v`xhH��ם�ܫJ�V��8��8N�:�`��}F����p=ЕJ�p�n�AK-�rE�n~uk�sx��/�uϾJ����8uZ[��]{1<���k�5Qz�s�����CU���U��}\�v����4\\o����o�������� ���<-:�U����;�{�,m���i�\�>�:�Y��0���O��%N��T�B�٦?$�)�nL+��C��܊�i�KQ %��x��F�ͻ�?��g��:5�|N�E5�1 \Y���8�OAiuyݵ��L��,������՝V*�u�\����Ï=���Q��@�Q�h,��d������<�/�"( �'�X����-"W��fD][��@��^Z��S8k���vcejkN�q�Ȁ��,���2���A�X�󓈧�n�ĢN#�G�֭�j�0&y�/gql5��bWߴo��D��&�p��������v��[�� !�L`��GYt:Z���$/��``p��#H����b	�����z#��w*5,�>�s��߽�Op�U�cvn���W�;���S������o�y瞍�5|���Ɖ�	��J��6��֩��K��߼�-��Y�����]?��?�q><�f3�r��)w��<�1'0���4�f5���q�M�ƛ���غ���Ǳ�:�N������)�,�e�!���^�����F'�S�F<��8�ⴈ�3C]5��Yn�����.�uL�u ���aզ�SZ[XR��6#-ȧ�1W(�P*��3Hx�I��$���sȥ|�X�u��U8��TE��-�)����!#�p�n���r<��c�Ї��S�e�Їv+!�.;g�׭7!^SN@�!������/��?��[>p����߰���[5?}���{?�xrr�5O�����_�bLO��}��>,�ߘ�^RX�����D��̍�*�d�2˂���L"$���{>����G��#���kg�9K�7����#�[�A�R@��W�� �L0݂P*#�o�]XR��.d�n�
p*�k��=�8)ЩqL��hG�~Y��S�A�T;Uu�݉��r.X�9������x}ٕYTJY���	����ǝ���,$����X(�F��G�A$ҽ�CW� ��nDI��81=�%�:�[�P�L���QX<P����m'U��Wo^6�6���)F���5Cb�S�J�=1�����5i۵�H\���F�-���6���98�{�r":�}������7\��=�F�2)�
(Ӊ�\C���!�l�q�ǃ�cwE�
[�at(+\YX��d���ȭ��C�Uԓ�E�0���II�����ݐ��/*�SE�9��J��9Nn��t9����Q�ń��p]���@2��ь�z�\�?����(�
��lB[��P�|6'��K)�t��J��?����b㵩!PQV��o��,���LN���p��b��F����p��}�z�C����M�jU�a~��E�$ø8L�U�])�D$�?K�ݽ�!�����ϙ�!`���l��@��bS�.d�RǾ���r��1��^�MMCh������W��PXNI�a�S*W�8���4Z�A�\@��s&�x"���ɉ�դ�D�Q,���6"0�M$q�^C��l*V���!�V*�xe���zPφ���f�� ���J��!�5��0
�E��{E]����r)���y���s�v\t���A�R�m�Z6���
]��g��0�"�N"���&��k0��8�2i LG�BI]$k���9&�c�<���%�����H���|aU߫X��JsqeU6�1�q����0q��W�"8����~{���͵��Ok�t#]1���'�����L2��=�v
#�P*���ī�D�����2��Di���Dj_!6���GU��ܢ���66]�M<�'f�����(���O��n��Y�̈́�
�(C}q�s�p��QZ���9����5�5ņ`yyQSXNڸ?��9���Г�a��A�?���<��1�&��Z�f�(�r�6�ҜpB�X�`�,��X�=n�fU��t�|H��K�q�9g�9�|�2]�<~sǏ��4�P��&�m��L6�	�(�j!��h��K�6����j>�D� 
`b-���U�q�K�y��=��O�Tex�y�O�Rn	�D]}�##�/ӥ �z!���U%�!��2D��3pj���}�s��g���8�����q6Z�"r�'q�����<��gcnv�ꋸ��w��=�N�%/�	���W`���8p� >���p�}��Q)��4��M7]�w���18E��ƽ������ؿ���Mu��&z�����`��F��F��*n��9x�_�[��cf���f��S�U�R\����V�e�@�fp��V|F��04؋�~Kv'�����P]Cs�.�ӝ?rVc�I�P���^�h`S�+,,�\D�&p�Kӳ3����Q�@)�*x�=��s�#�}f��Jd����C4�@,ЅLl];q���q�Ç?�U��� ��C�F�B�R�hT/M��Il�Y̡�6]x�k_��7��-��ߢ!��/���g?��f8��}��\y�ex��'�o�ފ���hJ#�D0�/�7�\��z	�=	\q����׿
go��B��{�� ��{���b���J�&��f�<5�;��fWۈ�FIuK�/��g�E�A�Ad�;�y0D������榧���hM�QdW��H*�
��Z� �'@2B<�F�W��#�@�f	�FY�`��
ْ4L��IZWN�<�3���])t��#�A�XE<�_0��M(�nw0���R�j<�5����
��ӁFug�`U�FC���졾B���-���O鐤t�rY	 �^�NG��I�i�7~N����[���J�)y�8"��J6鈎dC�bZ!����o��P���?z�"�憀c^wL2V��ߞ��C�77:���خ�E��B�beM�Dx|�u=n�0�j�jU������}�)���h>��Z7gY���7�B��p��95 ��)�������(&�*��r��i���H0��	��lb\+�t�F��_ȷ����H�`���c��H'�I�j��me}� �,�u ��P +ĕ!�Qؼv��z��dQ�5�j�_�M��D�r����5�,���r���=�b�*��G�����A������}�~�4$v��Z�+�c䡛nAt�-NmBTo�T�3���޵�O^Q)�g(ײ�ȯ��D�H!!6�	)j6��>wZ�.���{�uR)�^g2,��vm鶢��=�z|f%�5�A���Z&��G����
ͺ�N۷o��m�����氼�,���0���.{�M��0j""�k�y-��d��
�n��ygSI=Cw]S"(���>i�+M�>�Fe����g����8i�z#h����Z��P�c91,�]��@k��A���;1��(��~�|~?�S%M��A�)N�lrM`���׈�SN��E�W�Jk��/V��Yl4-��h��f��+N��Y#Q�%�('���MSb!�F�uBM�}A6%L�f^�p&��HSO>�����gA�    IDAT�"���A�R	Q�<�pf0��k�b��;��*9���]Fuy	����+@�t!	�2��I���c�PD%��|����2��F��W�Tfʢ�ר�?W *-H����..������c�S*��b��!q�9�6��\`n�")¶���<K��Eb���J��㫫�(�I�����O��z��Q?�ӳӘ^��Z��P<�toc���đ�aAH������36	!�B��6��<�S�x�Ǿ�_>z�U�<��p����4ιd7�����q!����2���_��R��܋w��_����?������|�'h�\�Ą�eUE쳮��~�;q���n���?��?�Y8p�F��x��J�}S�����"��ny��ַ�1������r�@��R����i�:�٥	����
t�wޤ�R�}�`tl#��2����t�&���n�`gO`N.�+��3�p\���3�@����`H΁j��1M
r�&gg4)�B��HI��<�7��Rꮅ��63���0��A�݉At�GћŮ��q�7���?�MLΒ؏v;�L����࡮�{S`���Gem���/{����wny��������С�|�+oٲg�?��������y|��_é��ǰR(�Az��3��}oF�FMt_���ع}ox��a�7���"� �6v��k�B���� @���0�,��=��3%�C*��<,ĩ5�@6<K��%�F)�mӬ+���֛��mሉ.�x����!'��Q�o>oRF��i+�5�Qǎ-��>6�x4$����
*%&�$2eB"���(�!2�[)��a%�����rE�䊨4Zu�}&L�k�R^E+��9&%��r(b2��1��b��w qC!UGŤs�oM�������%�Q��r4Ŕ�F3Ǐb���&�e�nN>C��{c��"N�EK��Ԓ��.��֡��RC@��,�g<�\r�5�D����5!൐�P��͙{ D!X�7�K�����¢B�̡��f��󺒲So�(�}��+ҽ`�JdFW�g>gŴU�j|<+W�oU�q-̊O5�,��TE�������\��ϯ7l"\��'���סx,��*��L[E6���Ԫ�oQ#���I��F62r��F��"�!�}���#�m��Ǎ�-��CU��#킩�F������MK����o�gs���G�5��xY�q�z����1^a�{�5�|���΍�g�+��l8oy�A�4"�<��l�5g��fg�R"���R�6����5�,,i_�&#P6	ך�� =������J��=)S�#7�QԞF�_v�ɻl���E�*�u��.�F�^�YZz}z��3�=�Q`�xoǗ�4�_�u)޹L	̉̚G�"�U��{��9~=�/�;)#ٵ5��e��|��s"��1��0�="�^�&O�/��X�aɻ\�jl�ia��Vg�YG	ȥJ�٬l�I7���'�e�{��B�B�5z�8���eMAM�l(�P�E��f�mk�>멚=��[�xI�I!�@�H���|�糺6�PTS��!���(�Kj���A]������'v��I�U�l�k.w��Mx���%n�p ��DN���׉����ԡIA|����8FR!�:��=� ���&���kNg2�^�s�j[FG�m���r1�L,��߇`���C��K(.-�������2��η*��P3ky��K�<B3	��+�H��XE_*&mƥ矋K/8O�Vav'}��e}R;�,1�L4�zC�n�_>+<#8=$�W����Qqzu㴭q鳯�஝�DX���ajn+���n��?͆���~�AQ�#о�3%E�#���щe|��_���h��h7�R>B�T�q�E���s\��˱������K��GnC)[@��1���ߌ}�����8=�O��%|��w�U���lƫ(�06ڇw��x�+n�)��s|�C��C=��Z��pW����0S��k+���,^��}x�_�	�]C�-,�m��`���8|�����Ѫ�Ź�"6Y� 	c��Ai	��ϯ
����Z��Q�%�.�-�z�l;����<��aR��QR�X�xRzR1W�VU�؄�E��w&����0�ܐ�B�^'�'�ƹsm���ۦ��CW��]��M��7�[��⋟�>��ocn�,�^�|� '5Y�p
O��3q�D��N��ja����_�����+����4����o�}�Y���HZ���	��f��̯�D�	���C
�U�HHH`�DӀ���ɎG�����64x�WM�W3AkN����>��ǗN!�;�Z����<���:I�g
.�34�!N�]q�]��_�XR��n�RN��N�I~?�����}Q F�Bک���}�N���W��d��[��eU#b�6�DW�###�?����!6�H/_z�7��ۏѱmBh(Z���P'��*�d�6�d�P���	iZը9�$LyOE�_�2��|��Fk��b�b	��:���G]0Y��f'�k�ߚ�'��ϊt�D�Xs<�]O�5�s1�
��!�������E�����I�Qf�_�e
Qr�1|�U��G� �8���D����RO�z���ib��
��i(�-�8z븷^C`�]_o���gZQ!�xt6$��R	
�q�^o���� yӤ��ζ�-�9������c����IRb��u@h��1g���<���fSs#�E��9;�h�6�F��^�Qq����t.�������9b���ʐ�����;S#a�՞Y��_)�<��  z�����(L�4k?pfq��,x^�����k��8pr�5�	{��$��n�p}y�6�l(��������1�t2�7_��rH��*ڣw�İ���0� ^G~��L��K���/��x��,��8�>,�Mxe����Х�&O���R�fM�K�鵜~Fn>	����u��O�	�]��]�M���"6�N����֦=�Ds��=7�8=	�&�!���h,([�b���oj4���p���hx�hB��/i-�Q��"�I^c�lKf.K^"��������%d�o#�A�I������!N��ӅǛR�P z���q?!�E�<!!P��"���֧�^�-g���UA�7�T�O�$�Sz���0x�)����iZhV�NE1�	a�G�x�����	��fW��<66&�%iiL���35D}y��5�ۍ8�r	}�4­���V���|��+[�H�X
��"��2�i5M��M3UQ�ɸ���x=�����8ꋫ���*U����n�
�r���\�h����?6���P0��b�TBm\����=:�R�)n{�P������!�9s�MheY�j*@`p��G5�4C� � �m;�N�㓟�:NN3�+%� �8�::Lj\[���Ļ��/p�uWb~~����/j2˽�����7��q�9{p��8>v�W��o� �]���V�}�^�����o�K�A��G������2�E���Xʄ���i�`���Tl.��5�����W�fl�1�م�ȗVI�P�����tȵ��Pa�W0�����cfG�-w��E0�C��l��,c�ܲ1Q��3O!��̀B� @ОMw����c]+ �K��X�f/Q����/3��ų��ҙ�s���q���� \<.��O�Pw��z]�s�h?�C�ڎ��.��|��o��wރ�K�9"����^�X�y���sA��k�������]��7�n߿^�s���������9�}�疛�B�!���|��V�1M�ָ���ؐ�OOx�xk먣\aQ�q���c�F�-�9kN"C� ��TB�^j��w=��O�"�Afp	Ry@��;�G.!s&	ț�I(+�r��Q������>=��o�(SAZ��Ŗ<�u�Y����Hr�Ѹvqnuژ�"(di��D(�A$f�-�zS3�ӭ�J��kD��(�VsH$�زu�>���,�[��3�5�,R-\�K^9�_���)�U�C{$�f���oX��{ra��B?�h��DŇ{X�Qm��H|��S�f�8��*�wϴG��k��A�?�l@�t��v��[���}���#�k���
��)��Q��]C�"ːP[#te�\�j��x��ZnT�!�^(�\s���G�QQ�Ę���%L��ZL������C
�I	P��cC�QsDGp\e���YA�5B2�����Y1&��RTD7�*�q�Ձ��k.A�T7)�M"�H��A8��:|�Fsה߇��Ffl��{?�H����e�!�Gi��Ī��U��P*��<k�"�Gs��L�|3���ǻf,��H�Mז�9�u�ֽǵ��s�v.�1�u#:��'���s��@���0J��
�����=19E���1���r�h0M;�C��k%��M!x��l�{��1i��Od��h��Q��i�t��ަ/�ӏ��?�R�L�f�VH �)Áhe�=�k�G�XP���_]c�B�BIk=�U��T��2Р&�j� �f���	n�jͿ�]{�Y@s_g�gSNF�i�v.�dkT��!X��꒛�oը�����11�G�}c����<`{I��N妆��F�snM�����5~_H9l� �w6BܜI��G�l*f�䛨�׍Y(�Je'A�h;�L+��e�ד�ܴFD�i�D��$�sj�T͛{�=SrY2Z%�%�\�����0�c��cUWq��?�]��&|B����!=7,��IJ!�B��}��0��������e!�[մ�;�S''�L��-2q�4b��k(�f�C|�n1�T�}<KHɡ�+]�H��dnJ�(;����#e�W�*Rn��k�iA:I��&��&|j��
{��j���YWc���X\]Q��T���y��s��>� ��7������Cz�*�8�I������sp��4>��/c�ԂB�X��~��`Ӈfv	g����o�7<SӋ���/�C�M�r�w�û��v\��+057�}�'p�w�&.jʹ��o�$���eϸ��߷b۶m��]��m��y� ��E�d���MRe
��]Zpj�n7Pɯ�E/�o�����]Ø^�@��G�'����8�(��<�jhZ��!J_200�Ɠ�m�VC>��C=�WFKem�Z�������(G��B�$z�	������d�jo�M{q������M���1��s����zE�
#E-" ���H16G��j4����@2ԧP�mCgcz<��o�~tϣh��ݛA���3�uS�~� ^<&�zN�Z�T\|���}൯��_=<���o4��>�[���;p���_���"���w�s�/>w72a+4�0:��a�6B2Lc�p c��܀9�c�?U����ӨV(��
!*���-��bxh�2��3?@�A��=�S
䍍p���7/����"P9D��p�g��
-Y�J� ����ƌ1�Z�l@\RV��ɫ��\��e8޹�Hؤ�@4��z+�ZӍq���M���Q�ǲ�b�̓��Y"�C4	��m��%|3���_.*N��f�E3���P,6���
�5�D����,!�q���:1��O�r�d�*��2|j��U��8r
0�łS<��`�B%�P
���C�MB�ᖛp�7�!89?����1�@�A�
)+��������^衟��U�+���;�km��si��0�o�w��%��MpD'q���Fz�**91p�g�soݸ�ڞ)ϓ���G������~kt����3ar�&>�hi��hx�,~?:%y�f3�˂X�I�(&�x�]�[{D�y��ɶ���~p��k���*y�(X�����!��g�='Q�::��B�bW����9|m�ł�C�u�h�����2��_�v�G�ژ*�B��ܴ�U����O�x��+e�I,:������y��C6��n�j4��lI�cS��Tq��!����ծ���9��[�B�~��K(�֥�j�_F�b#/�6�_�Q��\��a�lz]�=�5K�w�	��C� ��ߟ�Xd�z#�MUL�g���F=/�
�r��`p�����{��G�J�'���ߗ�rYr�@!�lD�sf2'�/���5lj�Dў�C^S#3���y�{k��FԪi�4�)���r�2l�.|O�sm�"l�,4l�����`Q�I�Lī���XT��i1�=�}��
8�#�/|�3�TA!��>��D�R�Z�`"�x���S�p�~��/�;Gp�=?���|�9�v����A����{�.��ӭ+���������έ�068�gg��i��q�����b�x��f�6�x�#��/כ&=��ɶ�%�qr�X3���¿��pfp�k�l��ISWBG$�oH��6�� �1<oXtrRV���c��ʫ���o|��&l&��<N�:���)�i�h0x��J9��عm���r���qhl�(C#{�����֏��Բ&����n��}m	{�ڊ��w��k.���
>��O�3_�2u�u�9c�W�<�:��E|�_��~x�&�����l�X�{�3�go�#�ڹ�����������P�uЪw$�U��I�M�T�8#��VE-���t���{�܉��I䊫@��|;����q|�8��5�y�h����appH{(����5T�E��`����t%P��P,��Ч{A�B8!��D�Y��C�j�z�:Y���H/�hr܇�3�k�\���"��@�����˟QmV�`W�j3�x���?��1�ret���OmEo|��F����w?����X��Ȇ�I��&��5Ά���7�Z	M^��j�կ���7��K��ߢ!`R�G���wN�/�����ܳ�e���(
�H���@�B�0�o�Lrƴ]-B��1��u����K�����S)�N�.��p��?{��𥟢܈�wlB���n�>"ТΚؕ`�_���_eH�G����.n��9���67���U��p9.B�t�n��F���]��F�<�;|a���������DBE1�c:������UW�=8z��Pc�c�C�W�J0��υ�Idl�j��x�L퇄T�Z��3��"R�҉��g�'1w�J��4��O�S���z���������W���T�h�78��'�M�i-�H 7��x�M�SCptrJ����CV(��B�C��x�펏�9
��c&:j�悑�Whڵ�{����1����a�d6�W��Z��v����Ԭ9�o��e�xv0�um�z]�P�
!�lQ�~��y�+{-V��pvBf:�z��^ʮ�&t�?\��]PD�e�	�HN�������S'B���2J��D�`gsO���$.�OAJ�מ�.�n��@d��� ��2�hs�����޽�i�P�`�jC����5�6��s��"Ͼ�M�4E�TN�M�6�'����(ɷ��b��"Ŏ��cff$� 1�	�י��deo8*S$�\G��sW�Ll.F].��k��>q�_ž�`�[��� �y�šw��|�t�=�ۃ�,��΀���Q����wUlcvp��akyX�&���P��)�I6$n��d�{�s�5s����&E��<�)L��v=w6��v�=���]�&1<m��D�,�5��u���ߢ��k�'f�e����/�f�(-���B�%6֜3���k�}Vw�5��� ���F��j��UыXs�?�й��E9�����}�4lL�h�(���i#Ѯ�S��MϺ/��*�EЪ5�|��v;��V�ަe4�>��b�^6is�Wq��8��fП����
���e���8]\YC�T��j&_3���#���N�.�4��%��E���H�MH�ʺIf�cP[4��Y��Q�X2�PH}��ղlO/{ڕx�o�Y�����,N�<���E"�"�fp+����AlU�����b�
n�u����C��/���&�6�Gf:Q��A�RG���Y�l����w�W]�ӓ3��G?�;���,u�.��3��y�[��Po61��G6_��BJs�h��� ≈�ώ�[�l-/�`qqUY!3��8q�R�]А����Y�FK�N�Å��X    IDAT��)\x��xӟ�	.}�EȕV����B=�l3���"f�f��]��ڂj^7NR؈r�fn���
����{咔N��,S�M*k�9 �)�F-�T/c�����x������7�8'=������5�v��)�����P�D�I�߯�c��M�?����3L��t��Ewl��1�$�!��7��1>��;Q�s���:6Ɣ�NZ���Yˎ��zi��B��/��}��×���##˛���ϿՄ���'>�����C6<28466b]��]~����XR	�%7,�]�'�C_�Z���۷��3�R0X8la����Ձ�:�;��(r� �#�ѕG��5:�Xa@�l�����fm��<D�a�DLC�x�P,�.�Rm�X�OvE�@D�Բ�QAb�'ȴBR����&�Q`U�
��X>�n��T����Һ�O�z�ʂ�,5.��P9g�����A/���%�isN/��	f<N������J�2uQ���'j	�OM`qr
��Y�U� �UC��$L{�ژ��Y�	��$5�Q��x(q�x�4B�"�3�5q�-/�57� �P'�gQ`:��.g��P;oZ��Fq�Įh�^u�D#�u��w����eC���Zw�q\h�ʎ��5^1m�Β�̽�k.HѰ�`�=[�&n���k(D�Y�Ys�>�I������5�ހ�Wn&�@�\^�ؽ�+������oI���H�Dj��@�u��U�(i 6^;��a�5��ă�E�����c����!�*�L=l��k�4�5��W�[A�A��6G�mW�{�'��O���E��K*F�V�v�y��>��������֐'uii����>����$ȡw?Ci��B�\�):���т��8)��4Q2@��*���,���OBZ�]������]�!G5���lE��q~�Ҙ�n��D�A4E��~�sS+�Ul"F�6�� �GZ���yϊ�{�5�^�Pj�j�L\8?p����`h�c�u���`sX�ЕXٹQ���kD��s�!��5ql"�;���	�i���o3 �k(��l�)�6*���sx�	�,k����p�V��I��D���ɣ�i�H^q�ϼ�97"�k'�_0��x ���7p�� 
�|y�>�l����MS��@��t�b�PXB��&Ͼ�U/���;�`]�>��~��89qچ��6r�sl61<�/��d,.
R�QG1_���6��������TWZ�2Ӯ�8p��xR�Q�hBAmN]�Ea��WMPt��/��M|�����2'q�:�{�rP�X�MM�����7��q�UWI5~�8�8�3����_�t��s3r�ZZZZ���À��.�������OM-�iaLM$���=�b`dx�)����1<~�$�u6�Y�p�0��T����?������1>~���K����#�-��c��~��;�/�w��"�� d�J�!>���;+���9��lE�ՆD��h��G,s���#�L��"�k�>�{��)��▗݌��4f�e7:���b~�˳X�-�P�"�=8D�O�=}���
�YX�C��G*���c�A��e�PO!�*uh�)��Vkב/Pbv�X�;�6L�7�4�q�4'h�9,�������Q(��'|&�{�ϡɃ�\����Q�E�/�x'��� 2�a�$��'�����;~���a4;q�~Bq�Cq�yt#=0Q�e0J��|t�[[@3;���W���?{ݫ?|�Xz�7m6��ߪ!8t�P������}�ɿ����C]\N?����)��Us@`�h�qs��q%�X:����i��|��/��z\xΙ���Y��I^ԁV�<qx����V(��B�w�pi���4VG�����\%���D�a����W�h���ڍHG����D��+�U���ud�z�+���=Nhˢ�e~�D�<7����&�0Z�-r�թlH8�0.7]�aԘ�hMJ�u"W+��� ׯS�C���uJ��W'��5Ug�ڕ�#I�)�W�6u�4�������g��'�^+jܨ���lY,ڤ��H�8��W�i��h�D���K�c?ο�\���Jc�TPCP+�D�b=���&pm�Hu�$�����ڨ�c���w�l#���:
oc��^H��?�^���@�7�V�xV��C�7�^C#�չ%yk�E��x��I։^t<��2y/�-��8{H�7�)�
_6V|����ikD�]�K���n6庡p�FU�!7�Q�!s&��i�H�4 j'�<t�gs����h���i<XXQH-�K�7���5���<]��(xMIXظ�3��#��o�缆`ݥ��2�����,G;No�Y��⏅��*%�	'b��[�[G�Yo��#�S"VܟxI�̺�3N��$JL�5��y�����6��haͲ5F�Tf��{ͨ�25�?k��{.�:�h�	=L���$��9��^�����,�-��U��֑7Y�A��P��B���Eٳ����]Zb�B��s����Ntnm��$�vS_�}pQ���}���#�{���7rqυ�<3��� �"�u�M���l�d�#���&�uq���$7�FǬ}7��o<���_S&�i���.�Lg���D����"�%�U���::��9���D�WKuD���(�_^�px�K�������S�Gp��8~��_bfv��V0�[�Hė7���\��dZ�6FFƴW�&��v�K��?ý���r�x� ���لќ^6B"��qN��%��+m4I�ؤČ7����I�H�4JEݟ��^���	����Us��'���&N��p�%�+E9jy�F�V��ر��{��mCW"��+�P�g�HB�}�c��C�����!<��(jM������hU[��r��3��\|�98t�(���o�{��)��i�0:փw����� �XP4�em3��go��)ڕ7A�\n�6��^�Ǧ�����_���p�ؓx��������N�fO`|������[R0Y+�B �ku����j�H5˭���Ė�D�!��p��癮W�V hďr��烩��zY�N]��pD@�Q����3��a4�S�iM+��NQ6����AE�t2�����!� J#�A"8����ķ��{೟���ϡ�g&]�l�K0��A�9,���8�a��h��@%����k^y�{��5���ӷt�n.��?�VA��������>��?R��hO:&��E�)��%�$mn��f"��!z���Q�ʋ7��^���A�������@�d�r�سX����r��'�����ca���?�p�K�H4��/*��f>�:*5�����핏w�VD�ZQ�?�Zi�ɲ�Z㘨�R�CruX���m�.yv�^�(!'� ��Q�M��%ٶ��h!�#��!Uǉd-$lÂ��qW��cꞐg9߰�k!���v�qZY�#�K�
H�:�VA�d�;�VBB��z]�J��RO4�XY^�\�X@imY�!&�qB��\3Q�j��B�I�`�/�4h��O��Ʉ(����������ٗ^�P:�|�E��������������F����^qh(��r�O���r�q%b�r ~-�U_�(�C�1w�Ch�{&��z�����_���ӏg�jE�F���'7�\�d���,�:�4kAZ�I��(@�f������ӛ�y� �x*e�H�:�(q�k�l:oiצ�w��-����%׻��.,L7�q���<;�U�g��y�F#���
yM�w��umx�{t#(j �wR��h<��օC{]�Ͽ�|?�"�~�2��B�H�$�t>�94�s� ��G�s��zݼ��5�E�n��������w�^M�����f��~%s�jk�\�,�����|x}ĹvT+6C\7֜l�ܛ>��:o��/�ݠg��߮�������L"<3 �V�MC�3W��#M����F�V�ю��������gD%�v@�{�k u�9�����^6�T/{��my՜�ꔖ��PL7=����D�8I���B��Y2�M������Ĭ�s/��	�f�j{�7�6���刖�����;��('�ԕ�Ѧx��C
e�Q��4vu��0q�&&O�Yͮ![���{��,g���+t�Ju�u��b���j���^����������#XY+ȍ+�[(�F��$�̲�âʹ:�DDSh�?�
�2p�sGc���OJ�e��fr�$Q~*Ӎ[o����$����"|�A���h�qz��� hçٝ�|�lv�2���s�Į�1��+��B6��P*�F�|0�L_=>���?��_>r��g����.�m��:����½x�{ށ�.>O>�;�?��^�L/�U/cx�K����f�a���@.�G_߀	l4Y��M�SdN'����������V�����H0SY �AZY�}��}�x>����o�ڪ�� ��{1�Zx�O=���,����2��
�^q
�AO/������U��,���۷��;�����v�/�6m�*z%�� :���>�P�}Saf����-�Mp�г��E�n�&j�*U��Y��$��u�Eӂ��v��Q_qZ�b�?̽g��gy&zWN�]�{r�(��HH�%��� X����&{���k�>���$�	�P�@%P������*�:羟��nq�?���K�LwW�����p�d;�5�1䓣H`�}�Ѫ����?��N�T?�U�(i���Ŏ-e����a�$y�ct�˨�W��o����o���7��'|�}�o?|ǣO�}�`494�n*�lf1r�U��Ӥ�4��`AUD�@�e��A*]�6�cm>�M�y\x�.��c#�.
ˋ"ʱz]'$�E��/ދ��|
M�!�F��E���ÈwS�$�ԆギS��^��[��֎�b�T��'۟�:�6�6�3����:�M��]?�TBB h�+��J'X�#���+�@�@E��T;Y�$[�)i�7Zm,���i-��`0T����"�t��^�dW��%�Y5gEJ��I$�[u�.i�m7����m�l�T,�U*`��a�� I��"	St�Pi��S��a���#�!bɭM��ĦMF�Z�f�@|��ظ}3�c\�J�Z�gQ4� &���f�q~��7���U��]���Y��3!P�8���^�f�A���x0�P@��!�\�����r���ѫ����(�
��ʁ��U�!�,pS\�1��LV�A
�!K���ԉR��i_�|��g�≉W��b &�$&����Zf�e�zUyv:z��A�Թ
~��.I��+�ϫ�
�B%�]�� ��������O�WH���`Y�d����ҿ"g��!�"�qO��l%�������%�=��I�k��m����d[$Yk{wY0�^��8A�}��k��x���U6l��IL\e(U��3e���g 跃���S):3H3�W�}.21��]��X"ʮ��>^�7�k8���N,)_I�W�0��Q>c	���X\Y�SH��hT�f�';����P��S�����9	\r�I����4��{Y��O�#^�W��h�9c�.��Ʉ�)����˻��C%�D{�.���!ut�FF�i�N��A
d_�#v[��422$%����<�KD=�6�P�Er�ܧ8\��D.�Z�%A���D��}({	}�:��s��>*����u�I%%���/��v���(�Lg�׾Di\ߓ��r���C�R�!7��V���j�)��҃�[R�4��r���Y\8H��|�.�LT�ok�c%������⋅l����ާ�����⢠R,���h�[u�����-04�~��6n؀5CcXZX|gddT��<��>�~�i|�O>��o�8�t��v&�%�yƉ��W,!xf�^\y�-���0sl�Z	������x��O�m���w��x`��յz�D̺[��'��]�v	�x���yz�x���vH&�VN�*�/21	߷G�Gg�<�_>�KL�N�ވK��Vt��~�iD�4�+c~�<�Yy�p�e\�dp8?,H�!r�)��ϊ��n|B��f�"��,�X����"��Q�hR���@+֑��`yV��9�|� �bJ(�������?��L<��ު�1�K�8��Y��s��3��"X�_���HG'Шf��c�p���a��004�V7���%i�F39Ź�S١�r�	:�Z�v(3K��ť?���}�����o\[���Uu��o�����;�C���Z���a5���� X�Yx3�A��x>mV����q���'�02�ӏۂ��6��u�X?�G�ۖK.7�j��r����(b}Y�v�^�p˃ȏn���0_�`viI�ch&�K�ə�/JlV��0�V�TZ�Ɛf��O�A�<�XJ-�B��G�s��C2��9��h��*`�NSMH�tti��lT0B���!%�d����m��F��"�d��)Qz<@-!�,v�u@ǩ�gɈI0�niU���]���@�C6``s)�K�}|a~Q��H����$�QbXIv,�I���j�*�i.��Z��X���12>�u[7axb-"�A���f�rV�ظ5:1G#X�VQU�A���Pywؓ�U��W��2����WND�@ǃD>'V56A�ȃ2'*Pg�E�V���b2s���0�F�P��ʡA����i�������P�Z��F�l����dV��bm뉶*�7nT��	��CG{A��_)NY#Y�*�8Y�8,� i,�:��$�d�m1X��/��%3���J����}�1y0f��t�LM=~��\=N�+J;�k��W:|L�ga�v���ú�Wt�6��$	�"�h��X�E��}+�ւ&�L[�$,-�'TB�0U�١��۪��1�.���m�$�����=�:�C�6��B`')jJ:��J*ufԂf%Z�Xݿa�eT�mUb��WKx�L�|=y�C�h �[�h���(;`-9F�9�9	������?�n�u��Q-'H�z��֌%Nt&.��P+��a��>�e��DN��xģ�P�:���dI��=V'`~�R�	][%�A�X��"H0���t��6��BǄ-�-�^'s� �S2d�� � $({I9"�H���A5�G�Um=x�HOJ�KD�����]r��Vj�Zn"�j!�*���<�dc��)~i/��22��C�*4HF�~ m3��t)"�%`	�'F|�wV%�V�I(X*K&�{cW<�������s|A����K�D��N���_�C��R���x:���k��g0;9���Y�c)����Le0�f��u������ظe=i�X.-#։btp��mB��t���G6�3]�DϾ�2~��Ø[*"Jiv�٥aW�N�ZB�Nė���8�����������]wޏ��ڵ
6o�g?�)\���cfn߿�Z�p�-HQ!G�TS��n��p����?��T�~��1����3��5Go�WG�l2�s1?��E~dhX�&F�'I*}l��t�p�wa��2��e��P�pt�0f�g��GC��|#�#�naqs���Q�r�I'a�ĸfC&C_��U��%TkE%�V�;�eg@�DW11|�8�L���w���j�� E&Jo-�&"C[7��4�b���E1�_���u(.&�����Ov��� ��!�@��E�!��G�:&�>�F����P/�VhV�Ԑ�T���C��o{ەgo^~U�@x�J�!��7o���{�+���!��4jى�&�hKK��6�X���-�}���Kyͮ`)�Hù^w�)x���-�J� (.�M�|v^�#㛰f�Z�yߋ��ǿ����Գ��B��}�`~��f���I����fU}2djQ���d�����:�Z�:��������]!N<%�)H��!#S��щ�R��F&�QFM�XF��ly����C��P��7�٫����aupK*�/
LǿW���B��*-�gVe����'�1���@�UCU�Mk]�E<8[M��寰0;��aif�n�&F��O�ը`z�(ff��ӬchxP��n�    IDATO�#k�
��Rc���L���mܤ���m) ϒ��t���O�1[(`��H�d���*�VUm�0����,,^P�<���� c�è]nD!P�D�p��e��'�	�*�l�20U0�.�%g�#�ip-o��O��c�W��+��^5ڱ�ڸ,y��W�4[IRԪH�Z�K�G�dD��`ǎ����)���˚g�jz����|�	-�
�;����eqς�:w#S} �z[.rm���p����J�y��6p��g����`s�sLF��<�����p�=�Qu�1�*ϫ�<�n~ߠ$��F�+}-!pO��f�@�Xz�����Q7��T�P<�B�a��X�H[��9f�E�VIw�C�#u荫mI��U��K%,����h(!�F%9NШ�	������)Bx�W�=�C��x)JH1غ-2����Y���` �	ǐ��8�˦�L	e��b�%@����N0�1Q�k��!���"ޠgI�4�G�u��D\�o�ާ��^X�@Ò��uq��(W���� r�w�������&�O�_t��.���D� gw��J!�aW�L�k�8��`������y���~/
�y�3��{X�+�8DIT
U�����/�[��H�����,��{~�'ۍ6�!�1�>� �sM�St�6ވ��B�G�x\VT��}&�ɠ^("� ,@ӿɡ)G��Ɍ�M F�vX���I�A���U��(��/��q��N�(�t�>�Q�����b�Qo�:H�h�/Y�!���ۮ5��pl���ڢ�w�zM	��M�Q�177�r��3y��z��%�V&ׇd6������Hf�]Q�T���|L���2��u�������N��߾s��b��N����7�?����.ž���+��o�]�G��s��-OO�1�_~9���/"�N�����?��GZQ$�݉��Y�X��d͋g�Ը�G:�B:�����e�ٺ�9'6l�#�&��N܆J����^��C�P��U	�46<�n�$�ݻӳ�8��m�&���s:C�\U2*�(Pm�Q�WPGu�yF��A��{�p�$�-.�ס��{� �K�J$�8�H�|�Yu
bt�xMӹ�R�Hv��@����_���?��ۃV#���J��u���������ܻ���A�e<˪�-f��O]v�y���~�{��)��'7<����}���>��?�Кlbhm��버Ig;(�x ��f��,M�}Œʸ�����78a�&\��ႳOF6��D�%b��b`���#7��?}w��Wh��8i�9��d��b�l}�Iժɥy��a���T:�5k�m�.M�ծkä	����6 �33�869�V?E�_2���_���Ϛ�@:��t��N�rQU!�7E�lp�j�``U,�0=5��%Sr���UMƑVO�A���#j�S$T�J�.��� 8��$v����#���� ��c�l�j�Ę��cX\�C�/���~\x޹Ȧ�4�������C�c�v���J����Q�X�N�0�R[��+���� ��T\���RE���zK���Sh�#��e@�s�7>�n���A��{vH�N'U~9���S��4΋��t��Ѫg
�X��J�Ϊi��靗T ������K\v���E�D���)禒����52$��X� ë��-)����A�o~R&מU��R�{q~���1`�r.��:�[.T��J�U�$�P	�ɇ���*�c�Ju:���1������*�P!�L%S��~t���\�=]u�"�� �&V����k���6s�2��x���=�����.U+���a�@��-�@�C�9	k��C�^�q}*!�q!���G�&���}���dӒX��g��cɹb�K���u�QV%��� �Sg��iaN��#r����T��^W$�����>ל_��j��\�xe܋.L0�}n����sHVXmΐ�DIPi�3IJ����� q$�������}�zw2��"�I&���x�K�?�ݶ�����{	��u�+(Q�@�a{�';��j�L?�.�T"�Ԩ��F�d�?�5B-��ٜ�[��,q"j�-b�C.rnP
~���W�yĽ�R�h�k���4�3^D`�V<�֙��a�)�*	/�ϣT�#�j�/ZE{�0N�6�����E����?��ؿ�"?;�J�d�!����XP�k���ɣzFJ�#�7�<�ѤCp��R�cFMь�����h���1>kq����_Y8c���м���ݯ�o���ޠ{o ��~O�wmo��^mO�f֦����S*���!%B�I2ܴ�#�,6lڨ���[Z\����gg���Qr2��[S�Z�8�c�0�t�h,Ma�v�K_��8�S���}���;p���`�Ф
7;O>���'p�_�CS���o�u7ߌ�i�H�(jRB4�����n|��G�`w�q/���������U�H�T?�ev�X�`Aa��K/!A��중��B�Y�Q$G2���my���s�߀����+�<�D6�BeY{τ�1�|ڰv�:��sxz�3R��:�8��y&֭���("�6*�"*墒�B��
?;A7�����h�e�A����kD�1��T�艔ؼa�M��@6�D�3�d��l"�Lz �� F��!���n�w��a<��!,OV��ax`\�ކ-[�;�{b�n��x�hw�B��5�k��v7�����Ld�?���Kް�_/8�D3�x�_��Cp�CO��?���x�
�Ǔ�<�}L�$1<YG	��,S�T�@�1g����t�lС6�t"�f��l<�Mk����5��01�-�cӆuF�f_����x��$��`z���%��EI�Ku,,,�&Hh��e�sX�~�>�����˪Z���41r}����fu �_*,[��JK����k�r� �M	A� 1��*�k��^o`~i�bY�!�̱"6?G3��ԼQ�&�>Ӝ(=�j���2��{ qqA����vpG���KD��s��k����@���tǎQ�D��SN9	�� ]���R>r� ^z�E�3)��X�����0�Ŀ�ZS��)/��\�R��H�Y5�h��M��C8��S12�/�?��}
�H;N:#�kT-�k4�t�\�+�a
������,��@�**?�u����*���r��Ai�o)9� =�!�͆���F�4�>%J
���ǟ��Mp�:#��ì�		��� �ڨ�a2�RvP<i�����K��Uh��]XR��=V$I��6�4's��]��MS��rn(����)�y~_���
��ڔU��ҧ���A��%�����	�m��)����$F�5x����\�`T5�*v�C��a�F%2B�	��+�eWL:�!Q��ρa4֦�tq�?���9�Q�D)�Tp�@�{r镠^���H>3=�|W��e.�#�C%��)	��1!=��߃'||*�1+��䌴I�a<��<%�LQ�9tr�X�@Ġ�k��� ɫ��g� ���p�L��$'�y�Ġ��y����]?���]Ak�q�����ο^L�������;wY���:.4{�9�`���H�v�+����y7�� <U�[����Y
v�	�Q'@�� ��1�q� S�=v���IRn.����*�i��0���5����GN^�P5b��/7m�� �	qal_�{3 �4*M��)�P��?��;q���C�p߬�2)�!�Y���ʥ�� ���9΄�I*�m��=�m��:B��������/�����ǑLF3�]/JrJZY�7� �����G:�L�U���H�H�n����H����%�j[��fEE�NiI^<���$���}��Q����v;���A]��L��E�	r��I��v%+�0��%����Y<�"��i�}����~'���<���яq�]���\Rc������i�����c�q�Oo��tf���0������z���.�����0<2�;������'� N)��a�j��hxǮqWL%@��������j����m�������sN���q)N:}&�b��Q�/cny��E�9G��hM����
3�&g�077#��uc�رy+N9�De��*WQ�_��d�X�����͝x���ϭ@%��(V	s�-���%�ɣ2	JP%�A*�Vw ��!�"�C2я�����O���'17Y�Q�F�~�V�;x'�~*>����8���F��އ��\�lc�d2�1����������ч�i��g�z����޾�?2t�O���o����ȯ���G�鲚�E\ʎ-�����%I"Au�	��ϙ����L	"v�Y)�۬�U�a ��5i��S�hxd��a�y�͎�A�:�nLM/c~���h��9�<x�4�����e>2ڏD������r2�x�Ǵ�1�E��Ĥ�?�ܧ$�M����翉͖d`�Z�N����l�3�-������/?���1�8H����?��8�^ͤ�W|�j�np|_�Kx��X_�b��q�����
��r9mf�cb�HF09yT-��۷b��b��;�#(��739���퓓#[��_f�� �I���`� '~����>��s&6�T��2\x�8rl7��s�/��u�	ظy;��(�(#k$h?p���o5\��h�-�u8�W#��CWs
I�%R�d�I�$V�Z��(I�ZwafG����LU�N�C#j���1WQ�'(��{�U���\�ܦ�է�ɯ[��h+��*=~���åX���d�B����N��\�ۧ�A���#����}�!*:n�������a��X�̯���{&$��$x���מ�'J5������<�}���ח��z���<a�h	�(\aŏj,$3��*�̩��ĞR��\
�F�� aW��J�+������U�eZ`�O��+I^u=�����۵ԙ	��ꍦy�����`��,�x,<���v7���4WԜ|\8����΁�O�=I�3 �?7 ϒz�	qp�� ���o�T���1.*E[K+u)�L{��ɮƤ��cV0����4,��ɞ_�Uۙ���!�����e�d2���F��U�1��r���v"'+�%n^&[ܟm^Ɠ��1һ%ά��9�sV�3����B�FC/;�b��Jؽ�z"����Ɖ2�u{�(2)�|�E�̟bA.���"
�%J�O_^�G�R%�IKZ���I���T�Z�#Y�jꀼF��%�"�6�,�q��_�S���};�ڹT�*��#��� ��L`,���3�+�f�(Tbm�I2��{�7���p��7�W]�F��X�����Dt��	M�����3�����w�EV�e��T\��V)p�|~��5����N�U�q[������Т1UgBp\)�0VI�����zC	�c��1!z�oj��3���״\D���R��A�F	�{6>���c��x�ɽ��w���w�+NB�T��m��/���<�����݄o}�����׃F&:�zTK��?�ןƚ�	�����������O��)ˠK�B�T0��5	��r���ю��,[$�f�V	�0�i��B���]��P�/���}x��X(̫�G(��Р���MU|!����G��bzr�REJM'n;g�x����&�d*ړk����j�����[@8;���L8�:#�'�����^��],���/u��u$b	��Y8N!˂�ԅ�*�6<��r�?K#�Nڶg�:�n?��ϱ��W��&6m�5�߆k��S��H'�2�l
ȍ���_�~�غ}7]sC!�h~���^������y����������w�c�Hv�:�d$9�Ĕ��"m���!0�w4��&�lXD1�sE4d8A�gL�l�XE�/�A�@_�p��@���H��0��(��8vtŒ�|xܔ�V�'	�mg���HM��z�V]r\������f�dΖI*��-���f�΍X���!��̉ō[Akh���O�*Y����4e���(f$VظQ21��� 	c�fR7�h�΢o��4=@�B^� A�a�M�AFh�b���km�Ŗ���ЮK�I�*!��I�p��S�X��5�v[8U,B�n�!�`��R�(0�N��d�7���p湯�e��Nt�	�s߃x���&�^�V+�J�/�a`���W�}sZ�y"�A�W?�a�P�{�j�.J��*Wܬ���7nrzr0�|?�dp�;��+!����|���\��J��p�e���7[�H�1�ܞ4���A_%@L�i��#UQ����5g}c�k�q*P�p��%e� �piEwY�8���0Ms�_�L#�ǫ���������_��ą'�J��3`�ݡ�}dW��.�^�[�QB!�0,vR8��jo��2�VמI�3�Ù		֞Lrl��?vlR��d���!��l�m�r�)y"&�@�:?r9�v���)M�!�������1'4��F�5ּ>�T�lhPl�`��� 1&�GvA�~�W�y��{�|���w�<�Q���0���m�B�8N�x]�+�8����тe8I�v�al�`�'3��upb��R6?3���)�rY�'(J�h����r��{���CI��RQ�[�A[�R��s�X�kTp ��<�k����ҫE�>��������g���O���C�����%͗`f�y��¤�2ˁh�N��c�J���)��+&I��u�T(쌼->+%�u�v�������yv�0�Yj�Vx��	VM��a#���VD�x�o^����Mؼق7�g%�����K~tg2i�A0N�o��Z�<2�%���4d[����#|����j�/J"�D����c�]ж@<;��3ɟ�?��N�bQ�P�@�C�Ԛ�%��T�����A���o������01�r�hgd:a��VS
D��kRҒ�⢠T��x�*as�]&�MK �|D^C���R��j~,d�����]�C�̳����]�o�M+�ر_�����o>W����ǵ�݄��y�sٴ���� �o��-��?�}��������^: ���b�n�Er;ˊ�S�EKY03v-��6tny�.�]
@���O=��}
N9���4�_~��xH*A��1f����ؚe��xS��Rx:z����D$�s�8o8��B���V˅�+˨6*h�<5N5;S��z�>�n��E�|rN�������sR0�ZS�m}}����JGM㹽�Ш�1}xO�~�П�;.��{����������&�'?��p��;���ŕWݨ��Q'o����}2��#��3�:�<����C�����>�k�n�j��W��� C_��������i�T�-��(��8&/i����To&��fB`�Y�X�\�*�l���E��p�&����v�~��O=��s��h���઩��9h�j�A��_97XV�٪��X�M��������h3�U�2 �Y����j��|�B9'Y8��O�z|O��]O���saUCFt`5�/�o�*
0Ƥ�`�V39%�n'v������m�M�ݑ� W¾)����X�P��3����Mt�4b�H�I�>��I�$�% ܭ(�ը6ЮU�70`�`�����dK�b���bs h�	�#僁�a����q�v,�*825�C��b�XA�;߃e�y������3�j������������7�{�/��x%ӡI��
n"V�Le3�J�[�C��fh<���iⲊ�?����&�=���4��4��-���🈰���(�-9a ����U���lϭTd&��P{U�R�1��F��B|xP��k1��*�:	0�Fȁo� �!:�&Y���7�Z�*��߮jdFLA�c���2�ι�� e�����_O�n�>+ry��3@��y��01m�B���k���
 �-�2h��3���o4�����
�j�N�<�u8	�>#�u�u�jl��k~��~����(���!��vx?A�\E#$3|��\ŏU	��`�fXxK��|U�    IDATi��;�����ý6�U��y����K��!�G�Z������{I����I�M�@vh&?W\��u�(���'����CG0��`]���ض˳����9f^PR��7�3��4ߛk�������}�Iځ��}H/q�����b]KB��z��2�tp~���xB+8�s�.W���������g�g��#�dI{]��d���{W�C݌R����|?*,�z�:�����bX��T����G0�Ob�ݷb��Gp����༳�m�����7E/�\��bS#�C�3�ߏ�����TT���Ȃ9}4"$y�	΋/Ə����q�xe���9�M�~e3�_^�����r�U�!ZJ��Q��\*z����R��"�}��E�P�j	�Oڎ�~���߾�v�2�!�Y��p��P^L�!�	�B�O�ga�Xo�<�V�4�N���{��uH] "&&�n�/C�	<��!|�?�Oo���Z'��_���E��"��B/��
�J\P����8���ڵkp��;�LM�����(�����֝�w���ǰ{�c�<6�N'"*�6I��]�궗��:���\ ��X7��l�o8��s2f������Qk��	` ����/}��nۄ���J�KK��<���9)=mZ�g�<��t
6�]��d˅9�t��7�#.���9��{��5`�S��ڞ��T�礮����R�*�Hln��#��p`�AL�G>;��t	�?��/`��6��?��^�>�t�|�~E�?�����N�<���j�{�0���Ѿ�oś.z����*<������o�ş��]���~�����o��o^��yi�����Z4�1]q������ԄP��k������8�Gn�j�;4GAv0O	e���eX�¶��Kr$_'�Uhy6���ҟ a�]u�jO�"d���
-p�W��00�,�����xhK�B�V�d����j����9��[��7����W4�l�\~������werS���>V�m�����c��+bT��É�b���F����*&T��R>���ˊ�g�>d��ޕ�����Ԟ�S���hbt�l�q<6mފd6���yLN�"'�º?|ͯW��3�̃�-g�Y0�c�)P'�(�{tI����M�\�md< 5ށၙP�T:�"a�V�E~+��ys瞈��5�<`�qu��ϻ��IbY�j m�:c9b��$g�����k�[R`��π+�b�	=+,�:gP����fn�
�R$2 ��*�N��IԂ+o�SJ��LS�a2d�&��a F��|�?O^�'�
&�ɠ�l�*��=z�Wi�z�O���:P ���q�`0"}�2�G�;,ύ�<q��Qߞ����`��a|�*լ`�=�o߮g�
�%������p�P	�Ǉ��H�k=�5�x���0G��4�K	]���0�k�jp:&��������W5?H�x�WO-�3.��e�~vp��G1��S�ˀ��Ov&�E�t5�t�#�ϋ��v8a��4B:����ʺ/�iQl�k�>#��`Pίo�.%=!�{>����EAcx+�=j,�q�� x�O}v��}��9V\J@{�S<���'D4��H*_SRG!$Y�N�Ln��&^7��`b��4���g� ��[�1� �8�f\�l?<ѳ�ƀ>�ʩI��*O
q�Ӣ5�@��s���Iӭ�1ڗ�i'n�h�����^�UA~bTE#�G�f���R�A�֙��1i;�3�ћ������̼������Ǆ�	Α�<�̋8xtF>��U�ܒ��u�����
n�8�.y(�	B,Az�kO՚��	=��o�9����#���<��{�$��Zc�x�e�ୗ\����)�Cc��,]O4b�UQ����fj�Ȥ�:����^��f2�^�q�F��Kt)�A�A?����7;��z7��S����v�,���7��_�K\r��9`]��b��l�6��$o96��\,(8��]�54:��{����<��{��2���+!�Pb���L+>ȏDP�2ڕE���X�e-�ص��s
r�iT��;�"
�E$9��.�2ff'�~�Z�8����a�R���ff�035�v���Tg��'w<6ML��9�:�ޛ48��Q��&D��k��q��YVrًٌ���&ʸKA?�@�RǞ^ƞ�/azz�J�Xù��2��!��	��7ކ?��a癧≗��?��?bl�Z|�C��M��{Ʒ��}<��~�clٶ�x�;�Ƌ�]��p�MWa����>��~�S�~�ͯ6�׿���﮽�o��M�8\���@;݇H�n���a0�Z�!!`&�w�}�T 
��V�cIj2�@4�̈́A�O���i�!�`B�(rV i�&�x����QI���FuZu���*��V��66�TVAw�L�����iMX�*����7b|��j�L_\	G�d��^a�d�P��TL�x��˃���w�(��a��y]F.cc7���*��*=X�c�yR6��L"iUp:FJ�;�<��}T!�P�8u�41�
����B�9��I��Z�"�����e��8���������y��{��0�z���kC��/#���P�@N! 4�aB�`����-n�RU�tQ+T0�G��9��?�/g���UVTH�}�~����!yqZ�kg@���d �����DB���A��B��CH��\o{�ǲ�'<x*$��ҝN�X����&G	]�x�m��JeE:2��ł
^<�	�Q�֎���ÒA^��-vt�%^?��C�&[��ڹ>y���u��y|�~{������y��^Q-�_��Y>ļS �\܂GB8���~rέ[�^AmqyY��j#����tH�@��㶙�k���@1�&��P�lvo<`�V�PE��#�d��л���^N��z����x�����@���U�=XQ�r�m)��Q�T���ڊ�q3��$��I��Y��:��ך5Q����@�m�&b��8ӿ����1�Lk��q�y��R7>9?���Q73r�-&z�PSj3�KH���Up�DL���d)��>�|=�ǋZ�ˋ�4I��҉g�߯���qN����4�$��*8�!9�"_�{���?v�ǆw=}W��N���}?K�=��w0����"ŤnTFW�b[&F�מ�H��[��
�/=��?� �g��~��E8��5x���:�|�����q�ӳ8v�(ftJ��i�.ǖIEJŤZ�ҵ���*����r�oøIgT��{6��[�����ƙ{��͛%�̿�y�]z5v�yV2Qer���:
q��i��qg���#y�"-pkO����?�j,�\n�W�n{�nT�:yQ�s^&��*���^g�0Rö�	<��~<��e������I'm���)\z��������j -($��F&�,ͮ�91h���	,;��"��~\s�u���s��,	�N#K	�KIXk�P�:*Ouq�2�)�Y;��'n����!?҇�3�P(/ �d;�F����#r�����w`d|Lh���2�gg��g�M�����l�׭�x���X�f�dM�k�I3!���<-%��5���n����?�j�ff�H���9<��s86I�^���8�<��,N.�5g���]�~��͗`~y��z-n���~����?��lކ_��>��7���ۏx"�|�ø�7���Ǳg�4n�����޻��t|����_����'I�������8Zj�_��t?"� �0�������7���̫cx^����#8c��S��5_��b��z-��5�֒e��-�B
_�*�R�-HIF�lYB�Ā�Zɂ0�>;X��[�ePS{1���ۤ�-�6�E��;�I������A��`�[�"�Jf�&�%<��c���lF
'��zx ��o�2�UZ?�V��������F)I�Q+��fS��L���DĂ{�Vu��2����t-�� �ɓK�*��}t���Nj;��2n�U��5�Q,.�����8��T�؄!���1a;+���{ld����pK
����o�nV|:j��I�xB%�!����K�$వ�� W�z���-�-OΣ5#���l������a�R�����3������a0���2����dPE��$w�W(��B����<���(�h�����സ\T57�?�����p�feM�c�a<����	�C�����t�*�w�L������@�{����Uqޏ'l� qȑ��df)9G��H/��a���n��t$#��j���ǒs^z�����4��y֒rw�V����)Qv�a[Y���^Ʉ��*&Gf�F9P;��m۪�"���Y���Zf�C�&j�3@OƤG�&1�	��������&~�
���l��7!۷nS�{>v옞9�����cG�0�g˪��,y�^̹ R���7Y{��^/�{$-o�՝3��imH9%����'XS3(�2�M����a�Ν�2>��ӽq�VCz �kg��ƔX�&s��hm8�z�%B|>����(��NH4a2��y��>ǅc�E%n����sA
<�+� ��_C����1�+٢�ձؑI�iu0�g����g�k��[+.�
Nپo�[�0;�����Bcv
q�����4�����C
B��0��|,I�!!N<Jߟ�Y�+D���Xs��Dȁ"�N��ύ&ɹK)9��B��8aM�B7@WA�B�I�!j{~��f�l[�n���K(���May9�q�Z�F�Z^qNhT��&�IS��p$[��MI-����^��w��<+��l��ܓU�{��U�Y
�Y�{t�-�
�-K���B�֭݌Z���r�D&�u,��Ν[��8.}�&fg�P*�E�N�鳑�>F�$"%�G�џKh�]*07��X4����ಙ���=��sE�ݻ�S���;�Ʊ�G��!����%�)�b���1V�)�̵���1�r��Z3@�2*�"*�"�F���%���09uXR�#�ؼ}3F֌"���7�����4�utjd�ql[��m݂��<���2��zC��PT�N����Q�sO���ۏg��VS,C�C�Caf�����/ř;�ć>�����H�������>��� .~���|[�l��n���������p��.�G��8��M(7��~��r�ya/����w������7ڦ��^U��o���Ӿ}�m�8Zj���(�Cch������(op׊F����[F��D,x]	C���GV��T5<�4k1w06dy�3���@~�s���W���zτ�P��Th�"gW.��`�
\�X�%�
!�D����W2݉ӯë���LQ���5�|�i��A��c5Ք�k��?1�j��I�WV�o0���F8��*�g��<�Hr,���YоRZ�a>2A�gĄ�*y����ղqrC,1r�됸�-�p��"F�ҁ���L�I��[�2�{��+�.�P�聲�8�=FM>L�N�|2Ą���TmiW�RE�?��A�}b#9B�N]!:i'[��9o��;��pg2�1�+���r��ʄ�EU� ���V~�He��Ԫ���4�d �˩OWRVP�Ҧ����z$���:5|~�|��k��Y`044�f�Dɞ�%d$5�!'�8�aʪ��( �$���d9�#�=�P���dr��+��|1ErW���!�Á4V����Wt9�ه���_���ϖ�Ʉ��4���(�c"J�\	���p�YE�Z"��ő��ίf��Bq��z%F��(�
�~V�W�(����ú��@�h��2XY�2���V�`k�Ǘ�(}r�X0���'$�2����#���f��׼#F9$P��K�cغy�?4����%�#��$�y������M���θ9�XնĨ)i?�CV�Y�z)
q�\�.���-U���J���C�={��Q��I*�֬�nk���#��k`hP��~� �z�|�<��k�Q9Δt��s?�:cLhB�c�� O���"1�&`���HH"c�$�;Ns�/uH$��6:Lt�g`�U���Y����� eF3�<��l�39�b$���^���:��?���t`?y�=�#ƹFY\���:��&�'�tӖ\*YUp�U���֩�t�6dU~�KM�������E9�-�T�C�d|�<��ha�o[�ƹ`��ǎ�)av�7����3������ӺW��{�+d	W��@�}P:,.��E�޳X9X����1�9�BW[W݋t��^��/U!�{��3!t6�e׎2���tSga�<��w���|�S���s15uO=��x�t#	���\-P,��o|-�v�E�"�<��7j�r}C(Uj8c�����]R���Z��+��cS�޿� ��t��0A$�>.���*���<b��iq���F�e�f�y�N��bvq
����3��M �R/��8;��ĺ	�ݸcc���F�'(-�(UP�PD�K��I�1��c��uR%"l�
�ƣp����[й���q�r.LNOi��+�F���їD������?��v?�3v����x�oD���=�~p�5ؽ�	틯����O�)֯Ǎ�_�o�:_��O>��.x��7�<�,�|��~�	L-̡/}�/�x�'?����Io��ʿ�����߹��������E�m#�?H �f�~=�L-n�Q�:4�an�7m�ʔ99,�P��R��2z����+u�R���"#,ː(@n��`�7X�-ᢖ�%M�Ӎ􂙫�Oą�	2�v������C(��h�~�t6L��_�M�C�_L:)�!��x=[��`��N���W�=�v���d`ɱc%�+����a��$Tὅ,7���`=tu��� ��"E�@�6o�S�#A�2��`�=�d���Z�+�%8MH�䨩�G�00U�B˛�A��$�������Omp����޻W�<0ӝ����B�WǜB�`zBƃ��W��mY�ƋgŐ8S�B�u&�b��>Ǆ�V�x<��0���Ȥ��'�7�I"�6�R���&��C��aϪ�А�:r�jys��Zx�J�C�*���&� �``��C/�K��H��wa����#�����ս�ˣ�񼲓d8c��*a�p����[�:ܜԥ�B]���s8ׅ�!�f��׆w8��KX���{L�>�c�b�%Z[t 'V5$e���9jC�^�r��z�>���wW:���S��p0��U���'��9l��9���x%�:ԍ�b�7R�����޺Uά����~x�Z��I݇�uV4����w~p>;>C��S���J�/�l������2]325�������C�|%�a�c�%u�R�'kM+ y�ǯM�s�6F���N�� erأ��|O&�jE�CCBy��ٽ4x�U�C��w��ã�DI�d(�0x旺b���s�[��U��eA��\�׭Q �s\�@&��gıd���I� �>�D�(�	��u�*՞�?odd#�>lߴ�Nzq��w�w�C�:*��rD�nz�x��{�R,#lne��D�S���0��ƹ�<&���a�|�&�M(J���f��.�T���5ó������A^��T
��:;O;UPJ&����GaiiE�4jғbd��g� A��_A�+D�q8���X t�yM�Xx���ÅK,~�X���7	��BR��a��~,�&��S](J�_�h���y�F|�o��w*^~y~p�����S��_��!j��J��V��?������%���?n��O�ҾC(U;��_�q;����_�m[�┓OĶ-:Jx�Q
��o�5�^��/��1�H��MU�X��e�=���C�;wM���y��ݰ�}:��Hf��g9-�E4[5T�%A��0�q=�mX�5��KR:='j�%T���بI�~p o�Q!�X�����B�Ji�l�V��X*�8L�1dq�d?r�aD:)L�Ğ��bar�7��w��y������g��O�w�s?"�<�sv��/|�Ӓ������_܍��?o���Q=��˸e���    IDAT�gw��}���l`��@��������O����`��?^UB�g���S�����Mף�cp,�B�{-d��!���ΘJ��>��Z�$Ӧ��Y4��U_�Q�W$ض� ���η�2��7�Ʉ���	�\|ʕA�^���qm�.�hv��3�J�yJe(BHE�-�7,�*�<�	�D�W<�RO�-ͭ,�`[�]�d+y
_~����}����NXUiS&%��j�OAK�9%�`i���4Ң�M;n~�;��@�)#����CA�_�ê��vYu�S*K����~�<��(���e2ƍ�;6��w��;Yyu� 8AH<D\	�]��?�d�V�O��Ǫ9��rf�;
|nL 8^�m�T�'�3`1<n�{v�\��&V2�f��TV�?VA��4F��E�+J�>6�*�x��)�n�dp���-8�Ӊ�#1��!I.����"�,�)�$�$n�1���BC��Xg�s7p	�K�*l�V鷷:ґ_����ܞ^x�{��L�e�a������E����������P�1�,��w���0A��\�<$MҨ���hx4������a��&�UYÞ�]8�C�]�N�(9�?�Jhpo��}��;�TVY�P#(�9(6܇>�:,�1��f�%��	#ׄ�ޥ����.��;���ͫV����=�1�
\��{L8^�㰺5�����ӡڈ���H�@k�$iI���~O�ezct&\��<�m۶mul۶m�NǶ�tlw�a��}�of�ܙ{~W�U�N�]�jX��?l\]�BTƶe��M'����KGF���#��Z�}
*� f�Ks����o�Ms�?�b��%���iΒw\���@�w�)S�����'V9�-�V2�h{\�B5}�����&a�.���Wd?�u�Z��y�/w��n�{(��X��X�(�g�n%	F?��#�H��������GQ[]�[�js�C��� ,�%By��3šp�Y�Q�|���B����qN�^ɳr�<X�����W������2�7i�����`LR�1u�y,����x����s�#<��������P�N�aXA0�Rf�����E�yjy��ۨ��Oz,��=ǣ��.j�Ұ��墵�r5�H���z�b�;D�޶�c�Gy�Q:��	��$������y�4U���q�z���,��d�.��b��\�����A�t�>ܲ'f���sө�8��iR�a,����:Y^��Gw���^�������M��j���k�mWz���޽�<؉�`�+K?� 0��u˃���w9.�ya�`/=Z����|<���F���.�b9�a��U��o��-ɩ�63Z��ۢ���
8�:1]Z*�ӡ��Yf^CH���7�#W�?���Q��a��a;����|0x���������i��U�Hپ�m9�e)~S��:���)S��pI%e��	ul�V�qs���sן3W�Tr���#��,�]�]������W�����
%���>M���^Qлe�W������)����W�xv��[���/(��ɇ%N\�ւ};��MGBS0A�)�a<�؂z��ʳΌ���E^�"�P�n���t�!TS��DV�|H���Ï�ͺ̓�h����]�yX��?afj/�JM2�$v95Ra��UG���d�F��v�ۆP�F����"����e��t�73���-|VL�gS�[��-��Gk>��N��$���W1Ibv��.������r�Q��>4D5���|Q��j�h:\b� ?ݼj���i�J�� ~0���3aB��n5�j'<O~8Pm;Y��ĥ��yO=�eP�_���80c"��XQs�]7����f�tEE*�����=��E,%����\,3 �9�K�q���#��&�����i�ˣ�)�D�_$㋵�����3e�#�Ƞu�@���S&���#4��.�n3�X���X�v�(�Ii��k\�MZ��'c�*���[TV�6>��ԇ��N���P[AA�
�~�\��WV��|yDf�dZ���Qi�aE..� ������߇i�}̿������X���y���-�6��a���Ggq�.�~U"�Ës[������X�������i|���_�4T��O�r	gPB���i;���"g�Y�ff�¶i����ؤ��w��{q����r��	u��g`��""F����^s��Jz�X�`�i�+Q'!$�x#�I�M��*,�nH���UYn��0��V߮�wY,/��^�L �!�mvKª]lJ�Y�m��E$�,ٯ[�`G�Ds�L��������"�_�J �ûA�nL?�X����P]~������b�G����L����K��AU��f��D�HV(�a�ǹ�]{�a.d�Y�"+�O��;�<3�,u���Z.�rX�ٟ�m$3u� �]K�A�{}���f�Z:tsV'��Ƅh/Ѻ:�T�E�Vꇗ�-s������վ�����*c�^P�|�O?��Z8�3Y	�����݀f\��!g[�l���5����͋���O��b鼱�\(���v���r�W�X��I/w���q�������]�ȣ�Q��f�&���|Bo�{��Myb�R����������`?�2w%Z+��X��&=�l��5}⸝.��ْ�4�Ua�V�*�=/��wQ���q�OG�:���&[Y��:�*�{%�'+ŉ�����p�;�Ĕ-N7Z,'��}h��M±ɮ��.���]����x~��s"D�}ٱ.B!~��D� L���0�jX��}�{�jGK�D���E ܎<���5��=�� ��5�u�ⴚuR�+�?h�A�:w���9
�|Kw��P�W�_ê0d!��#�mӝ�X{�� ������u�m�_,ˁ�If��Pm��=��ӻ��G�����i�z�ƽ�n��Ճ�`�QG��Ͻ3%������Ԍ+�UO�'ߦ�2z��C�u�9�"'$�ՕB�f�$J�"�6-�uƝuѪ�4�k��4�ž׆�b�]���~%I�6ߚ=g�+ʔ9�eA��:�v�J3�i��}k?���*4��hL%ʞ����g&����ѓ��|qҒ#�M;.��ҳb'΃w��RSFҤђYq̤�>�L��f�ҽeɪ�8I�b�-gƝ�Dщm��CyA�e
/�B��f򭝡5j� ɞ�� 7J��R�g�q'�L��~�Ъ}+I���,��]���,zR�y#�!'a�4�3�U�~tO8F���ogc��/�<;�	��f���Z">�b���<��Rd�� MYy�a�8~�9,�1J4*k����d27��F�a���ds�+眚L��C�b� X,����f&T�l��2��9;�_&���[Oy�thPP)䛾��>�뜚�c}	��V6a�賂"S��V���lث�"�af�h1BE�Ɗg�{���9�x$.:��/A����*�����|[��zϒ�^D:N�(r;*��<F,��r<!���Ţ�@(w�e�5U��=L��P��.���}r�yƧ�����8E�<�g{�X0�Y��V�=��6����2G�"ؘchà	�R��ȩ!V����gn}|�{�?a��$���'K���hL��n0�1��K���}�?�ݪ����%�$�bw9�F~���)d(BFA�CzT�o@��;�!�=9��7L���:'�2��`��'�>�fo;<BV�b��� ͜�g|E|2dY��GA��B��P.��ui�����e��t��EuZ���Q{Y��E8���e����D�����1,3P�V	���b��q+��;�eA{�����^�bH�!�y1�;�@����3=C�K�}Ō��Cd%�'xQ��k����d_w=*�i���QMHH���Jb=�x�dB�2����̑��@*�v=RgX<PC�H��S�wk2a�x�@��YO�x�B�"�-�Մ���M�i6}��r�ïU��Y0}0S�BC�?�*Z,0�>�˝�N&�b�.v���]EB{���'�="��{�sh�s��7�,��x�ґ2��A��r�Ә�A����6��8Y���X�x�w���Ϛ�.So���#�vc�	�嶃|�G�g�~	UG{|���5��?^VyoK.����Z�%9�L���{�UY��{#J���|?__�!��)��)	_��^��4�����'C�Z��X�Z���nH.���I5��μ!�:�Ha���T۹���As��j�ӡ��-��P�U�
�qB�C�~�k�禐.��ʃK�j���l���\����~"��!FI��J;�����go��t׽+o?���44��Y���|&��9�]0����?2�����aV�:�y�>p��e5�#ƣ6�Uh6N�?���s�Ѿ��/��p9���Y��k4b������F�o���"��"�%I�RʸH+���p�@W�v�eRlYM���S�<O~������uԜ���$?R��ּ�+���"{����'�/��(O�����2m���G�E�8�����[�ƥz�Ʒb��
�������(r!�*t�
tI���4��/�q�:�R-�1�2�<Jv�٫Z5{�]7k]�0�صg�0/-��m��ZucƗ�ބ��	��tf�yǖ=:�/
�vRc�q��t�� �X�㟹��uڦI��j�2��Vz�l(���X��ڱ�L�W�)/]�)Ǚ�n�=�u�YV�ī]<�V/����,X������r�Č�<z���IO>�n~\�n;�S�i���q��
�D�jԬ�Ք�^�aӉ�쮞�˰;r�F�i�ސ�M:M�ű�Z��8����6��-*�v�I�);�?z�oZ���a㉕0�p��I˩|�?�ѭ7]�]̺F\�휫��4ؒfa�b#6�OB b���BI��BCah��2������
I�QJM���趠	�k&ӗ��wj������i_�ZW�bLb�@���w�<v�������wE�#�0��ln!��i�A��u�$��c�#�ܘ��G.�B�[S��m&������5��hlW�"���r{S$G ҥp'q�W5�Ԏr�����G��b�v�o[�f�k='Ilid���W�	�c.��<���n�7��i g��]h�{�&�7�tQ�:�`�%ލ<F iV����q�T�K�6;�S�n�h�+��h�F<�eT�\�{�M����YR��(o,n$$��m�L��8^���	��]1�Yx���S<[������?����{�}�Zh$�c��G����c�GȎ�UBt�c�2��q[w���t6��zlF��S(L�*B%|�ez�3�#�ӹ!���1�oBֹ��l� q�������j�et�F�I}zl����a8J�d��[va�wau����}H��V�̆<!`�8������y �X��Yq��0m`�'���Fh�'8����/>g]�y���U��cTt��64�M�W �or��\�z#5��O�bN
�q-z'��S��"�A��b��>�c;��`X[������0ץ.]��z�ȥt�(���Ĵ�+�[oc���$�>$���c�pV'6����pk�~���T��	aV#�ü�W��i@5aG���_C,� �t,%
�Fi5����o���(������0����N������#���ta���	����[��c>	XFc{��Fܫ�)2'�{�9,��y}hV'����G�3��N�Ukp�����!p㡽6��钳���\�򾕭/���여�M{����{0�X |��c`�|�<۬"ɝ�_{C�����V�^z����?/K�懨�Rw(_>��!"���o �ˊ;|'�Ͽ�~O��������.��KV��rCNB���>�1A��P�ȴ�g&6mMeâ�!��<L�����b���8H���ǂY��EU.t���K���+�ct��A�/��F��S�]�,�4����z��6g;$��`ɽI����/ue��=�q���C��V����9�Wȿ��8]p( ����z6����=��}�v���0Y-(G����X�/T~�u�����s���T�%?����<
�t����~߿o�����<{Tص�P$|:�yB����Z;),1-���X;t������ qJ&Y1�YuW��ڤt�2,]]B۬��uMG�!��]��e�-��j^C!���Wt�o�3ow�R���ʺ��ͤ?���Q�[�
;��`��]Xթ-s�b>��f�)��Qv�'���ӝ�lt��K��լ�Q?�����Qh���}���i�ֹ�3s�꫟9f&�աks����ͤ(��g�ʼ�TE�y��jh��N28ȆF��?P����eW�"��&_�����:R!��{���G�[��P����ﶍ�,C�6��?�>tN���!9ą�'�Ǽ	G��Y��w_��g��n䟃w䩺�$�#�+H��G��zͭ�
�.^X���n���{�En�Y���n ��/�=���u4\K
��]��Z;6���<��ֆ�ÕP7�t�/��͍�	4��gH�Cf��%�M(��n�f�S<"h�|��f�� y��6�T�U��j���	��s{��p[H���c�?�JD�Cݫ�P{�J�%1���X�a:]m��ÈK�id���=�6�& v�����L0�%������fq�x��&BC��{���_A��ұ@��V�� ��`�bЈY��(��׌$(��ER�F���-"��@�)D��[[٣�̏�Y�e��~E��:�Tx����U�Jr���}/j��������%�,a�Egz�̿!8�����s�lݦ�?k�1wN�y�t��Ï�F�I��G,RQx�}
`\K{
�.@@�� ya���!P>!np��P���m���?ɦW���N���Ģ;�=D?x�l�B�L�-P��Զ+!�����{�@����B
#���<$tx��v��`�z+��خ�n�����!J�#ô�|$�ZA�aГ��S�c���O���y���q3����ʠ���샰)��B��t�E����A�~��#l��_����;>��:�v��n���h�-�� c�xi�Q������Y�{l��S���b���v��=��/'G���s"����]���i�Tuz�, �fQPX/x�6���RK�٘���(	��-}�r��1��^�9T��F�o���>���}���B������uB
i7�}� ;������`�H-�L&1!��]���dJ��0d�3���(��dc���O?	�؄hP��1��Xw9��Nr�Q�8��b%iae��-4�O�꽁z�4���y�͢��g)���w/K�p�K&���ŉ=t���yE���]����k}\�d��F>9��\���������}��-Q`O�9l�&��_����?�uk� �0��?��l��L�>��F��tI���S+�+�EY����s��P�X�6W7�\*������;�.|9�t�3+�sNX�����nS
ٻ�뜳V�U�5�=<���(:sq���ԩ��ڀ�|�� ȕ?:[tU�to�Dd�s�L�M�Y4�vo�I��>J�J-%)��A�b]��o�ks�ᦘ���K���{����[����AfkiP��.j�AP�=��a���v!�oMtU2a����K�'H��97����p�f�׃�_��O0���s~X>` �����%��
����8i���\����C��.c�<^8C5����0z�>5%%š�3�JY��Y���p�mE3z�:��C����Ii	�c�ʦ��Iמr�R�����7�;���oA@}����8 ̈-��g��6֒q%%�)��A�\bf��塠�iǆg��×�B�k8��u�[�q�ž��樓����,
~�&�ʮx�07+h��rSQ�)��@���zD������P}�I�>G��2����V&�)������t��|���ث#�T�t�
T��܇+����d˪�LH%pz���{��h��4��Р��k�r;* ̾\`*�T����.�6\>:ȉ	0���=�f9Ԉ5���^��K1L� ��
.ڤ��� 2f��/�堜��b�a�弖Dj�q}�4ّ��;T ���68CP�+H@��8'�e�K��E姠������'��K�7��l/�Qȃ�p��G_�����UϪ�D���R�9�j���u����ԙJ7��� 6z��T TH^��~G�	޺;�N��vv�j6���X���[���@�bcT| kgi�� �iy(<e���4�2�;�(]�a+Z�>�4l�����vd���j+�����;>��n�T2>�z�̪��wY��Ϸ�*�/r�]fPX"�q�( d��Y��J���k+so���w���6OOX	�z]�'ྲྀ�0#��<�J8�<$,:xU4�r���( ����e�F�ܬ�䈇z�l?Mx�|�Tܑ��6��^�Y�yL���-�cA��8T�	�}��K'�u#�w��ܱ;��a�u���ߺC��i�zYc���+�}�G�F.A_��l�G��@�/� �H|�L2ar�3�ƭ�o���b�,���ʬ]LQ�-f�߯�'x�����|�'���;��i��<IU*��Uק����g��FJm�#\DT}���%Y�'e�����3�/F�i�c<;��7����ݎ?�_�~��o6�P��o_'� �9��=*-�ħ#�~��y�2Z�'��.��Q>Sr�,��m�1�zܺIu�,�Y?�jR�)��o_�����/��."}���P��-��k�a?p�=��rol�
��Y�iN�f�v/*�D���.�әY��7O�Q��s�K�Zsi��n�y�SS�ҩ4u�Y��f���=o����uk��a�Y��(K�l�"h0Ð�"�x��h��&S'��Xle]ӭ&X0V�M�O:`���\W�D�轖��.�pA�h�xN̨m�~�J�� U�g]��6��|ŋ�+S�|G�"A�����S]��N���\]�}-��K��ɫ��>�N����Oj*�����`���m�1Qm����8���h�	�,��I��AZ��B	�K]�Y(1����`�BdkSڞ{W�|� �A�.�YLq��yF�g� ���� �PI��fl��R�n8�+�?o�&�����e!��1lC���w���*��i�pD0eԮҍ�����:�:�A���U�ӗ	L?�\.�'�3$�o&�#
cSj�Ĉ��@.Kt"��P�n�4�͊=�W2�?�ZѩÑ>!��}P)SB���T0���X8SL`�%3*�Z!�)��r�57-����p?%@Y\5C�m<n@�1g��a�a�u�-	������8��`#����F�)��x�bCi���Z2�����w��*�l7_rΤ��0;[�KRO+p��y���c�9�6�$�����ЁL �Z'�	�S�;����q,� گ/��a(l[b@me��Ψ�Z2Vf+E5'´D Y�1Z�E�-7AqC�y�|��b[�a�1h��r���H^$�|H���
־��Ê� 12}�22d�����N����{�F_~<�D����֠�6OO��\��1��c_Qi&�5v�X���O������R��'7���|��8a���yJh���,H�Þy�	��O���%�3�j�a6��SwGg)�<�$��8-���j���a��:���Z�QL��%Z�K =��ɀ�'<�#\��0h�!���j9����?TMbq;����6^�lQ�/!^�9�DB������e��ҁ_>A�=��-I��?�W��N�nG;����ދև����"�y�[����G����w�����Y�oS>Wes�7f<�GV<��c&�.�D�Q�������C>M.i�5�|�f<��N�"��s G�w&W�̘�Ǌ�DN:mZ˩��$�ŭ��e��Y�����14�7�!�g�������d��t+�U����q'jZ'�������t+	1��G�'U�#V�u��Q�z��)8QReի���ž�TC�c�u,���e��J���^�(�,j���\(�U�*Kx��h���8o��f�-��e�ַ��b�Q�H�,�J9�F��|(���:Z~��Jv˭Ӄ�t�2ɪ�l�Y���ۢ$@�̈�eu����Y���0n%/�{���֮A�����j�?u([����:¡1��iX�[�9"»m�d[|�f""�'kW�>-���M�	E��x�Sԝ����6�)���/��=|�5�t�F(��1�}�A���G��8P�������b4�P��x�� @16eX��^�Ÿ��aA�52��njfԣ����f��Kp��1��
��ǀ5��e�B�|�׌p �K G�XL`�l�.�8��Mc�}G׮7��~�\�Aj������M��BGM����e�$K8�~���r';=C���b��u=╇Y�	g�ŊD1�����Mq_�y8|ȩT Ao��]�����9�D �f�T��*47��J���(:��+`��B�-��oD ���(���$H�/��U0���X&i�g�[r��1���!F�2B�d��6v�հs�?!y�7E�aQo׸<Z�c5p�{�{ֺ֟��|����}3����+����B)�~x/���j=��#�l�2A�m�G��ξ$���-��#�]�UH�V%A�qz�O ��(�M(���a:���J�#��W�x���Ё����n����G��Ү�h xC��u���O7s�?Sߊϸ��	�������W@ҡ�����J�lӦ������P�+��a�~�v����������hs�;^�Rq���/PA�?>��e���ɮ}����c<I��������_�/P��x=����lEd��r;��.� �GTy�j㪯ɥ;.&@SQ+��1�b�t	B0�Y����f/k0���P���ݾ5�����^�ư��;�ֽo��wf�8�diÞ�& ���ҾҼQ�P���I����ǰ1����tN�}Ϟ\��V�k�L�8�8��ުEl�R�c��f9CoF��GX�>�.ĝF9kg[�[Y�(�Mvt�v��#�@�8�j�c�pQ�������:�*mip�s�o�M��¼F\����t�6�P�,XCM��N m��6С�y�t%rh���<�6+�^a5�R6��~pF��"6z�y>;��=ـ���:�ǽU�ɮ'�Q�(J�Y�v�8$͗) w=�m{�Kp���v�O��B!4��_�/��"[;Ǐ�	�z��|�9�a"��o���:���q����\r;
����$�pS=�T�dˑ�ʸׯ7����Tb0)��`	�'I����β���'J���c�N�@��9�{!@�X5�v�[�e�1��|$�%�Bc�1 iO�R`�%�.�!T4������R5r���v݄�fi�@�w%�1�t�Γ�Y��P��Ek��$b�߶��S#��sX�+�'�l�<��~�;T�����-ũ��*	�]8C�����:�#�\�W4��e���L��̱���PM��"���}y(\�0�g�<�)x�;/"<�ꖮ�_c����ς8�L����?C��8b��Tz�G��%���~�{IG �ņ�[p�-�3,T(����eY(,#��7g�r�ݲ�p����V��H�����b˄O�����=�i��t�V��0����|B�mv���w?PUcYf�^B�}�W)��{���[w_&=�<���5?Ze�����3Os��;̡�ӽ�kOH���{
����X&}�%s��g��vc�NtӄX�謭]o�o�t�ܑe�����IF���ۦ�s�D���oI\���AV�%�	��O*�WO�1��s�i`�|9�;�V�{=�Z��(h)ע�Nc��Lt.�Y���6C�o"c�5K�Pj�L.:�<�I3�k� ��Ѥt0�R��lF
�n<9��ƣ^!t�W`8w�2̦T�|�/׊�9
�Mʁ>"<�R.W
��[;�,�4� �@x���V����[&(H�7��DOJ��{�3 0X'�O��e��!�M!�Y�,��S���Yp�E ��\��&�M� �	2 ��AR�T�U@�2j�Պ��^ȢZ��(J�����O�vk�2�{#�-�ta� F�a�/Q�p���.Ƥ�ñ���Rh��/͈)�Y�j~k/>�J���K�RE�&(�\�dy2�f!�ؑ7�T�ڀr�0�˶	�V�����#���s�?I=���C4% ���u�B�J��}b���!!�2 �9:��3v��� �dix,w��޼�7'��o	�t��*�r~_db��
�N�(��wǌ�#6=�=�N�A�}�0�1!��]�GR2�P��覭�#��{/�O9�$��Q^���\G����� ��g�܁�	,O���ܭ��U����q�b�-=�7��y`	�"$��&kBi�����R"(F�u��O���?|&�q�Ʌ���t���=���s�R�O��Y.I���wT?�u{�U�����gg�®�?7�o0�ټ|� �+�u��9���n�]�l8�%[[�����l�S9z�5I����[1rЌ�.�������n+^��kGvk��:� ���`�^��m�$٢��fK���&��dev�)m�L���9�4�j��ra�pL�t� 쥺˙rH�C�<Ny~m���7)e,*���M�,bm��J�X���.+��[e�nW2����g}�v�ܠ#1w�jYM��b�f	7$Z��l 7�\��S�'-S�D4z�r�(~-�V�2{�Ie-:/odu��ٓ�β�*��,^���i/��	.E��K<Rk��t���Cw},�S����P
����b9����^�#�^}��&[,����G�H
�
 3�Ϗ�&���Vt�i����=�ӕ��Yq���;]�\.B���҂L�#	f�4Q�/>��,�Z�р ȫ���-='q��^9!�P"@l���NI��)�=j�4��2�.& �]8k�bfk�/1�ѳz�gˉ�N ���B�Jk7ˍ���ac��i�J%דd��h)���bt��H����V�jA*He��.�1Ĭ��}C��-l ��\�����H$!W`ݯ5�xa�;�@I!�Z���A�Ym��]�7����5�E�y4D^�豕����l�ooX=����Iť�C{���6|6��'���篋��2����Y��[s���FA��b����s8'����w��)�����=UBG`?e��Řq�?� ���rl[d�mG^ Kh�2�4_m�N�{��I�����^���ꫫȺ4�-��SGJ>2Um8+��t���Wq���=�B�=��+®L�cU���br�.��yL�е�6� /!��:S	6,�[@7�y'��,��V㫪h�`f����<���-""b2H�����z�z̫��I��$s�0���W7�H#JW�����W���l�")�R�W����C�m���M���9y��)+��rᤃ�
���rE�3F^M�
�U�h�r���@laa�9B��Mnؖ��a���2��a�(�4�m����K3��{� d�e�#�X2�j!컇���)�~U���@�ɟ�<�@��䐵$т��Qj� sd��H�ͣ��Q'��s�d^���� �i�U��9��4�(��?!� �Pe&b]�X<?�ㄑ��@~ɜ�
��uX8�����t&b���(�D���'$�!�]|J����|�,�A�YJ�kǈe;��-�(|"t�M`�`S�*��&d�ٖ�&�}�9�^�l�TG��\�@mM�a�I�:��2ؿ��7����5�a@B�qO��X�J��1��qFވ���X�|�УE�?|--O�pEc�+N���ߓv�Eqm2
^h��v�+
�J�-��r��z�>�$�~Jϱ��-I�j�������Z�|���'��x���(�2�Wq��l��Ϝo��E�U��IP����N����z��e&�:���s Rue����l���H�;�r-�5����N:�==֠���%9󥮠!���0�7xJ��q�e􅶨��ڠ�����!�ꦟ�n�Y7/J�PQ�nm��=/JS��\��w�+��F�,�g9��T��ӭ�E�	�9t�(�>�9�-��L�&G�^�8<����������}�����TKm�4�m2��ܖ��f�uī��Zl�ԣ�̔�T~�k���XEc�cz�Z�aU�����&�s�}#0
/fi�5���]�[_U����Ɛd���۷N�$l�g@^]㨐�Ț3c��u����!��U9�N�s� qDz�8%��E�WB�y?ȉN���'�=�ɤ,Gi��)n���GL�����i��-�.U�eN�2|��	_����F�u��Eօ�e�!xBj"ZS+\*&��׆[�Nm�NbzT��mh���"��n�o���MG�6A����4duU���!c�������a�g�rS��8�E�g���dy�=�C �IS�Ek�% 0l\^A(�U���7�Ma��<~��dn,<O$@�4& ��\�2���=�>M�%��\^9��7�����"��g�>���'���[x�oӬ�ܟ�[��ϟ�s�e�K'��C���	:�9��v������49��Ei6+��`���/�j��6�#�����|Y�S��nssO�4�/k�m��V�/�պ둮�k��+�r�5<�Ҳ�J_%�)3�l�+��L=����(C3_@�.��d6�Y{��6�hJ-9ԍ>�"������\aq�UWZWݵ���ϥ���Ί�KA��d
3f�1�p���#sFF����f#[�N��f-������y�pR눠MO�;��Z	V�h�M�6�N��ծ[��q�m3;��|�"٢���&e�;g�;��J'Gnp���RH:e�h�����d3��li��j�	�A��1������R}�<v�Ȝ�%^�����a��	nM���$-�,S`��~19Nx���6{ь��:�1'���u��>����#9��l��� �����:ZHb��P��@қD��s����J,��� ��������������:��:�ȟ��	C!�k�%��`�,~��E��ʙAr5��u��cw�^:��8|2�c-P^�\u]�>}p,��`�{<���E��	��tc��s����4���=Et�z��<���_��߼�)n���r�glb28~v���ٵ%��Ő@b��XjC�\�������l���քO.ǜ�*�l��[��\�v�[�>I�� ����/����~h��r���u����I�Wb)Zg�}.uzH^�:�	ǜz�E���e!̟�4����KiK� k��x�E�c�����o}N�/�/u��S8��`���U �2Y����V��_^'6[�E�nj�33�|�++jqT�;y��:d�" 2aX�q#Pc_n��U�5k�<�̔A�"�Ӈ�ϠI\g&��}G"�5�ޟɉ�.K�����>W�x��aV�?�!@�&�'�-ѧ�q!��f�=��W%<6g�X �Ѡq�!�~��T����M�Ɉ�ZLJ�+C��N��5�M��a��{V[����8{��?�� 	K�=�o�^k�^Cҍ �R:�����?�_?5z[�[	�>z�)
OH�9}D�|�w������`
ݿ0��m�]�*�<��"���p��mj�bwο��ZQ���\|����%k���#�M�)K�q�z�춠x7�.K%��"�'�l�ƺ���[��j5DH�	l �V
-�(��3���Ç�����2�YԦ�ӏDo#?F���yd�������!	���ޖ�C�[MO��imY���.p{�<�/=DצV~������rޚw�{
$��%ޚL�H�&�5���a70��TcƉk��;zZmkmkןpf��r�̫m\t�S��q�j
/B����7�ѷ�^c���bL�����%?������rY��e���N�{|A�N�{�n�l%5o?�uk>ks��y��tY�_|a�?ވZ�>�u�R��Ͼ�G;ט��[���a�q��=Y���#�0�]����h���/]qH�D�)v�Vk�g3t������w��c6TѲ0~��P ����`K���ʽL�t_�T���g�#�O�kΚ�(i@�k�sԒ�r��S�~�G�&ayz{�$~}Tc��HU]mn��N��i�܉Z�^,.��M)Yu�bmC2�?��Hh�f��9�Va��NrM�D�lw>�6F��-ʽ{WM�ʀ����1��Ņ�ԞZ(�ڱms\�R������ϞWk�2W-�����,C���l��ܮ�#j���R�r�c�c�	Z���w���l3h����BH�݉q��7��*��H}���ˢ,>=�&��llDM�f��mSm�%6�,���� �!m";=,�N��䲻H���ԕK��=������k��TB���zk�=����{HA��w��P���Ï�͞�w$"V+�c,��\��!������c�q���{o�D�ԓ�_����?����#��ҁ�"�����/�V���n{s���A��:&���ct���������_�Qִ�� �y��
bu"���PK   ���WX���� 8� /   images/596601c5-6246-4a4b-a4a1-d26711181a9c.png��s%\�-ڝN:�ݱm{Ƕ���ckǶm��Awvl������s���tV��1W�5�k���� �����7Di)q�o߾���la~��������}wQ��V;Kp��ۯo��"j��=^�^D����5�U-U��Y��0�$���H��r�?�E"�~���;E��l�k��&0�k��D졲��f\�^��՜��9|m~\ry�v���QD�xW�	8�,�m<�>徽���x�D�~��I�'
� b!��!����c!�`�Ѭ���7<�5���'��a�(�p֠����XZg��7�Dl�_?���������:���%
�!WROiijZT�%{$Kۮ�2L)\$o�����Nѻ����6�grh?�UZoI �%)��Yiɖ%ii�I桪��|u�SA��Dܵ6|ΛӍvcuJa�Sp�5�����HTt�u�ѿ�T�ho��T����_��H�l������1��3�uw��>�-�ː}gmՆ���/U�����[�m���i��^��qP+_=�<}B%my%��]=+�b2�,9��@C�X!5��,�H�U#4�Z���+��+��:�Z�����	��r�[
Wά�Tewe�a���!6-����{�H��Z�銹����F���?ȥ��P���0�@�vm^g��[���Fz=��>����#���+W7�J[����O\k�	�]��6w\�Q	Ԛ۷�*����V�ڳ"j�}��F��4�[��<�[��Bj��VC	����ﴟ0�O~/>ʇ���)�/0�ډ��Y7��uM[gSlT���������(��lc&�A\���6�;��f�ԏ�h�g^Csu'�������a���io�H�>£���R/?OX��ǡ�K�u>\�!�a�������V�㥕�� ����ʔ���C�l,c��hu�gkq'��;�x�1��ʨF����J�Z�e�{ة��ZH�\@�>&\ ��'|%m��m�� �g�ZUu����������B��z�0�ڽ�ռ8*��JauL�s�@͔^ݒ8�2x�>��H;]��J���F1�?g<)g��b��Rw	��Ѱ�C��ԒW�� w}�޻���޽J�)�C�jZxi`D���Sv�;��BȠ_!W>T?țh��0$ny�3�^��P�H��a�&�U��o|� �o��E$#RX��>����xSG7�����}��
U�[�{f�ytO:��xz�A���#��c�����9�ܲ[�O�s�u���dʿX��l�s�����!�,��I��I3/`<�"$]�D�7A6~�e�����B�/��J��S�d���.+�oQ���;]������;n�4�gn�
�|�V���e-jS*�d�rc%�#%fԏ5g4��~�;F�����Wݩ�+�]W��]��_O�8kȤ%צ�*��''��7����q\ѕZ��]y�ZQV�@z�Fv�(Ң�z;b$D[uu�Xce�DM��b���T���󌔣]j]�L�=�_�Q�vGԕ�h�N�bz��� �O$x�U�!w��5Ԡ9�K��w��ЌC�S��g*�2��_+J�?�I�G�(���Xy��jw糆iXAa�����	������K�d�=�u�'�  R��X���W3y��U53Z#�q״N�5�����+�ʪe�4o�6ʽ
�L���G���	'�8R9�~qB*����	O��`��J1]����?�O^E��G��r(�W4cܙ:g��Dء���>���%�hp�h Gf�!ՈpB/��lM8��?a��蝃�='��-��)iʀZe���4��a��Iy	���ccS���B�y�n�w��K�5~`XWi��vr�����S��<�ً͑_��>7-��	ۢ�̟S�WpM���>U���]^�Q1���W.�ji�m+�e�R\�\DJ�5��e�F�8i�U���'�~�}6:�a�!����΅p�U Nԣo�.~�f�bf���p�0�qX�{��>@\v�ز)kjۧ���0�h6g���������'lh ��X�І{DyF��ǮU�be�"��-,�l�c}UQ�DЖ0���궅�J	>L�R�ҏ�R����ԉp 8�2՗����tx���>��}�8�H'+�ݶc�
z��	iV�5�9#���X�:��C��X�V�Lx/U3>��Ph�.��I	�g�P��>�FUH���t͈(f��k�Dl2��W/��0J9-�b
N>E����s&#�Y����Y��)�޲��YHc���@�54��$���X��=j թQ�8p��9g�w�~Զ����k�uh숍H~>�pp�}yE��q��B:(�r�lY/��G,��u�O��R(v�EXe1��'��KE��Cʢ�	#�#3p� m%�L�x5��]�
]�8���<X؜�yާ}�;�m�\s�di�����6��?�l�N�O�E���v��g,�	�v��ǽo��>�?�`"�I�%����y�3��hE�#:S?$?/WN1 "����4:�15ڲQA�򧼩&�V�S��܌��̳E�h�i��l���_�hl���j��>/Wo-��-z��b_	����c.�����&^�|����q������鎳��hܯ��px �XU��ޕK�b�T��(��wҐ�W�Өc��Ɗ�����s��m���و�ʣ�z�I���[�&ē���MA4�@�B����
��|�L<k�͙�-�?�!ת��E@;��V�I���`,t��A��B�_( ra��ѧˠ�O� ��Y[U������'�AM5l��5�ә[ߦS�%tS	��J8E6�X��!��!�ￒtnԮ�����P �%M WŖc��vl�z��@,��%P�=���{.Qʩ�����1Ű_P�~����&)
Ğ���>���c5�!���P3S�G^Jd�T�}l�CVH�O`{��Clp��fw)錑�+=�g�p�����O����8�_:��ߨ�o��vM>>�ƪ���?�\�խw�\���bF�$B���r�S�$B�U2���B^;���6�����9|A랓[w���?�F�&?��pX9P����ƣ�'|W�^f�:���9�y�������q��^��&�x;���|�:j���c��q%r$Wdv��%�G0M�m�gٰ���z:*ķi�u����R.������Q|��uh�� ��.}>���:^aQ�>zP�W'�W�q�ۤ5F���C��An����/�Qlڣ<y�����U�3�{P�����q�֊�w�)�IM'e
iƨ�+P�o\ш%B��#(�eJ�:B��=��YɌ � ��1l�X�?)�yUj:\���	a��F�B����NK��R��b¿@v�|�L��D:5o�&n=cE~��3.����ga��9���M�z�D,9���ݕ^N�8g�����
>���0�����*����v���9���U�(��ɓt�v#rLN��3V�z�=��I�ý���$�O4���x�W�1��D��ԗdQ$7VH|FpIc�����������;Ho�/�O�@[� ��J4!'�;A������55U���Yތ���K���k�4��/��n�����&Z���*���cc#��Ĕi��������4U��y�[=�<6���x�MFc��.������
�~�t�t]���+�'U!�<���d�IP����mJ�4g~@�zA��)X��.��ɻ�P ��K,� ."lq%N�8
?n�u$��9Z%1�<=����I�TqS9��[obM������M�2���^�]�+9��'T�����`�ϋ6ƞ�pxF����+ӳQ�}�Wdm��]������5g��5g�	v�Pvа���j�;^���JOL(ȼ#Up�r�p'�iL��h���6w!@/`�5Vǋ�D;k��� VYI��HT� �.�Ɵ�8��!������;f�Y��U� �|�Ѯ��}��ova�U_�iB�0�T��ݐ��A�@���h�z��hQ8]!Y)����_z�$E��m��ȸ������u6����"a
E��K��$��^b��1�J���:c�E�f��зr.�ja̃����H,Y��~�1V^���ݩ�OP�GG��
%t�Y�p��2]�^�f��N�}}LG�ӣ��2�ꨬ�&����L}�n�$/$\���IV�,d�.y�K��lY�4o|���K\�}�oo[�g��}=��ǳQE��D@߰�g������9G�e�L4��$�,����^48J )|�HY�0o��+?���N�'��o)��/�x�#a��
�K
��;�E�2�_�|_8	����ʂ�+��9׸��v�"��H^��W���\@_m<�y��> �� ��A#qo�tr`�}�������Ѵ
�?�vޙ=��O��w������e����h��sym�r<#����h�5�-nК�F���EΩ��藪��g���%*��ɴ��F�l�09m֑���!�C�!-}9��1Xž�R-ioB�H�n�;�:R/7�Fʣ��kZH:2�����ڇ���ƫ&�hύE��CM�������3���D�\!S`o=E��/J�u��M��<ʪ��,�Aͷ
kK\i	�k�ڔ+��^J��و�?��yY��r�>s&�ɠc��?�#感��1k�h$E���.5d���)L.�8'�v2�r�a ~�QN���ɽ���pR^�M�T��脞��*�6r�o���6�l�BW������Go��ۣ�����7�p��vPn�Bbҥ<��i��3��1Ie����ͫ��5D���ey/L�{k�OĂ1�/�%��i�'T��wi��O|���i��
�ۤ�Z
�ܸ{����d��q
�4u"KPm��1�#?��Y6v�Uh͝K(�im�����f+n-U�$ʤbj�lݜ0�8��(:�b:Ϟ4[��x+�ArC8c�Νn�b	u�覲�ڳڇ�t3�3�t�f�:��yG�K\��z�f/�m:��&\����z����G��⿊ˎ��G�z��Vp��HF�}�*+;���:�춺��^�i^ώp�������l����
[�bA�!_�o&K�M��I��r4:�K%[�
w�b����v�?d��Ȍq���c���;::��;E��ڵ@�(O��;7���{��X&�ư,��<�F��@(����Y��#n����{=!�7�j ]F�ttyu���B�����%04����ۋn��PR�uJ7*ѐ������G�G¾��!�5�`���q�
��A�����Ն�$&��d�/�	��	3n�?�
�ͶE,pVY��0a�����kf]��Q4(�p<�$�h����m6��)�
P���<lb�O"����������w���[E�醰c�O�Z�<��3¦Y���h��Մ���8�g�5nW�?�N��7�*'�wg�}b�>��4����E������Ʃ1�BxĿ��^$&���`�O	V��`l�.!�M�6��cU��_�1t��0���X߫�-6��f�՞,MЎ�ԃ���˿=Bi�a��p0�|���I���1#���S�s<����.��b�d�P�(��]�|)��MuJ9�`o|}�"��������Ju��a���@�g�c8���x�����k��w�#��8z��v�W�����m�>~�2\���Y]�Y�	�"�����l�ߦ�����O�ַW�=��cO��/]��v� 7k��ӈ�I�f��,����8t�Ytnh��x�%�#"}4�������JqU��0\���wRJ+�W����ll���OB	8�T��KA�yC]i�V�X�h����_��(;�Qn:\��K��QY�����5�����7�K"���	�k����ڞ�.�2kЯ���)K)�|�ԫ�Щ/�2ԡ�
���_��j��8Cx�J�h�e&\�X��Af�U7�M&�?I0�d�1��X��W�7��l����>$��4dAE��bα�~��Э �q�NX�W�ܘ��>��4 ��7���v�P��q�lMK�,�}��H������^���7�,i�c7x��A���������l���&q6�	��:�)+2a�]��qKN,y�LZ1��Î�u�7TV�4�&42ISʖ���|f��Bސ�L�4c:��0�/�<�t���ֿ�a���
\S[ĉ��X���l#ť�5���t�h�����,!:Q=�O�7t]RO{tg����kz:9���]Xf:=3�K�)55�'=//�9�X�1U3U�i8�I��r�8�ED����rtyS�Z0ĥ���������1��y�j��d�t���%��O2w��gMKG(�&��G^E�$Xc.���V�3��?\��]8�f^Kj���"�`j��2*f9����+!=���Jf�5��77������]H8�2#��QUU:����t?�h-�lO<�O�U��,��M*j�>,)L@a�3�ΓV2��:��=���n�$�2X���C�N�`�2��\)8�W;8n�ew���Ʊ��b��Yˍ�n�2�k��4�B����S��s��o뢊�$uJ-4�,��h�^���x��h�J��B��K*8lmk���66?k�uU��bF��?!8:�j�3�����o+p�7m��2n�*�%�ό�g����E�9�SZT��[>@>}���]�<Un�T1}G��>�A'�8W�%������h(N�����Ƶ���mEU
�i⅝�U�4.3J�j�[�#�(�"�_�7bXA�(��d
�Ƥ���D�	E���v��I�3���4�F! ������橣̅���o�z��w!�|w����籴R��Ѷ���3�4y?/�N�jp]���Pz��h{D��kii%��"���/�Z�z����z�]�{~>�e�6��-����c�='uu�}������j5��@�B
%���D\���/��T���(\CAe�f��t�L)^ʿV��×��i�֍b�]]�
	`�2���5��le���ז���U+T�����)����9�g�3`��N����h��ba�"���F�˂�H�P���1�:̽���# �Ȩ'&��8�I�	1V11%��E4�p�S�"ggX/Y�X뉣��0�+�2�͈U�=�{N#鸋�"���R4u����3W��	��B�D�P�V��S�iB�L�;ޙ�B�|O\-��.ߚ3��i����0C��$�RP�u�r~�<��� �԰��D��!�*��Yt(մ]�����ٜ�
�jS��dj}Mz0{\C��Ȩ7��ew��Q��{hӟ��ڻ=��G�G��Gu �����X����"��az��Q'N|�	�?)���F�����6ɲT��ja�!f�n���d���Q���T�ݣ ����+�zm�󲷎�����?�����K-�ᘛZ�`�K!vr+A���ywU,�xVy!(vE[}?X;�E�k&/k��"8��?�*~�.$d���Q�Įī#um=.O
�DT��p�U@?@vܨ�:�}JD/SB(;��wP����Npy>8��_��U�?��q�����not��{��v�������zP\�d�>w�n'/t�m7|��Sʣ�����=+�9���`�KNE��'f���ˢ�b��b��z6��X�S�n`.���i0��$�#~��S�$�^^Sa����QE�����)yy�����'����#�;�Eq)����2����Y��c{�����j���a|jF����H̅r��\�f��(!r��f�)�U�&��8(����f��Ķ;��)��KkT����O<�!��;�S<�Y@�lCJp�'�j�I�	�13%^l��t,�]�߄�(��CZ��ʾ��, �@�yKj9�l�H��,��$D{��*�6,P�]B}��8X�I��ñ>�%��i��>񍺳�RJkցR��	~�y��{������o����t�g�{�����rvZ���X� ���|0 �u�qf�BޖQЄ�J��YGo��5c̵���M�� �E�TE���`)uR��[��|�.1�S���rLKz��=3�U`�Q���+/����3�uao13t���$P�̇���}%���xYZ]���|ݛ��<��� -|�Ua9N��X~���vr�qZ^���b�x��Z�_�ᓖE�㇝5�Μ�x}�/p��{h���Q���ߠ�	w��:������������ɜ-�"����cD�+�a�ȣ�i��j���1�Q�~T���%>[&�\?H�N7&��K�P7S"]���x���b4ݰz&�ʎ^"�7өIdYh`O-
��2�����㋩�.�(�`��"t;~*�zi������CJ0���f��q��9]^�CRX%����ňP�E�ttt&���z5V��I��Z����n-ҡ�ܢ[B�4�=8�DK®Sq���;�G�LĹȍ�XuJ�,5��1�*���a��r.����ޚ�51�Lp�R��J*bB�'K*� X8Ú,2M��X�A�t��
G���Q=�h>S�'>�Dt�G��+	�"S�)`�R3aϕa�C�H� �=�w��i�4�L�V��Z�]�>B�n+���/�2�|n�|NR��a^5����#�H����4s|�ܸ��?�i~��m,z .��]8��S��	�����e�BQ*M)k%ĲO;��%��R^����*2���3�ͯ�:�[�Jt�H��z�p�jpg�1.2��DO��iO�Q\v��Kg�gA��d)V�)���t{�B����!G�#{ب����� �:� T-�Nuq31�����ԔU���hݪ���������.��S�c���|.�3�����f�U���l�iyӋxqxp���j�a�_�歹M�17�(Ph�n����A�M�۰��G�����l���9��2�N�8L:��4隻h�d���Q�1ʇ,�8��YS�^����h����Iz��JX�8kIYT����ov/z ��@U���8�Ӧ������U����B�S�+E�j%d]]��;�x~Ҽo���"�4rHjp6G��@� o2(��wo�LERx"0-�yd5�F����H�F�Lϭ���WO�����W��ǘwy18e`��y!�yԨ���֫6T�R 1_kmK�)!�d#[1��v�G$-l�(�A�-t�1�cH��
83e�/��?�v=����~�GK�3\�Jt�%�E5��J���v�˃��*��h��'OO[7u�ڽ.�b���nkԊ8�3�y��D#�u"��ƶ�_�IX^M�Y�[�t\�ܛD�Sq���%�
B3x���ޕQe8ǣ,.�kaM�o�d�b���8� �Y+���	E�����;�0��S�H��F�up�;�Y{��n�X�+���y��׸�L?�cf ���L��XMj)�F���?%Y����k�fP��V%kfv���zgnWf!�d�أs�H#'xiK[W��*�?���/��Ihk�������c�����ᝒ�������,����+�gy���;�tiǇ���=�o�L��jy&?2W�x��8�=��:a �3c���PF�U�đcRk��8ǘ��
K�lvZ 9%e˛�����*�L0�d���"třixK�9�#E�4�D�m_���<�в���2�kMQ}N)f��D�P�㗔9�E#��U#�5���M����4gaW�q����J���,�H
SuyEl�̝�;�3�!�H�o�����Ņ���#$;s����u%jdf�E�������@✿�RWp��D���У�����:�q�:M͚.�uVڢ:h��*D^������g�ύ�������/�HHc�[����5�Y�r��v��,`ӮQ��@�,��3��ů��������+Þ��<�G���f���W4���q���ض��:M��eo`6���rIj��ל�.�����F�&G%��u~d;N�A�Ɯ�S�G4G������%�/,i�Z�~	��kޜG����?񂌻(�R"�j���H|�?O]��܎.��lc��F��JG~b2v���{�Z=h�
��
ۄgL��3_"�u5X�et��mn-��̲�Gy�
M���n�)��P�m��E�Q����ke�e	8�=3�����]��\|$�q�����Ojbc/C=>!|$�k´QMF�Bb���\�<��݋%T�ZB�������V�ӈx|г�����F��7�]b�ađ<r
�>L�ʍsS��e��s����bIb��U�JT4}�^��4��G�y{AyW��;z�nϦ����*K�4j���$@���q۔��_S-��
�j
�b�w�@S��C��� ��yIbLS��%ye�~5��j^�w�͵��(=x2K����cOۭ`D�r�~��3�������`�n�1R.�-��x߾B��B�L}�S���-�Ļ�\ xm�~Q\���@J�������}Q���~���
��;ϵ8��B��7��Q��{q��_�2N�8�V��bm�,��qy���xQ�̓XyQl
����0���ȳ��Y�н��C�����]�׭��[_s�����ɷh��b#��+�A|C��迍�i�p��n��j�lꔔ��	>�6��Њ���}^�>a��H����ͤ9�%����Z�&�%��e���rrN��a�:���l�5�-�|!�/��ȯH������!��x�[q�V��Hd�{r��4�e�\���* <h�ɸ�0�"��g���q�`Nh舎�a�|�|R��Ϧ��O����&yn�ӻ�؋/�)n[��T��,s|j�[�bu��X�.
�r{��^߫�y�_㛾�K|=S��:ۺ�NvR�W\����K��`V�#�)�P����B(ύ`�������#F��݅��=�OPV�v�Ę�K0+�t���(����Y+�����5�P#�$EC���v=�1�-�<��P��j�6��R�d��@ŎD�Ny������,��U����nGX����@��g���zJ!���4`E�J|��"���qJ��Ñ�9|�6&�+��1�T0P�c���<B���{t�#ON��� ��"�6�] Z��z�
� �e�Z�9��y���$�$��
�Y�� ���޳�y�q'��c�xǿ�{)�"ƞ�P7>��_���<L���wq�ؑ�M���=�Kˏ�N@��H�<��K��ь�ip���-t���q�H6-l3}��{k��}n��v�^b�}�nĩ�3jYA�޳�Y��G���bo�/�n`�0��ٓU�E�JOﰙf&&�r�J�|�Z�ʹ�����?;��o�r�5K���fu�c((j�)tg��j'~������Wz�opZ'�Al�d?�^���(�bo��F`�|���f���a��<���G0E��SZjc|	���K+�@��7)@˓Cr�VŲu��N���fD4��.8���Ua�*�ٶu&��0. ��g�y9D�h7�m�]�,ت�ߏY1�</�j����Od�?&��w��S�GG��u�LSp���M�@����W��Z���t��q�iD�>aӪb��}��i��R�*Pd�nⲡ�b�ˮ���4�i�ζM���X�c��%��Mq>d� ���7�#�N���~eT�'S �Ь���#�� ;���@��	�N��o��n�J�	�ke5�8=���k{�������Q���+.�E]n���v+1��k�g���p�-t����:L&)��0��#��
O0���I���b2����+6A����=�����nY�?���-�K���y�Fq�ޓD��`��^��ץ�,��T���ͽ�^y��WY���%�����v�C�^�˟����Y��;��wiI�ėq�~����V��?j�"��e�]K�-)\�� !��=&!�����g?����/��)8��+��#��kSK;��6�Epg��'EB��ɂ��l�Q�k� w��K���|h�z�ƒ�<X��ʭ@窆�ǡOU{\�C�R�F�겳p�x�Zy�2�Sɸ%+kk���MX{���Ur����d���� v!���I�G����:Y��iC޳�/�ZBtx��CW�)K.���5gAN���n�ZS�I��-6����5	�^�31�#�2��q�2a�A��g�pGnÿ��&��	��5X�a�������3W���A�ټ��I�����'_(�~0�_��i~ly�������;��Q��׹� ��w=�k�z_߄�`-=/���z�]�>�];�=�n�]�HPXX�L�i�<aי�MK��x87�2�$��Ę(��w��UѸ��=/{'S��Ժ!�Pdr�<�I0i���U�B�0 ���9{�������l0l���tx�0SĝC��ŗ�%1�q1�
����D.������{�B�A����zƶVw��"U�e[���c�~ʇ�e����q��*�$"��V!'��s��Q�R+��Q�G%r����I�4�B	0��{şɥ-��q>��r
ɨ�R?����Ѓi b���s��+��il2uBU)��C+�{S�:�d~!�]����ds9�hw��i� �������3��_�"�¬YUvQF��SQ��q�.6]yΪ|��sT�/� ��в;��*Z���?�}��ٯs)~Ձ>��R��M���<õ���kH�@ͮw����ޘ�R���</$X�Rz�|�i���v�����No6�1�U��ٳa ��{�`qe%ՏJ��J��]N�D����>�f�7 ����k����_���]�A�v�7��R����q�pNp/%G��b	&�)r{�#+%�$1�o�{<�/r���+�:�wɾ5���Ԡ�8s����qs�v�W��xs�'��=O�W��-w��_�*r�3�H	z�����й�x��2���w���|�%2���#�y�J�r.�p6gC���k��oU.�r�[Jl�}I�����1�S1�u�f��Q4�BI���Qf�ڈRlt9	������ꫣB���4�f�/�A�M�mѤ�_#���X	@�
L�nR.�����uB���������{�˧Y���
*�sG{/;b���-?��o˝`�F�GB��v�;�|����X���1��7�*�Y����4��'?��� �T���]��ʚ/�
�*�uнsW�],.^u9\�A��L//0�|�B����d=��_R.`}Â��w������C�ʾ#�5R=�ʪSԲ��!�Pfc(��"YQ�u��&���[ת���<r��J#�3��Z���/#)V6k����)��v;������%��pݿ��x8����[I{VӰ�B�
������1���)l'f�/�g�J�	Q@������+�d5������6�29��5@��GC�&^����L�!")
yčv���mt�ch���j��T��׮�����D�+eg�2�3��o�Ƅ�[��%D[|�L(rl#ݟS�
=-�V��5��=�j�cO���	��kůkh��������>'�#���&C����mo(z>t,v0��<r�����(7����.��ֆ8��D�E�t��%W��NʕFj���n6��.G*WCqX#�nb�frjx��Y���9�"�D�N �7�0�vs�k|B���f��X��5���T�������o6suA4�K�[��{�����9rS�	���P���k��݃hm�n
����0�v�q����4n]8^9N���W�L缾�Q��Gm�"G��\���\��L���%�t,����6/�V�Y��cn�pn6O��-ￆ���y����\�ES]�C��A�c�=�4o$�w�R��a�5κ�$I��jq����@�*��?8�,y�3]g
�U�"������s���<�~��D��K���ߔ3zD��{-'�iΈxA�%t�6�!���N	����ݜ7�6?$,{�hiʘyz�y���J�ϸ �m����ot($Uc����r�~���yb�q��u����cМ�^�eM ��q�ᢕ�g���2E�r�ĵ\��#¦�(%���Ln�C@V�f?�>��c�s^;�j�$qE� �/��A<U��ҤqY�-Y�+�"0��V2�u���N?�K�f�`0e������!y/�{����d�H�����7��ɩ#��t�Ұ:c�d�x�ʤ���w���V��\��P몓�u\N�C�4i�<Ib�*X��^J$��sa��8�#G=���{]������UI7���ck\w�hG&�X�vWl&vƯ��Vvٳ�(���`�!(�!9��a�����_����<�={#�n*�A��@2�������$�M�\H������KE&�� 
��d�=v�-�?J���׹���H]�5W�k��Z�92J�� �!�Ÿ�� a�OK�mYPOt�Ҋ�Ռ������������b�aQ���b��1�K�M���t�<c�Ly��NN�R:������aƒ��P|��:�uw?��N�m�&�p"��o�~U�,�'������ub���/>+>8%�Е�)ED4{rtp�Gc���_|��R�.������L���J�=x�T:ƩH9��H�C��Ti�<<���&��s'P���qKVg�}d��>�q	��u�����#��͡?�R�E��M��gW���OD�qXM�OD�@�Ɋ:DxC�
�xB��`���	��x>���WB#~�|�x��ᵞ��f|���W�L��&�u-�b��xbB믨��
�USfD�0F�+aգ?�\�΂�U-e0'Q"J���F-��mI����� w����cm�'=c����w{|�ET��x6EB$N�<��2Iy��I�,{aҿ^:{"I�{r!
���'��mSޚ�Ł�l8 V��~�ڌ�9�-�1���hjxq�IR���Q����j/��岹1�.�N���񵵓+����,��&3�U��tI=�3&ka�ȭ:'=�ђ#���cBS&��~�g���JY�|���U�e((?��{@+�<ގ �,.#٬a��WK �tL�~�&^�2��۲����n���Vx�h���
�u�_|+��D�B����P����Ԇ�p�%%�˳V�Y�0����58�-Ռi��X��'k��Fm���."ҮL5�ʧ?�q����&J1�浔~҈L$���$XOUp3��HYd�`r�����tl�64�,�m��\�~����]u7݃�F�<O�be�zu��P
�D�*��hY�T�=PL�#�07뚌;�u�E��ۀ*�X���Dx�qE��}<Ă8���f��7E�����n0O�o�%��~Cرdg>3��Lx�@~����_�=�"�&��x�J���u�a�����aFХ�O�������ۗ��-Ȟ3T��D���M�[�V9������V�Y�+��~�(e4d��C�ĝݏlX�*�I��D�p=In�|��vԂ����.;{;���pM߶���j)�:>[����ͥ������<<�l�={���
����kWҊ��W�'�Mۀ��o���g�J�?3	=��9���&��M�`�e�N��m� L���T�-9=�N�c[0�$��4�R��ˍ���	��ܣ̇R�x�>�}V�u�\�Da1����5�3j.��9?^��ܭ��a��y	#���o~�_[�P�Coh�����:�� n}3��<v��ZX�l�u#	�4o���(o�vd��T�%7�S�'*�g (0Jw���9x!��(=ȐX���B��&���>s �U� ��,GK�'�-{t���,]�'ʍV�8{��tx�[Z*n�5��
��q�[���j@�n֮6��Y�=k��3�-�7�����������5
˂'d^I�
���V�SI��  �J��1ޠŉYy�p�:�ж�N��d�GV��F<ٕ�c].`�x�N4��g`�9'�hJ��p(�K�*�e�[&�zo5ej7*a)��4�o�R�: @��h������+I%���ț����p���cIz-�U�*�'EP5v/!?�����}�χ3�1��B4/զ`mO8H� 4��\m�[�&�����a�������y�	
����؃W�WC��J{e�-m���H�mbg�P� j.��@n{-淩�.R*��1ȍ<�LFx���a��s�/y���%P�8�aoۈ�F����g��.�f��]��&�/��SBa�����9�7�e��5S��ܱ��pO�yE�)^1��>�k��.��-�_����|�w��0�M��G�n���u ��)��
�r9�B��G��?�c��!�\�^N�I6�!5�L3�tT�d��A@����F\��;@���fěk`c��$~	��9������f:�����X[\�}����Z_\�~����<4c���}������y����ڛ�`R`0��X���H�9��3��H_Q��H�<�1Q+ƓQ�0�X>��(�D��Kb�^ٗ��d�(��˺�7�)�|o^�%��U�����(Sp04Y�����@��=q�2?&��L�'N},���؉�n������6~����Γ�Sl�Wxd#��7�Ǜ����'>����{ۘ�bt�D]�2g3fMkml�H=���,5/j�'�x�r�5;R�[�ƓުA �SY2C��k	)2J>�׆��Y';���J��ɠ̿"�ѿEE�5��n���Q@���}���ξ.(��!jwE��'�4Q_X^±c�1��$��ir��투���Rơ�ox��
V�4�)8q:�9��"!˻T�B�T0i��S��Q��c�d*.͙kBWMr�B(q0��gJS�\�(�o2���mEC:e��}T:s��_�,h�/G�p�����(��TYq��@	m& HO��Ij��,�����r�E�ӹ�2�5�,�H߅�EqnLsCt�J���c��G�$�I��)%A���v�>>{����"w�����3z���t��9<e]��!�����v����Ջ��F�K��St���NN�Ŷ���G��a>��P��o%��/���ZF�,���V"S�ٚ�_�Y�W_^^�� ]�Ȥ5-8���;S\/�	M�D�-1�ĦƘ{�/IGTJ�b�ʔ15FGO4	&5a��ͅ�ˤse�{�_?�<�P�Z�ٰ����f��*���������	t�<;�&Q�#+:F���g����(�&Њ���;b�hT�ql�_�������{\��'��wQK#v�^h��D�^}ND�u�ԟ���ʧ�|��L��z��C3����'.����[#k������P�#���X� �Z6�gD�$*��JY�*�ef�0E�ʈ3zXlR/N��du�喝���b0���V6bLjd�b�;O=GF�l�.à����VF��;�(S�"�d*.8Q�u�&�X���F�2�ʟT*�`ur����c�ͅ���c��+x���յ���b��\9:��/�G�x�²���U�2h>�x�f#ؘ�L����Ӵi�=h4�u�T�'��O㭷��D尻��ф,fH=�#=e�w�r��]�Ӭa]@�"�a��ȅ��,�����&P���6pj��9�>;C)�����a^��&z0
��+�4� ^/�@���4 
K'�؜����<��,}��4#و�L���a)�*��Q�20["E��	\�X.������.sZr��'Ʀ$���$u,�"��o^|�:RU��A`a2؇m��1N�H��LzJ���uW�/�Hٳ�W=��FuZEJIsw����5���z�s&�c�h�"&ASX�u�0N�98���ގ�X-e�EԩSJi��'������>��R��U�אx+�8�� �ܱQfcD~�˗^���+�	��ZN�f���h	Z��~�{��Z֥�9N|�׾����̚�z�q:�$�ª���M�Fo���HD��SY�1e:�L����T_���ݏ���Q�\�Ζ�:�:�G�m]�e�Wꬫ�2<��/��n7ɠ@H��HFѻ.�(�k a�-����i�8ǔ�'��Z� IW	Zw�����9ƹϦ�WY��!�m�L+p_	+����|E��L�+��\E��.�����m�=�`�Ւ�`v�:u���>q���z�y�C3���w�����oM�����pc� [�c&9J'�=I�K�QL��Qg�����r�J�[��đU����V�E�����9m�f�s�n����ņ�T�:�y9����:�F
���)�D�9F{��=F-��O��Y��!����a��+xfԷ>:���=�H�ή�x�9�\y��ۿ���'Н���P��f
�V9�LQ�Ub��vD����/��DI>�↣�k�RxuJ�p4��³�(�?�]�)Ċ+W����B �b0�["�dk��BRZ��R��=�DUu�{}����]�Ѥj�[����1D�%��0����}γm��Z��P�Kȉ�9�@���N5�D�&�qM
���(� 02a�����~=���؆�u��U��y��AlH���[Z�,
�#�r5PQ�".�V�$��ܾ4 �]���Ӓ��n�d� t�!f:XEA�%�(bĳf�C̦Cx>��S�;���5VYF&�\j�!?K�q܃t
m������p��D�+*P�x%"�tDI5��K�B�YrL��Pc���B2�J�'/<���F�K��o>���v�+\ߛC�c\9������҄�Q�ȳ]ܼ����a��O"Z�*L����>6B+�Y����>���_���x��Iч�!.2�c�i�Z���.��¶0����4P �K���BO&Ҹ���f��@�D���J3�4��Lg��졂��F�FO��\~��%�n��QN7�no�F�aA�dߍ>�&Nw������@E���&0Db�P����)7m@Mo�p���(�IN��-�r���:�F���5�R9���|j��ܐ/Ab�;�1�#�H�봱��r�ԅӟ\j-�� F���P��̓��=���ϼ{}�w�Lq8�8�C�D*�v�H��b*]`E>C�̈́vϼ�ks�i�0p����ގJ,�	�92��Q��gI$!�&Đi��4��lin-��H�db$��$�1�z���twѡ��đPŊa��ʺ�A!ܘ�0q~�S^i���e"s�=׿���Ozx�t;������p����[��Y�I*��eÕ41
K	:!���Z�8�$(f��>���c�)_�g��9�fs�`!0f�݌�y�9ﭺ3҉S'����ap(����DE*^2�����B�BH�Jx2v�q|���8�ks�'`ۺ����R��zN""��� �@���!kB�F�\�a|��n���#�ZDM���q=*�A�<��vP'��˫�P�C�C��@Q���&�o�L����aIg���(H;=����h�����M=�y�|���5�����\8�nR�1�H�=�A���c��2BUY�yȃ�f֩x�|	�ñ���A j�d4�EE�x�E�c�)�3�j9G�]�4��s�֍}9GƖ�@c;�la<}�|�,�����v�k�}$�
��+)(^S���6�{�18��xpe���9�K�߁Ocfhw�2R�R�.��.�}�
^|��iv����(���8�w�JJ
��k�b���H��>�5���ht���v�!�Q6� ���Z"��)�2E��)�ؘ��</Y��?�?�Wd�jo����%m�+h��!k�<�������9	�K��C��)<N�N�q�ghr�j��9��嚟��z�9��͚?B�qr�@��Dƒ�s,1�Ry�.�C���=̵��u��<q�=}�?�!� �{��v0����7�>��{װ}0BZ���I���<s���PY����4���q�D�"'M>ƙD��B�4م�+��8ue<�!K9C�B�VH����Z.5���Ɉ��q'��g3�M�3������.|K�V�}�Lg�&VN�-9�l�m� k֟�be1եK4Ƅ^�\M�D�Ifw٦�;��ss�z��뿉c�Cw���4�ʘ�K��¡lI���$���/�DK�0"!S�M���d��c����S�'�h��G�p4J������0$,ݺu��v0�d��Mm6e(ʠ.�QcƑ�\gY����� lV�0Z������4�g�K%d���(���^�!e�I�Bh��=��μ���Ѩ�Q �7g;l7����2G���h���ji��'.3�[q��1!rF(YF��D(O�Y��M�ɂ��RD��<�ñ���|O�vavVZ� h�d��{�1큽B�t�~��l��x�bd)73�<4#d�3�� �7,��������`���х(S��2��K�{v\a���D��R{mOg%�(F'�}��/?���f�U<����8��>�K�}~��	��Y��)��6w�C6�F2څ������)W��UcK�����c'q��"���zo_~�2�G>
���)"Z$X�k�Ddb,�H�Ock�
��$�6���0O��v��G=?�9"�Xd��ɣ��hܸ6�Hd�\��zx;#��U�1B&+�����<�i�2��{�C�S]w�����S�$F�g̺ں���` �ޔ@I�r������[��2�ׇ� ��@T4�::R��H-�d�F���t8�Nc�r�,EX�_�9p������g}bnn����s�C5�;��oz�[_y��m���A�F�{�Bp�b��:��H��������2���o��XX����<ڝ��o���<c��y��i�ݽ����h�
�g�J�o$Z�e�I�8؅ȕ��9:�P-2s�lB�E���r���b�/�@��h�u�fԒ�9�G�@�5-��%���xŎ6�;�ɓrB�Opz�����w�ó�,ڝShͭ���fY������:�=�D�K&a@�cW;�RsĄ�/^�(��݉P.cl%��r��x��ǫ���XYY���L|1����-)Sa>�^��.�(�q����F�,�bT��'�]���No�	��Љ���h`�O �.3�W�n��z�E/_d[��3'�I���T�J.!�J�Fi|�Ύ5���8uꔠ�����Q2�f���"}:�X�,[��� q�G�#}rUY��Q�LF�Q��wºJ�ὄ�@`�ٔd�)�vnbwo햇N@"�\uJ���N0S7�D�K��,M�ܓu?eu�ԩ�r�Krq]mu��8/��*k;O�ܔ�k�U�ח���W�̚�[V�����	�4ǉ�'aWc�g����1qn�씸���ˀ�2�
H�p�	F�1<��x��tv��a��H7*:�_��*�l��e.*�p���e+�_��w�ΐ���k!&��<g��/r�l�g>u��Q'y��%���c�YM���T����Z��3��zz�V	~ aT�-�J{S6��t���ق@��8�&��}F4��ƼLޗ�!)6T�_�������ily���v�:5��t���)�3s�Mg2	�đ4���2k��)Htťj��F��)�E���k�9wѥ��ř��(C2�C�ȅ#�Z��X���4���3�>�a�y�C5���ѓo�w󵷯����!��ڤ����V�Bb��P���޺����=Y��īK��	��$=�[P1�P�L�(|Lxigk��Wnawg��r��$Q�5�(tvU&2��%���D��w!,Yw/�:bh�s4�u�XZ�A{�r�!R(�,Be�j�8٧t*Lnא��{���ǲ7��B�3��{���g���u~o�����B�#Q�-76�g�e[��t#�-��y�b�r��_�tI	��x�5���d�<7d�� !E1ʵ�}��1&N�=�]q��3ywg_����J[���e��Ls+^[�� ���G��. ���+R�Y��/*C5l��!�n�&$���a������)�X��~����fi
���4d-v�l��TrČ�5R[]]�.���@�.c �W��=�hiXh�Ln_f猠1��5���q�;�&�όZ���4���3�w�s����.����9Z%�dz���mv�<HY��3��\]�9��Ld����o!�5(_���������6�W��N>��ǐm�.--��c�F6.�$�ШӨ��T*q��(sF�t�N�<ךb8yO�<Z�.no���Gᮡ�}��#;��O��oc6�������l ��~���|K�r�M�+t�̳�R�B8�!�pd�i�+�^���"����.,�%3xMI�1bt,W�s�G���K�F<u��	�Y:�2@��&5p��Ncks�YTԀD@M]��(��D:;&���%���Ά�O#��s���=k����`�@�ƸXWs��� B8)�hEA��>&R���R�o���GJ�<W��}�э3 F�LݾO�Zq���f��/�9�l��B�L"	��sI�r\i3)����vK䳼��;�x���� ����P��`?��ի������.������$S�P0Y�������ʌ�߿"����,-�&a�)v���Y>�u^�!�,����{Wq��f)��CU�E2��C6��?ܽY��Y��5v��O{�&nt����Y}�˸%�w�����H�$,����iH���dTTٮ��&��"#n�����w��7�Z�^��ʩ*�T'��9{����Zs�1����Ѣ�N��v�]�4!pZ!�UX����"�p���N�s�{�����̋�̍QV^,Q�����d�`·�Z��Q8��Ղ��>�w���J�K�v/�`4�d.Պ�`4�!:����@5�����\���z�\���<�3�+�\�~��$����)�tE��n>g6��0�4��EIE6A��f������_R��2T����*|<Z�?@��v W\U��޴����&���5+3��`畂-Y2� �K��lA3*�x���>��L9�m	0��f��%h�;օ�J�zhyd6'����S?��	�Zx���"�����<s8H�]�F��� ��>1Cy�	�k���{�"�^� 8_T��k��c@���8��s���Рxd�ޠ�|fd�J���{��h�3R�%		�"�,�̆�+%�rq+�R�łl���"%��s ��M�Fn6OS���������U)u>�To����+k��d�G�]-k)���jh���X�O>�l���d_�y�h�l:rR���te��O���&�mEM���<Rت�T�5U���G�>�w�D�Y[�bW�Κ��,�1��<��̎g� ���s�Ĉ$b0J�Vir��h�v4q"q��ف��`�[1,	V8��9���Y��-�}T����"-�W��ǹ��������j7�+�\@pA*��s�tE��,��~�|�z"��l4t�?U�{���i>7�yhq8y�JY)����J#�u5�RBA���a�Q��S�� ��\[;���_Z[[{���?�g>�`�z��O>}��G��?TgcC�.L?�E�$�!H 㐁]lv�riE��~�'Ow=����S
;�wl���ʘw�����d���A_�����=�&&9�ﺪ�L-.-M]����զ����"��3!@���^��B4�����^����J�OCt����Lr�4�F!+3DM"����T�b_��D{�ӷ���%�j��:A3U%5o ^��f�A{��3"�=h"�Ύ?��ή�e	�>H��}��K��dd��������b���g�޶���������=߇6*�KɁ���Z�z�6���R�i<"J���x4��)2�1�3��s�}p�E����F&Xŵ&7�4L��, b*�Z�1ĺ�34�迻���8�ez]�[�~H 8Q� 2s2
C�Y>�{A�"B���Q�z��'��d Ͻ�k-�0�kX;��� u�6l��'�ݩ:�._�����h(OB����H���MF�*����q����b6�P�{�K�!c�)U��LФ"��W���6��pȒ.Y�t�ge��Y�5��j�ۡ+�[7nK�S���կ}Q�^O��`��iq˕-W]���j��]-gZ.N5_�b84y�۪�@U����,�h����]z�բ�{��N����x__�Χ:��4Z4�^�������    IDATEU�}�,)dH��4�R�X�%W�9�2}��r�	�I#�
���" ����s�%8��5�a�2�D�g^�$�|L8;s��Eg���U�(dl�8D�-Κ|n�<�.>CNl�����'�t��<���[o���fh��5�g>�y]�sw&*ӘZ�f�]����ؒ/�K�����q�S����e��_�l����=oY�̺s���\�t����������l�ξ�����{�ɶ�<�ޚ=X�NN�:�?��'����nG+�����>�G�7���E���J�����K�7Ԇ$U��?���@O��ѣ}��?La��Gv`�-t��^z�VW����J�D�Ұ�&P�PY�9�F_湑��T��������C8�}��E��a�����ȼ�*�O����_����P�����H�eQ�P���((�Ž����MYy�%���"�~�T?��O|���oR�8v���E@��@��g	��̞`�x�h8U�
��ۼ�Z��R�G�m��U�\���%uz=WhTk��Ȳv$�4�Wt��<�*���q&%�L�΋� �>	)O0��Eϋj�`��|�����v!�W(�"/�`EC$��	�G�l�l��m�g�g�y�%6���_�ו}k��iTD�o'��z`,#UO�9�w��	�a�\���������K5����DC�eg:>ڷ(�t6T�ϕ
����+C����X�7��i�uDnh���aR�l+%��V�Q���z���hͦQ)rJ�]m޺yS��������W_Q���Ӄ���64���o�j�t�S?�X�J�3-�c���ը�]�߸To����w��V;muZU����zE���O���vO�-���.��ZQ{}��c5�/9�8`�B�����,��x�[F�������&�8/b=gr_��I�6i�;��3��<a��u��<&����O����7�E�J��1���o��$3��_�hw�Y-�S
�	b�P��p�a��� �彙�5���F�n4Y^��(&Np��c� 8�a��N2��I(�v�C�d
�H69W���%+J!�����JO׮\�O^�����E���3�k��?;{��w?~�����vVT�7�������)4#�ʥ]����j׋��?�'�>��ma���1%g�뽖�7��|eݎ/����N��w���ܣ�sO� Z��%�]���M���-����#���&g��I-�0Fb�@}�v�p��`D�v��Q8'�+3V���l��:/J{�2W�<Q�p���P�'ߔ
[*4ֵ}z��|�FuŔ���C�p-��׭�KU;������&����?�0��U���ֆx��l���X���چ��b��&X�M#��b�g��ve��m�t��CB�u�kBBs,�`��w�`�(U����=��|_sФ�K5���9�Q9��bl!����0E`~7�A��&�%H�ʓ�6�a�ǙHr�L���1b8?�Gs��b&��%��BRU-�qd�^�|�� �q�����V)[�	F&�}fV!Op��V	IC�J
ؖ�?���`���_H���N�#�WKe��#-ȉ��^p�M�����A#�3������f�������+f�'�~�^��j��^�x����'��oڄ��_�����U�� ؎t��C���X�©��h<	�4�R��*�ڥ�7a�Sf��R�m222�Po�j�T��?�@��H3p��P��|~���k��J���ό��ԪʉB3\/��h��,{t��G%���*�+Z$���^0��Y�X�y�&$,$?��Y��?�܉	�>'L8�8���1ߞ����z�z�Lwق%�'`�#�l-!=�b$�.�D����Cߞ/*c'#��ˋ��B!��4*��B$>z��ޣm�+[��IY{��+��{�\�{�$l;����{�����O��ȿ��������w���=�� ��U-J5C�'�=}���y�a�Pҍ뗵ui]+=���������c3�	�k���������ZK�:Y��b���G��=��ޙN�&�M���h*[�Lp��`����#��y���5�,4M-'W(�q�`��š��X,�J�k�W�V�
��gߓ��r��$o,��H7��L��P��L����o}���7�����<���>=H�C�#���pH��$,��������w����8z%il��;f%�J���/�N�����
����C������Lm|p,��[�
o���T�~.�����j�m�PW�_����e!�H�/�b�J�@��3���]-.�a��� )4��/�� ����H� }���l�@ܗ*��ȿ�*��<�������	�=�¸��ڨ\ �E���f�����X�ӛk�5� �P�5�.s��M"�r�3Ѹ/A���>�0���C�E��`oǁw:�_Hx��d�,�u���j
򼎭���~���A�A�]=��}x	������VǑLp�cr~r�u���/_�ȯ�|Y�bѢ�Û6u2.�P�b�k��{:��T�ٱ
�s��&YZ��c}%UjS�����|�.k��V�^R�Y0��Tmi4o��������P����m�m����s&���X�L(;h�Q$L�R�I:�.ݫ}� =�,r�
̞�E>y~�?���<��8|��:�$Q@�)�1�8��	�&Aг�H��C��ݞ�J��f��jΊgDP�0��E/8��\�33�ԲL~��]��Q��l��i�xu�7=q���e 8ۀ�c�����4e�bn�S@�+H�b��D��(�_��W����?�g>�`K���O����#W�mf)�̖:=X{x�w�D�q��U˩Q�l�{�=ܶ6-?	vO��֬q�lU5�m����v�����1*;E�q83�k��5�Ƶu�t���X�ؒ���t~6v�M al(/.��L�	�$p� t�T�V��8��J�����A��u��ly�r�X�W����������V���������*s����3l`�jŌI��y�-[�=z�H?�}[�e�(�lT��b7s���R?><���-���t�F}�,���b����e��]�&T���! 9"B�#1(EE�G�ר�u��e��I$8 �9�����n���s�ъ�E���9ԚBR���u	����D!��0������k��*�k�|(���N k�Є>�I-��FV"8��C�j��>Z����\%�v�s�-���L��ST�B��Xr�q027	,�%c/Z�j��b���{N��볓�*e��ЕA�^P�=���{���|��J[�.m�����ϭ���Vj�4íe���f�M�_�c��(a��#!�s�E<Nw�W����ك��k^��q�nhr1>�Ï���}��'*�U*��E_<ty+��.mu�,��hO�YR��0�kľ��j�!I�U�m���}��ɱf�KZ����ݐ�$ha,�	;2��r-�9�l[N���U����b�x%�DA�<�`Ԃg#Y@�N�1j���&k,�R�L�cS�x2�p���j%���\
Ҝ�8�$�
��0�Y�C����k̜G�62������aW,��1{#�Bf~�~=��D"���s )q� �ks`䀯��h2sɣF&=7�\@�-�D϶��Uk ���7��T(\���?ǯ�5�����{�~��ɞ��C�0�i�\��?h<����荇��ϓ�[v>�R@���ˊ���벑��'g���C�<_˯�Z�3���>������T]���uݾyI���Y�(,=|�X��:;�Ĝ'ݑ>�Q��q2k��9ż$���4�D/�E���S H$���<7����yĀz*����s�|����胻�|�Qc�����FjW�Aϟ� Pq"K`�#'g�(�Z�����w�g�F��s;�D�b���p����PÂ�X%����YS���tV���mm��tʆ����!Z�u���G&Hۑ�b���tO=1?��a0��ZN�Y�G�$������E�����*�ϙ�����cw��_m�ŵ��#*ѓ�+�TQmi�	�m�G�9��&�*�+F`�J!8���>؜`���מ�:�HDz��,�9m�DvIs�������r�v��Ns�Ǆ�nQ���J-1	Xh�3W��
�ۅ�7:j7kf@O�#=|��P2Z�^���$���40%GQXAFϖ�V5q͜E&�E]�tE���^zq������`��e�fE��R���~�����m�P<�!�G��%�tc���a�To��1���ޚ���|k�U�jK��^џ��~�ӧ�4oj0����hu}�m�>�*%T<C���Z��^`V�#��ӳs�jUW�$)T��&�q.�ll�G�e�ӭ�E3d̓�o
�v�0���?�SW�����Bk��J����c؞�j����x��dd�� �FŞ��R�NVz�3M�X�FA|TJ:�|N.Ir�~o�w�e�ӓ$��� ���لǀ�Mt4b����	(σ���|w����fK���W�����J�3�9~}��v�����{𣧻�:�����<f4{� �1	
��:��
���דǏ5<����F�m_M\^X��sΟ�X�n8�k</h0��dyZt?��t��\��BW�����k����>'���<���{O��s�q�S�:��-�A����G2"8�(	�F<df��b��W�I��
�3M��c���f�JeR=�с�m.��/_������k��Rs��T�g*�cp�*��n�ᓧ��g"nv�HVzY�>����E��*;�F�G��\$̀+��o��5&�,���ݻ�ɔD��[�^Օ˷5.uڟ6��uχ�F��"�����Z�b�&�5=>�5�@٬&�d'f�K�%�8�0!�ѷu�^L=��ly''�~��L��B5�A"�2Y��/{���y����T����D#�0��h��+9�ġ2�n_���c��jk��>gט��c�5�<����څ�u��Ey�D��y�L����^�}�^T�h����;�T-/�������с��Sk�$~�0�������'U&�{�Ͻ�j��ƈ5[е���V,u�ֆ�6����#���4*�ڑ���сv���=��T8Q��9��|'m�Z��ha؀��\���׻j5�l�\jQ��M�����R���a$nm}�m�=b���։���� /���m8�x�?�Ē���g�^��ͨXN8y����%��U������'��,���N�h�䗝~���X�qfe"�]�R;�3��`��D\J�[�<[�u�J�ɳm��ud*�Xp1`�\�0�]�Z�UG,��G����n)�vr+������rz�K���}��tz��FS+�6���/��r����s��q��_�_��vw�����O�;�-���hLO ���z�,Z�w��A������"	����Ug�d��<��C��޵�9}.z[�����>"dFf�a:\Z��VO/ݹ����g/y������~���5A���aRYa1DO%���������)��Uт�fZ��tѓa�r(�o�f]B���ED&؎G��\�o���qx���,_Sm�GC������y�
��ս��Z�D5kW�b���d`>��ѩ�y��q�y,�yHֽ�D��ل�a��:^jjw7�l�i����\՝_����Nφ:=�j<e&5�w�a$Ţ��l����_�HD��QS��٨<sW����s�B_�z�Ez�)�&������d@Oa���x��.HF���J�Z+2�A���I��"�)_a)�d8>��FEQ8W�E+W�������l
�9���hR����q<�ٸ>��Q@ٞN�������L�l>�l���֦XCXt� 19�xt�f����͍��\]�t��ӧu|�jbc�B�/\�����rH�q����FI���c��C۰ݸ|]��P�ځ�^�j}���xW'�K:��4+TTo4t�����j|���鶤3Uk1S�#s`$_��T�3�d#b�:��uu�u�q�5��6���ww���~�j���������kk���ؚ����"A���R���5S`��N�Jvz9H�����n$ey�D���>s�)��ٛ�fB�A�Y]�S�Y�6������ܽr��3]v���	|��Iv*K
i܋��!�)	�O����yA�֛e
�)����ovb���nʜb9Ɩ���hAb�]U���9�@����}P�gH��BI�Rɕm���K�o��v��*����k���;�������ۇ0gj���L���27tq�^�<Va���+.4|�ڷ�li}c����q>!;>>:"I�c�b#�X��Y~y��6$$�Dnݼ��UFL���{�����]=y��L�������I��'_��5��F���`����͟+��wu�o�	�X�&	!�q���;����w�����B����u�-f�;<U���|<��J[kk���7�����Z2�p�t�u>��`�P��ַh���p|���Ԁ���.nK0hޱ	9\WT��2^W��VouS��^7�9���U��z�/6o��L.:Yn1����`��c�Q�020ߣ�P�/���l��h2�7+�uaiƲ��Q�ED���ڪ�I��5h�5�=���0Énq
�����T��4O�p?m�@�!	9W)3��|�沈�V�=��?[`J��v��{R�u�q���W�6^���u�m��<O-��n��e�k:G2�F�|����67V,�_.M���t��F�s'*lhf��}v����i���?c�H"�{����my��-t�����m����O�u2��P!����LO�}��ў�����6'9N4"�Wt�RG�&F���րg�be�jk�Z��R���>:�7���J�+-�v(kt:L�����M!�n	�Er�J�~l�D�`��Q�]�ZXu�	d���(�y��T	�'P��3#�����IƌL��!)��\k��=����'=�|�9OB/�I�����7�ϕ�mN�9k�x�{>��d��/T/�]�dc*eFي�l���;����k��@1�^/�����E߻��Ҫ�L�BI
tq��=x�K��,
ь�s��\�����[?z�mi2/��~���d8���{��y[[Qasz��p]���u�7��[]�:�4�%�����mvY*�/<m��`m2�Ǹ��҅ɷ6״��o)mo�꓏��`�X�1~�!������Բ؀+�Rn;�K�ٮ���ᨒht;�ؘ�L�Ҩ���z�Ԓ�gj7����_����ӟ�\��5��R_�&j�ZZi7�����3L��:><
�i��	a���>><�~�;�<l�&�`�P�R��>�ՍMǘ�
�)�T.m�պ�jeM�:P���/��Vbd3,�TU��	��L�"C�`����C�3�Pr
X3��м��JR5g��?E��d�K.s�u�O6�V�U5Ϗ���υ�H�.�O"^���#�ST��9P�g�+Aw1Oͧ��MCw62��l&���r��WH���!��z֢�T��w .�pD`ϐ��`�×����G#�J�_�H6�-��B?�N��v�h�e�  ��b���P�GO�t��f��ץ� ���	��IJ�A����d�`;��
L��jθ�w�s��M��u�&&E�Jg�u��]l���~���i��=�TP�Lc��<aߎ����U��j�^�+�a��v���JI��Ted#K}�ɱ���O�,nj��jQm�h��N�٧���J�qIḺ2��H�i� E�v���s�l��X�<�ǹʼP�J�s�9<��%�����	3��L�+���s��`e��k6qZ�m] G�fe6﮴o��R�ͣ8�����,xJb>��pȌz�2��P݂��V�|�IV����*/K���������^�/ɴ��	���h%W� ��F�*��ѽv�ї��E�m�������l���������ޑp�[ݸ�r��Ó��������ƺ�V;�s����ybG���am�[���ىHV����p���G ��&���'}���
��    IDATd��x*�
��<}�v�i���S�c'�6�@�� %XgH%W����}�Yd��ć*'m/��w0|�!� rx���|�_,�U������_Q��~򓟫P�������D��\�暯�۬��ұ��4�f�>>w�����#O��g{�>�!a��@��l��C�-��"2w��h�n�Q��z풦��*զ^|�ݸ}E��P�(��a^HP�ҳ��a'��L�ǝ%�Ph����EUi�W~��Ȭs�6x�� 	4mVwѰ�E�M:�9�xB��Î+��`h��x���:���g-o71D$��I�\]$�����I�U�:sb�̱�/'�v1�~�ǁ��(�D+�9C�U*a�`H�ڤ0�{Z��Z�8����`�S�(���ԂlV?IYY�FYW�����4;~1g<�DG�Ou�lWW{j��=� >@���s���73��PN�o�f�cL�Zt�B��X-�ҭ4��V?�+/]1\Xm^ҬI�&E��^��o���g���F�#�zс6��2n���ZK��[jT�����n���+��]"�/6��G'�ỏ4_�4+64�5�1��j0�����}E2/n֤l"ibW+!CIki<]���cy/��\Y���ps�h^BRN�U�aפ�����Is�oK��=��S��d<�!`sO��t��fd	fz�Ȱ*��D��@��޿���C����\h��y=4����8��}��(��$Qc��'�}�F)�{o@�5G�t�?�"dD���XW�� �Nr����~�W^��?���}����O���ޓ}�G5{�*W[:8�kg������X+����cD�����;:>�`��,�`֝�^&���2[�a��uvr� ��hxG�m]V�hպ���.����,����
tba�̒��������7B�Þ�� ���B?���l^��p(�BJ1h	�z���׾��َ~����P��Ხ�!����$)8\з������q��ݷ�!w��P<����H���7=�}�8@���"����;aE�F�G�q!?��Z��Z��p�̊�x�K�zc]�ѱNώL��"�*����d���� ��D�;Q��x������%,�Ҩ �6T�<_�WK�l��h�{xv0��{�)�0$���`>��3�{u��o���ȣ41���:Y��S���e��ah`x�9,�*�"+������N��i�	�p����oJ���T�:s�E��$&�H~�-](���T ��I?�h�����ǩ_ 1��Pם��ToP�=*3��i-0r��xL[ׯ^��3�{��bv�67�{��s��з�%�n���m���'z����P��^S{�.�������?����X�>����|EUAj��p����z=ie�ι�L�o�K�7�V��4��.�z���6Ng]�0��N݁�d>�E�����$+��V�v����Ҏ�'��\��,��d^b�4ɍ�f�lr�Jթ�sZ[�2�b?a�f2���L�_F�SK��#)����EAr�+<�A�	�|�P��q�_�Z�!i	��v3��!�h�T��_�� ���vm@��DOַ%`�5a��X8<�d�#!�x�� �l+!�wS����߻s����.�no����>{��G��యj{E*�ut6��щ7��J(B�W�e�%�Xĺ�O�qQ�2O�!��(�v��2E<U��}`KL�B���9���a!�BT�b�#�<#�`�N���N�*P�c�j��:E�����;�9�<-n�K;~��_!x~��(�,�����ٮ��+�z�x����7���;��H���k�9>���4���@Z�����A�Rh�����	��p�-)T�rO&��l��*�$��k��0v_,�a��Z�T��kp0��^z���4��?��ҋM'9Q��tv��h�c\"�L�
1�j��p�u�4�ϩ��0n��,�(Ȝ��x���� ء�$�*�,��l�
H-sx>FG
i�'Xd�A4��ωT�q-
�d;9t�[.Ԭ2�u�`k��FqPf7��d�h�}a��aȿ�$n�H(聣%��^6��>��jN�Nfo�+��'����u���-#D4�
�nl�O�lTu��5�jGd�^��������~��4��h����%�~\�+vNe&f�ް��wT�!!0�u��3����l�O����Z��]]��+�U�,a�2?���?}W�������5_T,�A������U)B�*��k�K;`��n+��
v��m��R�j<��?~��h�P���e��!�P�nf5d?>똙l;%�,��pש����'�������m�N���,�m�>�.����5�Is����!c\������x����3yŴ�f�f̓`v�cj���V��FCB`R닿�}�xV�à!�-�'���h],�C�O���V+�|���T�	� �S�: 9���|'1�y�E�։
6��aʄ@M�y��Q���woܸ������~��O��}�3�;{*ԚR����3���&q���-�)c���o��uB��Y�Z��b�ˇs�`���f�s�Ⱦ�&NO�U*׵���j���Au2)6�e쐻ö���j���Ւ���K3�`;Z�y8 [��E�Ep"�V`N��8�=8�M�/������f�aQQ3��8>R�6�o��kZ����7��j�����x�i����pb_^���J�(�Z2o�.��:�������-l�L���6HR�IU�	@?��t�;��6U.�i�l�\�B^��Н�����p��gY
�;��'TWx�f�� �P��C&,��;�)�.#0�zGٍ�{�Y��X��gL�Yo�`Wp�d�Q��kZP�d!��A�
�RF�¨jb����p�Y���=F#�N�TŁAK��u��Ledy����C���?��e?wNK���pO�G��$���'�l$%=�^�`r�O��­h���M�`A�(Iǂ�i���--u�ʦ��l��Ug�h��=�'���Ό�������6*�����=�*�0W��F�R�VO��Wze���:خ�zj�.��������tU)ڳ�ho_������}�y�MC��yz|�Y,�}i���#7k͔-�H�m6���^ok4m��?���H�U�]���Wg�-L�
@H"P��y�
��.�IaZL�3#s9r JU0ךIL9�fd$vs�ڡ���ל�9�4�>?��s%i�;`�K>{�5�ϑD<��fw��ɉ�ǅ�$���/��`S�x8�-"y�,�^븀�����Y���:R�U��k�͝��D�wplH3�z�m.���P(�[��U�W=��v�B�lL .�͐���	EF�њ]��zk}}�������_~��'�!����)UJc������/&�3�4��?8��ٱe�2y�,;�[~�i��=9>teB5������~uK���`�rp�Z��ɥ��?�p�����7�x��vux��>�+�x�!�ѨX���&3;��
�4c�@�ٶ�~�-y-����)�镊nݺ�9E�w�`P��?P���_��_Qqz�?���R���j+W�ɓ�BK��XUg�R��PB���T���J�#6p,��Oe������tɒ0�Q�2�PM�j�(��P�Tn{̊M�uyS7o^���pt�6G����]o^����c����8�3��Ts��6g��|�$�o�g��|���!�i&q��/q@��J���$��P���s�Θ/��\�һb�(�n{x���XKC�A�\��`�+�ܻvp�(T��8��Ę"زv�~�3�`��V�3�����r=f��� ���Y@��@�V}T$�:RaNL��xu���@�9B4�:9�C�6ħs�Ҽ��&_Q�f)���9����	Yn<I"�ǌ�-��/���l	�o�~Ǫ?��Z_Ҭ�����I6uN���������\��:p�j5���:3�K�n���Z��Y��J��ҍ��I��bC��C�Ov�*�V�n&#C���*��%���"c��Σ?$�La[�("#B�Bv�s����=62a���j�!,	�D4��.ƽb�܉U��٫;%�[dlML2��Ř�}��n2�u��2��ѻgLdO�m��m�m���Oςmm�񑸛Ę�ˉꕅV;5m������vu�c����ٯ{4/�PF�gc�r�^����X�`k-�FӺ��D/��MT����k/��;����_��Y^����o����?��ގ��E���Um�=��~�Ȕ�4����?qi<�Go'���є��B�cX���z����~��fz��u��U�n�`�¢��^��{'�����v�\�n���S�������&CD5j�Wc��F;U�����{0 ~Gg}�y��@�&�� �"�0A����3o�˗/;�f����ݘ��˚������:+���~S�>���`�f��6~����g$���#�L�-������9U�w��]��N|�㪏({�{̘UlA�R��b������������+�|y�..�� 9�P��z���� ;Q)�=��F&��o�H�`��c�4�Xy���ΑXA����r�5Q�d�!	a�ڪ����A�[��4#��b����^�ٿ��,��d��g�"6���r��6[)f�X�٪�	J��<l���9�Yau����9���䮠��,�����t~����^�Qz����To�u��Zu�����qo<8���JŅU���W��o^��#QN�3��ؓ'g��*6��I#FLi������2�>����N�Ӛz[oi\hk��8:�$fӉ���?�g�~�b��s��N��J���f[kkܓ���.b-��\�n]���������~r���ʭ�(�L��}�Ao5�E�xF=�g�;��s(j[��9N'H��X7&-�p�Y��-J�r&.��X�6�-�R��3K~���(5`����wb�o"F�r��F�8y��y����~�\�:HO-��y��}�g���bb�r��VY��rK׶V��b@z��j����?;��|��yAG}�[C�jW*�\��l/	���0/�*�� �S��QG���-�v���n߼�_�Yb�/�=�k�}�d��~��ӯ�hW�ǧ�3#�+F��
lׁ���P�~�}M<�7vkb�4���e"��Z�'�p�"����ƕ����W,�#��JO�s��Kz�w����D��5����)嬛��d�.Dٽ��J]����r׺[�!=Y��.�&HjD9seQ�w�i]���+k�\�Z:�X+����o���َ����Z����=F(d�Ta��F��4�Xx�,6nf�N㐆�������w�����)5~>غ��P:>m�i�*VVT,3�ְ���k�zu�c\�J��3�?�ې�3|i�ڥ+W��ی�Z�����[��͌ݘ$1M�@~�1���`��`�j4��zV/UI;�Ƭ9���|��9�/VyQ�P�"���҆�[�����l�� U��T��F5�����q6�X�5���R:>�6���a� D�|y�u3� �]���( c`C��h0���ٱ��,�hiL���xaEY,.t�rO�N�������%�mOu����2�~T�T��gH�����c�4�sX�e@���&�b���k�O��d��z��U��tr&m]�UMK=� fcfCS���Cݽ�c͗��yň��rU���Ҕk�-���7W�47�&r��t�E�\]���X�r��{��]-Q9sЌѯ��~Q��!�@:��,�rJR�=�|Dp�T�ه
Y�O��Q��h�+<�|&��� H`^ǉ/`T�;$�9Pɴ�b0��;�/;�������S�ct2?3"�+ڋѽT�g4$����T�$|$��g;�q.�w���_yK��nh6>�Γ�n݄��23�e�����#���T��i�Nu[(h��rlQ�c����Y�G�m7�n�<��������{�H �����l?�����m�������R<�u:8�����)6��c�ր��	�C ;�p0ځ�hx�_��z�擾6Vz��/�ת�g[).]A�����^��p�w��=zzz�,��
Yp��0/�t{F��P	���/,�n��k�/i3���T����!�0B<�a�G�,���x*CX��@i }o�_�+o�8;�O~��f�--kk�>>բP��J'����zjDnշ��(fU�:=>�����la#{󑸧�(G����Z�N�#��Rq]�2��b�nH�_�k׮�Ǵ�EU�W�<F��N.?|>l?%fv1��w�ѓ�07cW��8��m��b̢�`�A����T�ANlߗ�%\-�'g֘ǳ̆�ʰʸ�{<Ahمk �8�.��%�,�'):����Vz����r����X�J �`�w�{S�s����	��#V]4Qd��UQT�Yc���gچ���a� �p� �S����f�g�X���"L���V�]6�rv��F�1v�Œ�����[��l�W*[~%��>�&��G@�=��� +��K#Bۯ�����O�{�~�W���h�K�S�_҃'6j �l��#��'����C���JTTT�ބ��By�zc�v��f?ՅZuf;Q��YEˎU�u�|�O��{2V���y 2�\�+9���$�Ct�S	su�(�I�)�,�Ņa�s��rd]"��`��W��0��E�Б��I�����L��8�4�@ӄ16�'a2��e������M*�A��X�!q��Xo�}90r 6a5��hK��3����@H22n�R�Z5��/���W7T\N�����vT,T����k�oke}Ò�}vO{�g*׺���T�45�0����&�rH���f\*�:���z�6����ҭ��?K��E����{{o�p���\�9{t~��;�z���ó���Q�z�é�7�QcbB?�H@���q��3i��>�]��z��֗���d�l�Q��#g���X[W��P���?zO�=��d��V�=$T�X(g�����}M��Ƞ�U�RV�m��[�ɏ 3�pZ�9&db&G�`�3��Dt8��~���]�R�/����'O���O5_^r�}�wh��j{�=�R7�MlPf��O���{��d�lh����s�칂L+%�p�9H�a�(\,�ZH(6U�D�-����*Ǳ��KRx.��>J�o��%6c� �%���`h��P����ru��9{b>�3z~C��Њ=�-CН
'�9���
����U���t��C�]���y�綷w.�u�&��tJE�>�<��[��\���|0e8=�������ID�gr9'�I� ��S�y��� ->z��֤�&��>�S!����$1V��o��S�S��iՐ8횉ܪ/U+�u~~������W�\2�L�1�QO0e�?��e$������F��l�$���嗾�5W����P_y�:�������%k��٣}�H:� �������'{j:9U���R�J3z����u�Qu;X�a ���v��h+������'�;.i��iY��?V��u~�$~�� ��L�}-�SA�(�2�	u�z��`Eu��>/��sf&���%=���ae8%����@&)ԙ��@s��Z/�{陂�n����pw�y�P��$3�1��5�S�)�{q.g^M&|���s���t�S�D��B/�pC[k-u�������6�]m]�jE�k76����Olk4.����i;A9Z_]Q6~��[�j�z�=]n�Zoe�iw��+[[������\�����+?z�O�O^|�dG��>u�v��@���3B)�����G��E��a��ɢ����4��(�0e��&gz����=�Z���՞�[�����ֶ������O��G4���lYf~:X�ӑ�zx�ӳ�4��<7�(�����0�_�����`6���3�ċ�1���N*Q����EݻwO~���S�x��/�zM������?Ѳt]��5=����`���%U�U-�1������o�*�e3����N��e�}�����W�d�g�`E�X �!��S���ru��(	�����7�jkk�ڳبq=�	>v��2k�~��j��ȖN�
6�����Q�$s;�CT�����D�m�/�_    IDAT)NK�_�`y�S�g��D�c��-�	_�~X��fӃ�TI��z��Bp���=��	�bD���d��#a2��i1���M�dF�~i��H���D�YoW2��r��Q�0���8=�X��쾓M�1�szt����,ˍ�ބP�"��ɝ#���w�Jy�Q�н�juf7��b��E�e]�믿n� ���<g:]�ּ_��Y1X��4�+z���o��Vc��O~�/�rI����w�jv��R��>�����V�]����ѓ���ϬjU+�T]Ԫ�M>ϰv,jm���u��j��-�9��M��u}�G��?�hQjjV����(]͆��L�?G�+�Z��U��Z���R&@�g��*_B1-�;��1;=�L	��G��^��s���f�s��T��f�<!)N R�6��ٴ�חU��(d8؞�	�r�O�g��?{�i���D���������+pdK�j��f���n=�KT����P���N���^�T�Z��G�=8W�
g�n��J�:�j0�G�A��8�2�UW�QR�����n�o������_���l���ƽ���ѽ'��~���t��ϴv���^ߦ�3w��]���LJA�/.�O��FZ��6Wѳ#���"���T��mݼ��Ŭ�ʈ 6r6zF��5�R-�spa�D��SF-(���4����P��WԮ8���&����d�ui�����o�r��XP���A���Z�pнu�'���'�v���߸���꽟}��|K��[���51Y�e8o>sU�����^z�:Ҩp� E������Z.k�9�>x���➒ 9S�T�����b��r��[�b��&���D�z���5��WR���E��Y��\!`����e������r��-����U"?g���=���oz�O{�d��*?�a��:x Ӧ@约f=A�������V�|f	��^H� g��U"� ��>}�R��c2��瑐he��W&6�γ���8����d(=JǞJ�$�;�	,Ge�����SL�#�E�6�C�cW2�
�����f�cMGG*��j� baW���FK/���ʵ��$>���ۦ���v:;g��R�\j,��ٹ�ܺ��^Y�G���ׯ�=<���������'�$�� ~��Y�����~�}}��FT���g;�	��^]�^Y�f\3c��f�5;m���U}�ǟj0nh`lM�FS��T��]�F����v�� ,xJ���3gbg�Hu�	G�g^�9J��E��ύ�2�v���b=%���re�4���g)W<W�#=��D�o$�Y&ДǯԪ��>c�W��v&b+�V���0'���e�d􆳓�!(�So o+�
���@>��ֶ��k��JQ��tS��CsmŶ��"��s���%�j��Am9��6�4j�������{�k����'��>�������?��ɹ�+����c�
wd�����������6�u�����LY���^�/)��Z�mH���d��p����g�6L���%���uX�ѧ��X&"N/�g�@�yoN�b��'�^�ge�c��k�4>��� f���®�h���F���\ԛ5w����zI_y�g����~�j��J�MF�Mjŀ;rq��E��o�=H~tr�
(�C��HC�W}���ٺ�M�X6X�B����f����e3���s�b�*|`��;
Ÿ99%oǠ~hU;0Y� �p?2���$`9s��C� �!��]	"��3)R��	j��0	XF������ox�1�
^�g ���`$A9;>��2�v�dtb���`���	#A������O"�T��4��J�I;��y���.k:�.��NV3����fT'��4�he�F=�=��̽���3s�<�c�|8�`�h1=W�)u�%���tr�n^2Ɉ1;��Vt�6�`���n811`>�	�@sH��a���s]����^E��w��_z�,��:�o�T��ݏ?��u�^{��豷����������Ç>�V��R�奺+L�\-ը�-ratաƊ��>���OO5�b(RW��ִXհT�����yI������j�P�Z��#�-����������cm�B�HUb�Hi��ƺ6g!�Ӌ��w���<��q�ԯM����m6�P���3�BN�B}�����BJo摌Є�<����LF�N�h��6F"�eNB��Y���s<Z<8j屸���p����h�,�vc[mVum���l������?��MkM+m���ԫV�R(���H%.T��j�7�q������_�`���w�[?����w���ǟj���=�%�I5L���l9��� r����dFV5"��q�,ؾ��ؠ��ek(��z��<Rc�-�Z�=A2.�l���o���꭮
��A]�����l�a�u�yz���,PK�R1A9�����Bzo*2|�����pg���kβ�9 v�o�?��jA���W5��o_��*7ֵ}x���Т��U9D��,�Y��ny�~8�j��@�څ0��%l� ���{�ϋ���\vM��ֶܳ��E2 
��jO��aR�R��\S&��3J�f�GJ\-�i:�2b�}����r
k"�fmV6g�L 's�<p2l"'^����B�B
B��)�s���Yq��\�lG1Ve�fmGs���O~��F@�Y"؁��dy�\��E�6&��H<L~1���|�<�D��z��jUQ�J���a.�Q�J�$�$��;0�kJ�0�p ,�!�a�ld\�>���~}u��u3?0t{�JO+�������^�����sp�N��_>W��`���3���C�>�ǭ���i.������[wti��'O�Ui��RmK�=|h.�k/�ѯ���t��5W�������7OG{Mдog���Іh�j6�KBΘjkU瓢>�lO;�@��g���|�F�V67u���߿���Jg��<�}��W0y�1�:A�1��_�o&��\�:��i�P�OeW��,^H��M(�	a������I^Hj�5�%��5-����3̜�Y;�%��&g��5qb���kO�:+Xe7�����&
&�4JDی}�|��0Y��8K�0���b2�a�f���zS�7���kw�� ��۟jT��k��˕JE됣�e5�UUͱ�t�]��ֵk��l>�Kl��e���������?�T{��8�U��9؃8��҂j#t���F�H�qH�[CH�E������;��,�S`��GσyZ6=g��ں�nm�ǐʊJ�pxx�jr��HG��L5�x~�P��Poc���6KF�t���E��bR�s�ų�Ţ+�F��K�[���l��p�>.�Vx�{ݶ3^FF�˅\s�z�L����H���;j��ѽ�����Ț+��M�����-t\�aTe�J�/�J'Ñ��9���I���K�i�=�R6rO*��c��rlTw4p��|�%�M(�#=sH����P���d�y�$�(6w�D����qh�^��[����b�U~}Ɗ��B󱀒����3G�@��+`d����ZU�Q��9x<T����@�|]���̑��<UFfC�5��ه0��{��C4 �<S@,�q��:ۜ�e-l��s��b�t��mg,���g��;݁t�؜�9�<S�{��V�����Hv�5C�;;O-�ꫯz�D��&��~#�-���9�]'��M�R�j�U��+�ըNl�~뎃���@���j����z��W�9��������;����O�C� Z�V��L�U1��E0S���O���������ǻ:��U���?��WR���~��v�����`���n��ӎ�*�J'=�>.�@C+�� �5/!��ݟM�vџ!�"��N^�zp-x3�ٸ� g��3�8�b����6�#�:`-g「bY2D/��� l�$!!��@n3����Yk��#M78�sO�/]v���s�� �r�����\@m* �͕]Z�h�Y�W�|G/�xK����'Rsê_L���jZ�p���y�EԼs�k�����/����@��.0������������w���`�3��J�L�s�@h̭!3��9S�"�ȼƪթ�g�׮;c��ӏ��艡�+�/��iyޕ,�﮴]]z<��憾����O�l�0t�����q��#=|�H��{���;:8>q�1!D!J5��� �{��<=>�X��5݆	'O�QX�\�E��J����g����l���f�����q豠W[,�Uց���������}[��j�����c������n����q٠GX�<�Z�"f�y�	O����Gi{{;���Atb�s�C�ֺV�*W�UA�Xb���k7���K!�?��6���B��g m#��#��o*[*��Fr�B�X�ͦ`'���{�
=fGC��I��dT�>{�;�8EbOb�� ����	��/�D������x�1k��d�ʨ��Y߬Z\u�S-��촨�3ٶd�	X������G��k[������z�&�ʶ��z���`Kekq.��,R����x�8 �� d�{'Gjf#���G&*K-ɃN���[)��g�:ؾ��[4������D�7G�E2]n��׃������	�_{�
R���\_{���]^���B����VupxlR�+/�v�mTj&Yq����w�{���*,Fբ�����q?�jR�B��W�ù��'���юΆ����k��"��$���݋��m6Z~n�=����l ��K$M��A�K�o3Iv��>	�ϋG���a���D�2�T'Y����5���_ӮY	���:�O&4��Ԛ �®ϣq&h��������V��8=�j�F����s��qKː
;��9�\Y�~��U)͵������m������Zi�h��R�8�k/l�o�n���?֬�S���5��hh�^S�f]��UMSp����ݾv���Kl?��������~����}������\�J�C�E��y�@�����;��`G���)'á{f�k��-Uk�y�n^�n�/����+q ����?;�Q��Ʀ0���ik�X�d:�x޺��Gz�t[�~���:<8ָ�N��vwAx|D��z�D��l��e���	D�2�ѿjhmu52��B��3�G�;x �c���a��i@�����~���P�4�7����/��vK��wt|6���rٛ!�ׁ�!@r�ФZΛ� �f�����jgg�BJ�:�Ϥ�zq��Z*�*��Z �wUĘ�V����=�D�s�`T�vxˆ�]"����3�4�3�Q�3P�Y�A��Rٮ� ���$A�
?��^e�/�H^�5��VR�+[�E�D��pr�5�Um�3��ƨ��f잳�1"��)[�nX+6�y\#��et�\�᭟�ѬP �nH6�'�Ϗ"�/�3�!��l0�U����lT;|?A��J���9F�U�ɲ��1t���f�s�[$ACU+��C��s#2~x�����v�roo�{��h��!h�f�	�����6[�MGч�w4�����+o��WzM�Z_�`���ٹ�ĩl��o��I����b������?��@��T��-�-4����+�N�c]P��0G�X�����>�τDA�Ɔad�����*ԁ%A���ϜZ���,.l)�n6��Q�I/��g��('������%�o��v�7�ap6�b�,�;�?����a��g�nY�-� @�$Z)A�4�-�8z;�b��� ,�g�N'i^<��^�F��F����e@�f4���NQw�l��*�?���NH�q����Ӯ�Z��fY���7�������_q���k���nj���*-@8;i�x���_޼v�?�Kl���{��~�~����U��a��)d�bE�VK�"Vp���4�l[�=aJ ��dp���o��7�_ѝ�/hsk�� =>�G��yX�?�&.�%��^χ��0���B�Nc��-�]�p:���u����G(L���޶G �@�@�;��17@��?Oʇi��X�#fUɾVV����L��r23úU�F.�င�!
0��)�+G���|]ݖ��o~GK�ȫ7���T�C�*5�`˜*=[f9$�{L0����wo#Yzf���qc�#������v�d�#q�y,2d`��'�oҋ˰�7�!z�G�˚��1lk �c�Zg��M��ޫ�k�̬�3#3�}1���?+���9l`�$ͮ%3"���}�;�X�Sܹs�=�L��]�$iO��J!�ɶDH�Ϫ�Fc��_�x�B�IN���E$�qY�Z"���B�,��_�tk�iq`�9�h2�p�Y���qV�xjx})ӕX<yX���M�F�4ǃ����/gL|�%	���$��b�co@S�a��S�������0����?�>���Vb���E�|e��;���>3ٲ؊��x,�2����[58"�Y�=��sŖ��'���8��R	a����v�D5
���v��x�|Ld#"/b����ݯ~�~��r�hȏ{���SuO����<�Kg�8bnq��W/������]|�sX],`<1	���'��v�E��|��_GLF@w��w��G���oc�k"��9�8�k&�PV2�>��%��sgq<�:��N�~� �`�TA*[Ĕ� �-��P�b�L�S�'By��P6C��l���|�%s���^܎i.������S^-�G#�W7f2�?>�҆�����{�\2�eb���C�}�����Lg���
�Ki�3͚��<c�����l�\�ȫS���[��"zt��51W���0W�λo���=I�"�9������ �^�u��+��8���H�6���<�J>�j>�
�*�����"(&�ouy���R���N�n��ﯯ?���;�����sT�aw��8�n1L0�B�H0C�XQ�K��4�{���*���2i,���ƍx��,-.�桉X&|�f��ԝ7''W~ѷջ�xƭy�
h�)�~k�5�����?:��~w>����H)�KK�
���F��B�?,˃˞;y3��2�7.a�j��݊�f�3�'��h�h�රpn1�R�>����bh~ﵷP?������y���f��L?�/��/�M[���z#���C��{����O?=ỗo��m 8YF�Fh_Gmm� �X���w�
����w���ǘؑL�?&��z�g� �B���AF�u�.���@QN�f�A$��l�%֩���D�1W��b�����Xt��7(U��r�&���{hJ�/�GjmccdsI5�I�!���%�Tl�$BYԟ��l_,�:�a���z^;Q�Ѯ=����V!�
�0�"B���y�\.�w��!L�N���o[OֳI�>;�r�}�;�d�f�
u�2�0��&a=Y�R�nGH$��@Cyr�76�輾u�>k6��jY߃�%5zZ	�v����=��$O�����s�b�i�Q��[��B�a�^B�F�ݑ5��kW��[�����iZ�>�z�������`�)R16Q���6�L*Pr|�M0�g��O���E��,F��$F��<܉�Qm�>�a��y?X��k(=��_����h��,��y�P���^�����S�l`���
��	���a��4K2f&�{�<�Yt���Ş��3�-k����՗� ��ĂkB�=��pr5��)���>�G�_9ƽ']�V�&�(��؈V-%͚t��恗_8/?��u�{���?~��@��\��� 7/f���\�Bi��m�X�*�m&�@�+J�Jγ^{�t�o-ͯ���T�v��k������jʵ�>��� ����x3���2�����Vl2�D�0�^״��8�U��+_�������FR�&f0�M�,�$	��[����?�]#���wǛ��闣�FS�Վp��=���{��㏤�]�pA�g�����6�ݾ�Ah� v�Ab�ȑ�HB>M+8�s��Φ���D�h�8�Ssz8��cC r��o.cn>�����fq���Q��?��*'��?F�N#��,���,��{2���8��Xk��)���8mBv@�    IDATu�6mA��H<%w/��sΉ����A��SV(����x�Lg��!l; ����#��}?;�[|��n��+�-��i�R*N�&["+�Ŗ:S[����ܺrxP�������u�adL�(3"���5Zm�[�S[��пXf�?*aɅ
ж�̮N�'RªZ;�IGәM�l4�8�PM��B�����ܳ��C<�rNEm�~�����qm����v�JD�)��K�=4٠�s"�Ln�f}�iKK�&$ލ���%�Lz#e�Q�0/���V\&�1C�:����R9@D$�X�75�����u\�:��sU��S̢0�d����0��7��կ}�T
�v�Q��~�w�	v7�I𳥬e$�G>C���LXlU0{��G?�/�0���s�F#B�YMH�=������9��5щLd�C?�陚8-8�a:�9c~�P�su����}��D.�'WԽ5'�;'� #@ܿf)Ex*�lv��P!wM?{~jhũp�"G|]��55��S�d���>����S�G�gn���ͤvl�jC��C�У�M3��P�:f����:x��"���x�=����M����q��^}y��t�X{{ml�0��g2��Ȗ��X�_A.g��Q�$��������)�ۏ߹��sﻭ���hH�>��g��f�Ǣ�Q���� �n���Q�t�,�-�Y���.C"/ޥ���ƭ[x���HD#�t1�ߋ��͞nNv�d�����[�2�\���O��~�2�4d{�E��<��vw���o���W�F�P�?�Q�.Vs���^��Q����05*�|B�q��E�n��R.�ɖw��v���H�	���&^|~�|�>��ý(*�G��`��a�%��p6��h�@�2>>d|H�r&�M����Mv��͹�i�as����x�(bT,^V��EB5LssUI>h��]3��=�$֧|�Zei��:h���y�ӿ�I	���'.eqR��lMc;x/�P�:�EE�[dl�2t���l�<��O�$�K� 0u�	��:Vg2Ǩ�D��A�\՟ow;*�6���`�CG��yy�tF�t������w������6qr�=�����P;����?�I�������%l���gc [���OM�d����a�g�ƙP�ZX� ��=�Ѥ�l*@u>�A���Ο�j��b�@�D7�WVљ@���a����uj&)G4�I8:埝��뗐����;�ꭋ�x����.f�KMs8j�%3�z�"^y�e�/�w�OPo���~��C��L'��Y�QƙI{.O�S�-�?���;Op�	D��Y�f$��n� 5���?�rm�]9��)Q�Q�P
^o�Ü]���W��k�XZ���EW�k~��5��w`$��q�4�?�>1�?4���޼��Ĺ{Q�5"$#{&8����YS`@�8"��-/�r�^|�\˙��[6��o�l|Ϛ��&lO)�#$R�X���#i�HL�vpi%�o}����:ַ�����V�|+���*^���+k+")�oֱ�?Fw�D�XUhL>�B9�j6�9fy�:ǳ��߮�V��/M��������7f�b����E$A�]�����8i�qx��6��X
D�j���_����q��M\�x%&aP���y�*�ԠZO������P9cz�ҳ���S�'��^�2�$�3���#|��m|��׵��W�Hfs�����Im"		��#dBm��,.�;SJ�A�-(<K3���0�9$XHX"H�(I�ǭ�/�X���'��R�%���5�H%�Q���#W��v�t���Y�|(Xl�0j��	R"xy8�O���8����>�� �!&�ON�Q�A΅<���k��/�U����y�j/)	D`��@���^:BgG���HJ����eW��'�)R�$�[XCC�Kf��~4� �fS6�y��q�N)>̂��4=�CB��$��{�3'�����C�ny��S��։���ÔN;$�PZD����/B"�H�k�6�A�n7�M=���ߏ�&��وSF�0M��?�����΄�Yl��fQ!��e͇ľV<&�hp�0�wn.����K/.��`�!ݠ��fҸv�P�|�<�)���DFo���?������d4�g�kz���-�ȗ�W��E��>�Ѵ�ͽ=��+��+�����G�?��qm���5:���bQ>t#يm2��'�m,]����O��ُ����,�=�pLCc�[A�f��/*��gv�܅�b�D�gb|�_Eۡig'[��G��d&�m�f@�~p��﫥	�"a�"~��3��ޓ<|��&&j\E"t����"W�z�5�l�h�-K":�F���5�41�/�ۭ`��6kQ�[L;@�|
��	rHRg;��K�|1��j�Dz���#<���D�
�(�.� �c}����!:��BE��t"*{�y ���e=��b���˿�KQl��_~���7NN�̅���!�AA���)���$1�0|<�f{�N/��$���6z�8����0_|��z�E\8wE
�u���yF����&���O�g>VM�Z��2A���ff��r�k2��/�@����z�G�������6�_�,���4����D�DOI<p�W���lJ�|dVw�-��h�d`�\A.�2֣X�}�&���W/"M�����үu��-2�c���4��l:Ԍ�{a��n7Cr�=b6��w2����
��~N$&�9]���_`N�	����}Vl9ٲ�r/|��E���X����E�9F��mZ�r���!��ʩ�חȆ�)�gd����MG��&���u���f��s�Ҋ�D�M��\����U<Lx����ke��vO2���P�rҝJ�����s(0����$HO�C��a�����e���(�zI6XN�-�+7�Z�3��~'�nͱ����b�u�&R�Fc!Ҕ�@�A#�g������Cy=��MS5�a
*W{�¾��p�g��X�½޾L-�\YƓ�w,@`2B>��s��Ԏ�&z�0pN����f����χ�݉�2����o\��d8���q��V��B�Xl��"�k5��������Ulo�Z�:vw�����R��&'H����� F�N�un�aWۓ���D��3��(�1y%�ОE��k�q��ۛ�Mn�#!�<���:p�t��W5��H��ܝ�F�TC�/���s C:i�-�55F��uM�qc��{) ��	X��KR��rj�_�o&xVX�M'6+�|>�<��1��3�2_l��Rs�J�ؚkZ��D��	zT�j��F��)L;d� W�W��1?���"�Ӯ�!�\uZuĢS��U��<xr�͝Fщ�HR$b�,�+��.WLZ(~�\^�O~)��ƃ�����{���E�!b<�E���]�+CM(�h�8;f�x�7��`�x��2�]���n����RI��Y�l�)R��#O�:�}��/��)��z��Zl5��p�3�D?��g�.�tfND��~|�^�-l(
����۷���$ߡ?gtf�� #N]�@{N2��'H�����.V�	C�����l�x��W�q��O6vTl��Z���ӳ��N=�����[���u����9R�D_d�#�T'U��#�T>�u�yD�,�8�T2���
�s
! 	³3���d8�A�wx��LtVj{t���hW�?�����	�ʁ�5Vv3Ā��@S.;·<D���Q�O{t��u1(L���~�~Wqvl��h1�.e���ɿtp�h��@���)�8���-ͦ�!�4<	��'��BD�=�}$��P:ȑϚ�X��ۤ#���{��,/���AƱ��Qy
�t�)��~'O��X02�W����8�$ad5 � "���<A�G����x������l���%5і��nT|�-ڒ���hH�y7��Sݛ,��P;������&�����#W��F�#T�6}/=��B��}�1���n>��{��oՐ��%��*%�O�#��S	2�$HKp��;�iK`dUl'���>7}ήaeQ$t�{���ͬY�xh�B؜�_�L�Cs��H��N���f��X�D��"˜d!ک��YX��N#��qOD��WH�I���
��3��O�QBVT����<v0��~E�r�6>C~�&	�_d�kW��I��e�����f��i�#>Ic��!�R-`::D!,�%�JG0W-I�����Rl��y��Q<zr���1b�,���և�Q�l�\K�
�,����KK��D���K��RM-��GW?��������xl���Xg��$\���D�T>R�G�9�&�|��?�ƥ+_�Wo}7o<��jEnH�By6�zF��3�i?������'��9�q~_龡A͟����������������vK� ���Ǔ�mtt�}��G'1�fPv�h"KFN,��A�t�def�rS��n�b�F�=��)�������ۋ �Y�7r��Ef��L�'>�>�h	�
�%���Qߢ����AJ�������t�L '�u|�S�Uxiޞ����� z3Pjc�G#��H���z}�jYly��y�NSIt4�q�Pf��q;=v�� ��Y\G𠑀|�5)����v���B87�2�C��J��$^�φЦJk�X��~(E��Lg���Ղ$�Y���=�H�d��rK%��H�li�����z,G��9��ݱ�h�����`�����d�u�6��<8%��qgn���hC���&!CΖ���ؒ]�YVlS�������1r� �R��-��^x�">��>���R��?��t�|~��!~^JRv�uM}�xD�ݛ���|�����X\Lbq��1D��P�\A�Ւ=�/�[�������ױ�~��E<�Gt�A">A4�f$�L:�b��3�'�b�H�_�ࣻ�h(�K������y������׉�'[z��m?������a�n^�F��q�Z���p;\Y���~u>�>��:��Va�%�U5o�h���c8Tq��6}����5� c��+'w>��(��z�z�K����u���?�3SN�����gw���~_�s�߳O��`rZl�4�/�}�r)�r1���^n˭���<���Y�����O�٦�BG$�L6�\)'�C�=D	d�E�Y,�Q���j�r�+���ΗXg��2��'��w��w��s
��r�H4`q�����W�]ìC���mC��+��e���+(�K��"j����t��&[s�_����3���)�-�g���t�������s���;��8�`���~��&�c���V�B$^0#�H=�� �Ha�P@1�,&YP"�騅^g��+/�ZM���?A��F����f��6�,���ȵ��=tk��6�;a�ّ�6��07�	C*����h����^?uNs)Dc����<ɜ�k�ŕE�9��mk^\S���m��d7�If�`�P��$���6�Y�9��e�o2+��"(ա�D��ܑ�2;�Tb���13�Vd�
Χ���a��� ZN����I�� ����ͺ��,M;RhS���]&��M��C��<�e�%��"�-�����dИ�f�r5�����̦�wB����<q��f����԰�ز������9�1RR��к�n�g��2D��!R��Mۨ�8=MQ;^G�⅛k��ѻh5��d{��%[�N�6��|��"ｃ#[��0�ɂ&���T^[;�0N/�-�χXẒٚ`8;���54�}�>��5��0�q|���'�bg{�L��H'�H��'�I�8��1">�l3E�����-��1��	 ��pb00Ȋ�?x�iM��{w���&��\�?�5QZ�J��u��'ľ��B�د5��up,�����N)SKXSF�"w��``���*�����WX���O���"�<���hg�&n���AG��\ۘ�����Y���/�g�'!U:�Ҙ���)��D/)�T��	Ʀ�ܔ
�\�s<�	�F���uM ���^7�3��,.T�0���Ҩ34�{�;.̗17_� 3Y�.|=�)��e��/����^|�蓷N�7�"�
r�]�=�����b��W��tJ���Q��H���__y�K�:lH"�����e�p���v�E���U�C�u��/?�:2nw�)�X�\��>�٢�91�`8�ko����>:�����-B+Sۡqҥ�n�T,�h{��3�[XB�P՞�_��a��Z��R���6��9���h�٣F�8��6z�˜M�)�=l�`>�0�@r�`����Cko��������-Y�����hg0���b�*���
*�¤��)4M�ڿ�qi86�)u�� v��f@���MQ�ͻز�-�͓S�`z=��d�hS� /�7Y�⾘Ŗ�$I�.�C#�p�H�dM�
*�Y����L�^�����L�h��m̝��R$�p�JR(9B)t�`q�#��C�v��v�qJ%�95;H��*OlG�& g��sN�(����Zy��}ĝ;=��p'\�AJ�4���#�5�p<2F>$��K�D�.�O6��6��WV���o���HE��Sf1�`n�������[�_��6j'�1����R������cmy1�BN�4��U���o�ީ [����&��I�nWV�t�-<}� �V���HG�6��N�-�'�d�t��>>���f/���q�َ�1��B�C�50�V�L��k�T�u��B�`"Nf��E������.$#dl����Y�؈�i�DPc���p�d>0�=�Y6�DC"����;���Q+�3�]�2�p��L���:4���I��pCn���|vB��.��83l�`0��X���7�T�Y��8��}���{��7�/���;�KƑ�E��������&"2�A,�v��Vӂ9ίTq���v��6�L�)5�<�h��P�bya�,����R7�<�K�l�w��/���b��h�5�!u�3��C��-�����.E�%�����7��W^�����F#qX�;�$�s��Y.�����[Grr��[�״��s��t���䅬m�ܪ���p��C<y��Ǜ��m�� ;���'��0Y�r�T�|e'�:u��\�T0��${�a�Ά�t.^�����!�e*�sܴ�of���أ#�d>@�l��h(�R.�$#�Y���	�{��}���'a~�F�R��%�a�'�"�XV�ș|�J	��z�(g \l�B6U��S�g�2�!�KY�q��8q8�c�1F�,ʧLa�Or�����96��$d�l>֭CIP�l�$��tH0iJ�Ȭ|SK�b���!a�)^7Ncb"3/3m�Al�q��q�����%$�HJ���~��F�DQ�fL,������H��a}?!��瞝�9s۲�zF����f����H�2�M�3M��+N""I�O3�*ϋ0S~616�	��VW���h�����q��
�~�5l�?F1���v����dV0C��D�^�A�m���^7Y��dK�`�D�ay)�R!T�Q��xf���Z�dA��4���q�����S5��k_�m<W�w��L��ҙ�K�pp������Ic0K��-��ͤ�O���t���\,	��3�A`͌��3ř�J>lpEpJ�����x���]��2y}�I�W��1��/�R,��������C�k6�>�Y�Ξ�E[�m7}�V��L93� rE6�SY1�)��״�PN�{���x���5��&�M"N|/�o�|��$�����%���m)���'����9|[��M�d-�t��Wqum��>Z'5L�1������P�Q�!���\e	�KK�W�ߎD�I��Ҿ��b;����^{�����N�ݦ���>�������@�<0��tZ]��\�_��~�/^r�Y�s��<��E>%��{A����U�N�j;3�^}w�w%[�!_雹�p<���>^{�ث�vr�Π�V��v�Q���zKH�?A�PE6W�d��&��R���|�A�N�e��n����n�����:��Ջ�O��9�a%�q�D�[opBO�tR�<p��9�}�
�e� &y��S���Ӝ]!}�%��Eo�"b�
�D�t�=�ܛX��:�����^�K{    IDATHL�!/�����GDZRj�H��9��,�m�"홙F�28���Թ˟�DWl�i:��A_ƪ4M.u�lH3��:b���ힰ铇r:e!�L�������t�=s&�r�>SVz���w��"C3�pӏ��'�|��X���e�'b�M�Z	��;[<1��L�U�]�`��v{��5M�V��ۼ�ݾ1�e�Hϩ�p�^����!�h0F29E�Ȣ�&'�ry�|Z0��.M.�*�4��u�S�p����y&�Q����0���k3��T�8����`<8�{X;_���v;GiT����IEFr
�''ZO����u'�S$cD@�(�Rʯ�Ԯ2��{GJ�bH���o�G�9N)�g#��@�d�S�2C�xh�OC~���c�"t�Ƞ��/c�4�ϖ�y�5�'���̈=�N���U��5���&2$��!d����8O��n�}��0���2BikF�Ԫ( ߠo��l��.n�d��B�-�K��o�ݴ-X�&!����7�H�K �(�A��D�K#� �9��ΐ�A�+�X���X��r�l̕3�/e��s�06����
�YX:/���0"w�L*�s媸0+K����}��Ԑ/�g��b[ۺ�����k�u�����C�b�Ѩ���{������5���x��W��o}[�I��l�V�}y����E�>_l�Vp�������
"qNR?�g�!D���?z�ܿ�V��I�P^�{�t
O7w����1����|^0���!R�$��U\��"�0e!�u�������%���`�K#]XFw�A��H2�n5��
s��)?��<�_%�s	�X4(?Kv�5n<zl�w���i����(�2K�ED��/ ˜�=b��8��6���R���1؝�5������]>ITc�u�1�i`oNH��C5��u�
fW.����jcʞ���!f&!\�<F����O!]A�q��H�J�L �t���&OB��s����zYh�E�\���"fw�Y�g	%&���=��=Y�i��MX}�?�l�l�o�-^�i591�~�9Hy���)MHZ!���E�g�6���d>��A�X\J!�w���P.��j8<�C��p��VW�����0R*l]���dE�YG�}b��}#�̢$��u���e�&���)n\[B1b������9l��sH���v��N���	B�C2S����Ɛ��E�bC.�G"ERY�X&�����`�nA���,�����\�h���ؒ%��͌`c����c1�	_;ƻ/���� �KY��g�@g��:�$�2+K��Ŗ��;Q?m�%rş����"lF9��H;��.�Qz}.
�[i�o�~?^/#�{P�����f���+�>J����E�1�5���b@[���>�(Ⓢ4�����������'Rp7�j5��(�(f�q�*�����kwp��e��"v�"�B�T�J1����ŕ�_����/ZG�ȟ�R���o�������u�v���u���#4�S�jV�+a~�"�(!���w���e��_�<w��C>���+6k�_D��w;K����|�P��9�f?�	�yꌶW/�`���>�w^�.�����ci�ӷ���B���>��O�=F{0Eo,��!�/���H�{˥2n�?�`�C@Ӂi��>�^]ƍ+�x�Ul��9tF1�Z�t��g����d+�|p9�r�᎘�"�'��B_�w�c��(v��:�%Y��Ԡ2f�jk��bU��Z�O�/^�t��a>0�wJ"!F^�b0�p�� ��c^u��|M5b����۔'�:jr]��T����n��Gh�]>��ͭ�lgMl:t���6TR��be�L�hE��N~F�Ÿs�-N�k����S�=&�}�6�kW숀�3���J+�6	��b{k+����v��D;�8�V��K3�E�����dK��>�����8M�N+@������rF�6��![�Q,dQoc4����.]^C����q���
�hQ�%��C����ў���k�g<ʵ�P��4�W���]|�7��;{-l�fW���+�v�Z�w������@ؐec2N#���-l<�"�!�<�d�P�����Үqc��b���Tџ �*4�a|�+����<��"$q�=;����m��n��=���1�g͔��.v�7��=O��!�����ʸ�VM��:gs�����[?-��C��Ho<Wup�1��j�s�y�$.��s3CC�t���<����ͅ����l+�z�b��g��0'w��^1�N���#2S8�	wǌf�O������ϑ薊!W�X[�ô����S,-�C����{N,�/a>��:�������/�g�Ŷ�9\���ۇG[壓<����Q�^���ܳ.V��+T��J&]��IG-���-|�֫��. ���N�,��ߤ	0>W�~�O�O����`�!���ԍ��>��ϊ�Ʈ=�"ǚ��������#|t�Ct�}EV���_�K�;:��_��3H�
��-�yR����9�|�*b�>�̪6����޼�����F��̼&[[rKy6j�&�l�`��K<�l"c�����UWp��=ܿ{�R��>�7��z8�k�E-�'ZF�,�a�|N�-�TB�!5�$?��czb���{��"�4��[q!c�?���:r������|Xw8i%��pph�Kyӭ���z܎����6�^���?�0�n�_�}�r�����0Ⱥ�b���<����it�=c�
zV����YD	��`�u��No)�g�i;Έd|3�(�	�����f�Ab�ɜؒ�d���~y8{����>��W��f�@TA��d�2S�Qʞh4������F2�������6.^<�ã}L�,/����K�Ŷ�-��~�8Q�Ȥ���׏��k�b���}-Ic��Q?�D"���^�!�������Q�����=��r�lO����&�SF�@R<��L�hK���l�L�[:��^;��b&����{?U��U�S��3`1�:�A��<ـqZR�s����mP
�g,j$'���Ӛ>+�~e��"�?���J��v�d�ۿ9٪K^g%NR�q�`zd"H�ٖ�IIƄ8n����%=0f���#7�E�7�wB�jn]�(�)�2��*�d�LqG��ٹ��YU>�!�Y`*�>B��Xl�1mz���'�t���陙�.i��<��c��'X](am��b:��ځ�m�����z��̞�X���-�������%���_x���6�ڇ�o�v7��w��qC��J���0W�J0�P*�%!U;�,`{��d��֯ai�R�����p�?����k���v�È��3]�4��j?�#�M[3�8�����+��G�M������������4���߻~�9������m"W�W%�	#2����I�ֵ+H$��?A���7�ṫ�x�ͷ1꧐�.�=��N?fK�!�dȈ�I�l�X<�J٢�"k<P����C<�{�l�|�&�K�!��w7��mP���6�B.�U��S#W*��RN��EA�C1�Y0mj�0wk�h���A"�p���r�Qg*����˦14�vx�J��z&��Ro��A��yd.�{i�u�*�����`06[ʖu�lm��ih�����3ja��gl>	��n���H4LW��W��,ac�Z	S���K���PD(�2xM��u�'�������lZDH�!�-H��ab'tA�d��u��D1�3#��GX�O ��y����M�"#,/�c{�)�X֖p��%t�m��m�U���a�"�f�~�`�w�g���T֎q\�|��u��|nY2�۟n`c;D�z�׷U ��%��lm�v��ᨥ(�x���!�L�I���Fiilmg�b�ͅ*�L����Z��A^�v���o0�~�O������M�H ���f�b���,;y�xL*f��/�g��02��?�Td�K):�v0�K�M ����G|ʃ(C�u'���9�>N�]o6aܟ���F��L�H��w�ȧ�[H�1���?ϒ�,�B秇�]���C0=���	��g��f4t���?b�q��� A�tI��'�'�XJ��|s�,�1���8>i�3aqa���_&�C�:���+������~����Ï���;����Si�(���͆�ᚯ����E�6fS��#J�2��o�����֭o�����ek�����������A�M}���7�ى��,?iYݷ�E����|Zl	�p5U v��;��ƽ����Qk����
fMgڕ�i�HQ}2�]	��q�`�/_D��<��'hu�p��y<mEŶ�K LΡ5�����\e�)�9a2��a�G	{���áb{�>������c��wc¼F	Lg)�2"r���u��
T+�x��mq�����Р�z\�� �Mh��e��3Ss��{�������_�a9�s��Μ��;~�Vӌ<R|>'� d�������vQ�}��!���PQR��k�)8~0��|�5�r�}Vgɽ'���S�t� �ײs�2(�l��ب(RbH��̘�~�a#�UBҭV[�V�n ��ܞ���&#�[-��Y�-���lĦu�V��l��H��x�t
���|�`�St��XX(JN���!ҙ�]_����N��B�$o�I̤{$�����~0$�7�H�V�1�[M��/��9@>���+�����v�r��W�ѧ����P*
윜ึ�	-�&y '�	�q�j
�����t�#Q��!r�"�$6wZ���]�zy�����f�9V�c,*>f��}�{�߯����d�k�w�n?��b���+�=�7�g��,ɏ1�y]M;m�u�c@Ձ���b�����	�M�k݋Ϊ���e�IR���{N�m�*a���ZxH���3�)3�ǥ�l�:�h'Rb�`�(��<�6�]Ģ3ՎB&���#�[-�霔�9��Z�aׁߓ��t<�r6�J9���B�$s���1]ʦb�/-��3�D^,��rq��ykʟ��~��v6�ſ���������֡겒�Lp�<m�z(d��"�L�tL�ݡ�;�o}�o`i�qo�o�և-�b;s�w?�;��V��g:Cq�a=���Fw7��@6՞��q��u����?��?��x���N}b���H��Nh�0�����`��Ƥ�µ�X,0m��k��j����x�<�����v9�Tl4��6�~g��o�Ⱦ��I�)�2X�X@5Er�8��n<Yǀӓb��m)���9�q"J��r�ep<�m�\B�)sy�T#�@��"-��bˊbݰI>X����>�*N"c|���~��*�JёSؙ� �n<����c�%�Չ��2�bks���d.��];��<X<T�Ʉ�e�ג�J���(�:FF�:M����4��[�!j�;��5R=��m�e��u&R�)�i*�4ݷg&v��������i-��B�'k��!k�Gt�2;A�K�Kٙ���T�!��F��٤����������B
��vdq��E\X#Ԍ���g@�Mj59ݴ����M��%I���k����F�p�ZYٹ��b�(�0s�߾�f��j���$�V��ųE�!2��� �}�'��Q�%�ϥeI�R."�H��扛l�D��0!��;r^�'��Ą��Mr��V���-G�
$���,7}A��+��=���D=�Y6|��,������h�;���4�?Wߘ�u��Xl��p�B5?á�	~�LD���|}|���H�;cUI���B��:��U�L�&@���숯�ރ���ǚn'���k�qnu	[O7������6l����T
� !�|&C6�J��R�%��e�:�ޖ��Y�U�ۦ���dro�.^��U4���9K�O�q��V�_������vwOd(O�Tj��ky\X�`��Ÿw�|J�w��$j�@,�ï��o�tfeqG��ǋ-����w��b�JR�}�կ�q�������L��ق{�3�c`%�D����/������`b�,�~�L^R�F��0�G�T��f���z]u��.����f�z�c�6p��^z~�|�	�}N�Y�'t�1�"N�,�d#��AOtj�V-3C��d#D��qj2�㇏����~��b��0=�U!�.�89�i$�0�F�\D�\@����M@�eJW�/��d;��n�����7v7H�����i�sd���roG��m�l2�(��p{��fl�������,�3i��e� �i��K�M?Y��bgs��1apN�c���s��?��9�N�l"E0S�f0��V���f��y��IC���_ȓ�;��s���;��ڵ*4 nF�|�<L����c#��u��������-�2�d�
�ϐhA�nN�F�'�N�r�47E�,��}������|�.]��"��8쎔��B��bE.B�?4�Z`��1�2lS23��ڥ+(��kky,-g�ֻw�d+D�tY�m��THx6�s�@���0N-/���b�Ꮰ�O(+;�RJ�T�"��I�\\)�ؽ�!��@�$�b_�v"�����bK�(N�BV\���5�I�0�#������/�~��I++_�<����)l�--
��`^���,�2>�V`���X��:��)kb홙�]�����˸Npϖ&K�C����Y��V,?{fHJ�}��
��+'l��!$i6���Ջ�y�V|x��6��@v�#��tb	DcIi�s��X��<W Ӕ�<��h��3�%��rN��d2u�X]����?g����v��q�����ѽ���<L���L�p��"�H<9F0�c�k���H�)�ތ"�?�[_��b%6�`�AR�����@�r��������ݝTu�.���z�nP��E�������s�S:㦛��������~�z�z���I,,��~�t]j�EDC������ʸ]*�p��*b�&�6�O6�����'ҺV��posǭ���8�pz�	wl$%3�z�y˺�d�v�����l�nlbs}�`dA�6��ɖ76#i��J.b!1$�l��l��yB02Fv�|�:]z�����%j�ulZF�
N:ER<�D��;s 9�9V��7����M!���X8֤4��4�'=N�"s�Α�w���q� ��ϒ��	A`"����"��Np��̇U�mͅ�E(Y��=ML�NS���*V�c�g�EU��C�5~��hpB�������f���b�W|��-�Shp�"y?�P�ul����0�G�<$�i����c��B���7'�I������� �/,���sΛ9�v�'��a}N���n���:�5ԋ�7�L�I2�W��"=��J�)���#<X҅˸}�t��*������`�h@����(f��|�뛠�Q.g�	ӈp痍"U(Kg��G�?
1B� 9�GZ2��(��z���`R��[��Dۭ;�L�����R���	ғ�<��� �<Ȥ%f:eޗ2����i,..�\�����!�=��������'�{��?۟B�\���D/��(�;6S��wk[~q��&�5���$�zO"ś޹�<F:P.�qnuQ�~~�p�{5ds}�a�#���~�$J�@&Lj�-eE!�r�U<�#H��J<KF���+�<㇗V׾��U>����O�[��b��w����|��b�R��Ͷn���4�*1���btx�(>��i�!��P�^�_�U�XiR:��v�z�����9߁/��>E��mY�I���y.E�[����]��g^���4Kl�)���G���}�=�p�k�{�Je������NF�#��Hg�hwprp��?�2��[A���1�-,/f�^��O>E-�\��G;5�Ȝpx �i�9���(�Ŋ��`�h����>��3�Alm>�'��십��)�g.�+����UǤne�-Q,�-���Ȯ�=�c��m�m(���#�C��Skj���������wa��4��/�>$@;�3"�^L�qLH��KسB	��0�0��/'Y�YԢ��
&���&�o1'V�"����MC��pz�9�;?;?]��Z�w.�Y�c���4��gw�u�nٔ��)�����3����$1nwl�9��R�    IDAT�@�c� I��u�� Ȣ�I�H�b����#2��
N#ar�J9�ag[����C��-��Ν_�Ҳ���&Byr��&[�'Gh4X��l��<�A�c����9�<�wP�XXL�O7�d'�X�n�H�w1��D�}|�᠍):c���a>F.E�"J�~���D4�f��LD�/$�-Wq��.~���,"a�X�H��@!q���Cݫ"�e�s��`42�<��~V�]�_x��!�?ˉϯR�}��{:�Ҹ@׏�)�%,�|l�y?����[Ζ�1��(�R:_���F�{�{Zck�~�n�D˝�����uϯ��eJ��'[~/"Dr�RN70t������@��v��TZ�w�>��>��sEE�r�2�İwX�����8�F4��+X\;�gR�ɴVHE�r�(�w?�b���������>���o������G�՘Y�S�)w1���b��)�<�G��ف�7v4�ci�&�]x 4@˿�tU��LFN�������?g�e����;?ә��&�?����� s�Q�}�֛x��7dj��{~��(�|��G���p�)z㩴���<�ɬ�ۻ�[(g�X��Q�M۠�fmKi|��U<�� �	��2�[h�0ۃ�����1��#S�w�$�	J6C|>���666��{�� �_4��n8Q��D�1����RΝ��\��u�3����I2�c������l���40�t89?سSV,~,.�F�NG�R��w	S{�(M��D�[M���Y�MǚV�����3�E�)C�$˽��4���~>?1OH�d��A-�,O���$FKg;�c3T�d>"��󛺿�]������n��_#�����4Ȟ��_d�+C~��g�Ό/2�^to�HsJ�KG�5����c����#�1�>���B.�L6Ĺ�e��W��ӹ�<���(��S�p���]�����7�,[�k9	19���y-��u,��P.x�d��y�b��p]�@Hm1��I�~�=���E�����H�@,6=�l�6`�m* �/`s����]G��G4Y�8��-�r��Ŗ������~����������[C�Xlcr�{�\���O�����[;ۘ5�,����Ѷ����@����,b����d���I�N�+'=�ŖϬ�~�#�7G`�{�hJ/�3����=AJ����y?�!�X>+�Sz �z�����5,��nw�l���L�A.P��T2�K��aq�����5||w�HR:��a�U�M%l��z�x,)��\6�b.�B��0����7��s��/|�}������`�o��٩�כ��I�3vE�^Y*��O"F0_-�\.��"�gq��(�W�N1���i1Ӛ���T�����(�v�?�����l'�g2��� ��ĩ}�G�$���7��y����RXM��|Il<����1�4���U�Q(Wu�qwʽm>��b!��b�~͓�U�x���x��&�4R����Nd`!Z�����a�Ύ-���N��v��?��;�a�Gعb�|J��)�Ñɀ��L-���]&��~6�	���R�
�gi�:�1	�B��^��!a�g��f�!v����Ӳ�A�E,p��ܠ9g����^.D�v��:��7�?2��|d��f���m�#��FoN�@vN��c����Ǆ�V>}�y��� tCy49+���~�k�/�I;l@��k��)���L$���.S�;��Ȯ���SB���ז�P:kɘ�bGk��S)�xx��'B�S��q/#WL�ҥ�[����;�0�G��E��X'��w͂r�Ҽ���}v#q\�x�F��^)"�ak��F�i�6��i�M,����79�!%�hf�6Jt��3�I,T
�ZDd� ���������d[F�Mk�����@��F9��e[���l��wk�Ŗ]���⡞E<���Yq�Uǳ�����H;F����CY���y�$dE��y*�lf���f���lG��C F��?�*�^��5ql�=Y�?Ӿq�����I����$q2&T ad�t��˫Y|����������z8<a��x����� �ڷ޻�1�He�jb�y01�ŖLzj�i�A|,��z���b6�b�)h	,�-�͕�����������ޠ��N�fWn:��Vk�䄶m�VR�ٕU+$�ƳR]�7^�KHg*��%�ԉ|�ت�����YkO��}�gE��$�g�R_��?S���	��~����x��7�t$�j��Lżn�N�QSc	OQ\�/�2����C<y�P1ys�<��eT���ho�T��k/]R��l�E���Z{�bKkHA�D���ȲX�t�� s9=$���ݎ(�~�ܹsO=R��Y���u �h<���H��0�Hc���X���veuA���F���T0ha"��� $���ir	o���!�Y����\v0� �.Ϧ3�#w)��VPy�y���󡧦�f<�����{���>�1&��ŕ��4K'��ə:�F�'�1IR�C6����ͳ%}��Zvؚ:	����b�����,΀+�N�X�Z����n5���� ��MQ����Yl-���61���+x��H��HHl������T�I��؜jYlYH���b�M�^]���!.4��F&�T���Ӹ|e�+��灞
�cj�>��ټ������W��O��kR�0í_�C���{x��ET*Q4�{�Es���޾
w��Ĩ���7����$�G<$HhR��"Ld	ȝm.G��35�QG�	~��}4�9 ^�~J6<�D�V'C>��ͫ���qєj*d�Ｋc��Z�����|V�<�c��5Y�����('��o�=K[��׷2~O�zC!RV<�yWl�$>c*�ͨ�3n� ��~w�z�;~�sN���;�H�˵%�I��N�>� ��yB�C ���Y��v���2^�u��Sý�:�jtG	}�|&�VJ��+�Q*��p}����b�լ�}�� J�(rY�1��5�3*d\_�<��4����Z[\��_������9�������pt��d���{��q���ఉz�#!��ɸL%����X^^����C,T�S��c�S��3��+nuQ�P^?�}���Vw6��~��I����ӿ�^�X�F3�΃����{���1j�mK�ʜZ= aR�w�r�*ҙ���w������v�tkK��e�k�P�m!����c��sȗ��D��m��&[���R��39d��r��>����ّ7����L G#�ۦ�a'�HR:�db�h�Xa2�\!��Ŋ�jgFL���p��d���1߻��Xl���ӏ�>*����}-)�V4찲��)9�M�����)E8bh<su��5�_O.�$�bK����b*��A�ݶX��8NZ]��8�o�d���nU���Hd�8k
�=O-X��Q�G���w�����hſ�v+�g��L)RĠ�aψ.|���?jJ-8��B�&��;V?�S��c�������(�O[�f�j�:���B�d��X����{趎���+++�2X][���׌��`�H\��F�Dg�I��P��M�4��Ԫ�L����1�5������ʸq���z����wC���0��w��A���= 6B�Tl��RQ¨Vl���L�bFSN�*��v������s�9�ĕ�D���b�(�Ԗ���=��;[��W�\��4�ld��~j�g�������y�T�"�d`��-B�k9^G�Raj5�Xc*�~�������ʘ�vh�u76�w݃�׽Ζ�)5®��Q����)_�^�+��Dv_|&�16=��5��p�C6�ƫ_Y����"ll��O��w2�4V ´��˙��7.������x������|i#w�//,��ϡɌ�Ns�yD�9���/�N�Ҳb��ϩ�/�OWΝ��~������/���~��{��?xe2nJ@_S>��� �'=eCt�;1�����7�7q��Y��S���4n;A=S�(~�k��O����	N&��������w��>�jl>v��]l5��v�?y�u�����8i�Б�(��F◈Bt{��d
e�>p?>��#�� 5��a<h㨶�B>�n��9<觐+.�3���LojN\,��^tC'��d�H�3�+u �iu;*
��''X__��b��-�Nc�Ftg�^J�$��<�ʵ-�X��T* _H#�5�pD�8���T�¨}���A;s�n�S�o��C|:�JI�i�L�u���ƂM)�WT����0����;XA���2iKy�z]�#��-��Vt|M#i�iy�h�{��VR1��r���t�[VN�hŖi'�0qw�v\cs�g�)]�m�G�'6.���l�qFv4�RNVl��&�l6��g�҄A���)��_�I�BvV���,'/:G"���9��N12=o��G�xG;Ѫ��r��-��J����������f�����N���#L���o����)��wo�&��_��q�{��by)�W���^w��Fh��=!"�t�ð�A�ݔ	���m(��L�"�L�)����4��l#�%g��G���x�N�$�@+��Dޔ"�H�d���?km��V�����4��u!�����Rg���P�'��?�x/s��$��;ڤ+ܞ����Xl��	�a��۩�ݎ�ʑ���Y��E�r0�4��ϟOg)��R"(��imYl=�2�ri�!��s�҄��G':��c��������+K�z�F�<z����}��V�h	��0��QH�s\9��B|rw=E"M����^�y+K��������Ve]�lv�NeQ��S�f1�dٕ�17ws3�=����ܷ����b�I6���$P�P҇����@��>�SЯ�}�CF�8ͨ�ӭ�=;�2�r��3c��}7_�s���&��"�ʁDfFF�[�����{�����Z����ų��ӯI���mq�+���o���_~ލ��}H��>Àr0C�;C�6@�C����|l�#�%�����~�wTӐ]�{j���˫2,�{��d��`�wQ�������f���$%��D-��i2��7�8j������W�&3礏�M��a*�t&P�������V�Xs��l��;�:��{��ӸzeO=F��B����,�F�'� B>d� EbI$T���[ُ�Ȍ����c{{[��>�z��n9��L�4���b#�'�A-��_���;m�D�����Ǡ�J�X�bܘ��Sq�::�\��1uB81�m��g�Y�����)2%���(Ş���9�fj
o2B!g��<xI�R��IѨ��Xe����D	����r.<�f�>IM1ݬhg:����sy�;�Ȅ���P?�c#~�C/�c�2g�y(J�6N��Y�&~�6�/R�o�'*�݆��[�sK��Qp?m?���Y�$�?�7aGA�Nq��{�����CU�/"Q+��a:õUG6MY�'h���1e����XZ]���*Μ;�{���A��Z͚�<&/GG���`>�9pB�\�YJ���KW�{]|~�X���w�{ln����b︅�=~��AcsJB���%(�Y�|H�y�s)�m˅<���LĹ�<�)�}�Ǎ,�̜F�w�J�F
ZD�
��L��_�{��78��Qc�Jp%������B�81}r# �}Iu(%3i��C�$�Ǎ�G�֖���Fmh�'�&*wa���hl
P|ޯ�T�x2^��C���P��\���Z4�(pI,Mxv��=d!��ul%�4���7W��
�GΧ�85����4�C�Zu<yQÇ7�PD�sr^��Ҩ��b0��3+XZ;��z���9�ꕗ����KgN���3x����ӛ�dzS;��_���S�bI�������/������7��8��ƾ���?��Q��0>�#q�[�}��]2����ץ"�T8�x!�}��c,�l�����@�
�!�΃��,�	1%��}�kL���b=yO�]�B�L�o1�'�f�����	[���Kޏg*%'�A��_~�	���?�}V�����'ì��+_�˕�$��ϟ<E��=�t�W��X*�ש��<F>\����[���BT�khvf�&��2���(E"(V�D�	!��w7;�=�Vvst��� uttd�,dS��J�}S�a1��0�d�_D��cqy+�VD~�����4Ly<&ӡ��&�}�=�
�����Kf�Svb��N�N��M�Y�pg��Z��0�M#�Iژf:\�cr��p+�j5��7���Bd�$��\���b)��:�}�$�Lԏ7�GK�$�AG�/�E��3�/T,`�-�!j���),a�e�t$3�V=����$Pp5��a޻lU�T������3���{��+�Z�@���3͠�#\c� x�D���6�i�u6�JW�R�S�Vqjc]ϹVob4 t��ς�Ҭ��3��3=V��b��c�<_���i���/���+Kx�����a�a��#��kf�=�i�Vu��8	�t�*�	�(�\D'�!
yZэ�˥�8_F����L*�C�5ç��5�a8�3��*'������Vq�[���$����x;�x=� �uƗ�ގ���$�[��}Ȝ@	�u&!|�	T�:�~&E�o��(�q2L�1�ڕ����{�0v0��:dB�R�WA2k��<'���D[t�$�e�M,����5�f$%���X� d����9�����{W��1'r�g����V�i	#/�v/F6㡐�QL��9����b����1<����YY���o���nyKF0��U,��i�|��a��(_T�e2]ɗ���KW��WP�-���w����>�<�/൑�cA%c��X��m�(K���g��t�I�����c���k�`m㼬���Nt��hċq�5��-�w܀H���4 ��)}my#��eMcgO��[���/�\�q;���V���37��̧��H�C:_,)h<{���#�'SD�/���bI3iq��(l�^��'[��o�q|<D�;����C��1P<D�@m�,����H�Y72$��9����
~9>>6-]�oɔ�D�I�+,H�ћ~�#�������{|�<�D�VLa�$(��F���T���>�^�|�*H��bIj�fKE���{��aEi�I�DB���d���1��lU�R"�a&dR�/{�|�i6�:�X�%c��8��j�lb�4�'61PD0J��<;�d�F��U���6�� -�oSql,H�U;��.�jT�%��eF`{��(ߣ;���D�LUjS��	���9K�����Uq3���L�,QK|�ɮ�~�XH��j�=y�׍14���>�Y~�D�	���V����t:�$��Q�!D�2���ٻ&$��	��T/Of�?��I�����p���yc	�N����{8����ϲO�1f0���Y�!�y,�B�ii!3�)�s4!�P-��F*
Kצ���4�F���͹�BL94�u���,2[���p��kh���rXK�ص���d4���HG����Bͮ����:X5k��#�{I
tg ���1�M����k�g2��%�},$���L2!���,�P{9�� ���B��s����QI�Ff��3��~�ͲZ�G�{],����w/`u�,��_}���Ec���`�4��i:����mbu}�>�����8�SKkx��&�^8�/n�����++X[�@!�x� Q�(62��R�ϯ�����`��Ώ��n���y��md�>�|���.+&�񈋋�a�,����$�^?�\~����b��!r���@2؝���t�7���Y?��4f�z��c��mquR�P�U��G�&z� e�k2 R����٧��Ge���H��/�>C��@H ���+X�T���h7�b�Z����d����+g�m���ѐ\X0�,u�3+�}'͞�GfYg�g�[BJ��Uf�a��6��b�+ ��!W����N��.%[V��|����T�:A� ,�$� i���]N��x��jc���R3�]M��os�X$�'��CK�5�F����nyOX�x�R�����.�Y��WSU,�o���u=S�%5z��$@�#�wK�׮t��X�p!����HV!d��F4aR�$D���Br&D�D��$�s��d"�ե#	    IDAT�2{���=1}wS�
�W�*g(�}+v��6{���"Y��΀���'`O�/7���-��tD�:>��\\^R"B�q
�æX��E��*{�L�Tq��	��}��\���ӧw���p�l^����.�=l`�1ad�uӧ�Ϥm�֟)�f��Ŋ��շ�(}�K�W)�$��7W�C����_m�э0�"L)�/$�W����=[�"���3.'����]��z����ƒ�t�[����LyC��H�3��SA�[P.���Ҏ�y�'��
��a�������<Z*�sZ���-5���Q��s��i�5�]B̽��
lm�=Z�{N_;��I�.�$�
�%���?��Y��V�#����n�Ⱅ��+�a���(�=D����:6�,�7�ν�x�h�6pisW.]�g7o�����"VVV����Z�)�El�,������������~���[�������F��������gP���R�2fʸY6�Md<Q�g��ӈ'9|��?A�z�ER�R_���*���6l��k���6!����%�753��h��n��|�_~�):��)ڃ���܈m����bd�$��('^����l�P�X�/c�T�O9�G&
��{�1��*�1����N��wDF"�&�X��G!�3�A�)1*��s`ܬ��n|���g�N>�%	}����O���|����d�t"���*�a�ʑRz�\�BA�����$JE#W��f6R��oi�f�����4l���f	m[_3I�l���~���y�
���~Tv�X��� {�6�:����[��8����n��l�T�2P$,nͩ������d�($)� �
��I� �I]�}�8��?ڲyh'��A��2ee�ǛlI#䘦T!5�CZ���@ո�;hy8��������4��`�)DϞ�ʺX_)������3U����������y�ӿ�ȗ��z�����6����g#�hx`��V5����o~��o�
��Z�v�vv��f�'��}�3�Ar̄r����ɗ�`;WM+�F��!�|�^\��z'DL�l���<�̛��fL�X1�2i�>�x�D,,iH��h$�dR�*IW_�Ɇ%>�7[��������8��$�2��|�g�BI+�Ml���b�2�cr���S�����)����_1��糿,���!'��u(���_A�B�DJlUa�@�o�*�h#�ʊR�|J����rz�������K�;|��[����C����ϋ<�V�l��r)�Ba��/�an�g_G�n|�X��o���g��ڍ;�;l��Z������768�G1_I�R(��W��Я�}�h��}��?j<�i6C�HRQ��N}��=�=9wi�J��JS�U��y�9,/_ťK?D6�(*e��ył',Ȳ?��4�u~hۈ��F�ӿQ�&��w
!��Hh�?�����|�����_�_���=l����L����M�#0�~-�F9�9��N�-�(o�E8����R��p��sl96��P<`�No$�3}s�4��*s(��(�"ɺ��Bכ��jP�Eu|y�KU�Χ]�6���&Ǚ��e&K���$ز�]Y[�
��L�\�Ԉ����L��VV����욌l�[�1��tlY1���p,�����)73�I�	l�J�Bf��50�P�G�7+�j"rBv2�����Lo���$�0��c/�
[��$%�@�w�>	�ڸ�~W� ǂ!���4Ǡ��C�Y�k�*�$�&о�[��2W����I~��I�Z�5�qV�fM��۩�CX�ql�g�d3P�~0ؒk���~����"ܠ��������>QV�@�SS�]ZYRCFr6��"C4�A,�@�����YO�yJht�Ź<�q��q��"^�D�m[���G��b{��8�!���M�8%�MR<ǪlǱ��J���$�(�sJR�T��g����l��l�L�&$A/�U�+���)cBcɴk�9g-A�J*����6��D�r=Q�K�?�E&b,ҿN1˗�M�F���3�Ȥ}���p�|i���}@���ɟ2��lL֟cJ3IY+�OdI���j�Of����~���65$���K�-���6�%LQL{(3���&�|m��>��K|��c��D�M�b&��g\93��+!V�SD�N,0�<x|��[���w���ͳ����t��(�x���c�|!���"��ʵ�\~�ݯO������^�s����=o�:�md�
%��Y6$�aL̟�WBsC�Ӯ6�l�C��� B���7�/}�)�N��sV{r=ݿ�O����M$y>؟L�8�7�?���/�
�fK���Vm���>�rv�4�eP�ϲ�Gqz��Q�5��c,��X[�<b'#�mc:驲;
���5��w���4��mƒ�*|T��.��̓��D���nJ�y�>��S��^��
h�aH�(v�a�NM��<��ױ��$&�@�Sh���u���rY�IV!�c3\g��>�#:�^/�*;#�F8E���c����dF�V�%yP'�6�z���8��\�N�<�͆U�|�2�7�|xisJa�����!)�����c���:z=���"LL�	�!*������1h�G�_����K�Âb@�(eD���*'#�$կ�$*e���V�����x�)ΐx�R�D�'R��8=E�yx���(�%�z�F�r�}�)���|���^�OQ���u�/T����{B�{�|a�>_$6w��M��R����q	���s��I[b.���|��l.ă�6~��g�x���VO�1ip}�:�Iq�*]��"���	P.汸8�6B�ٚ�k[h�B�@RTF�-�-�yL�y}�l%���a�Z|i��g�Sd7˪J�U|����a����Z���^��L���N�l�Q�������|�+�T	wT��j�#�q�ްJ�4�e�"�<|�DA.����D�xI�%�,$ʙ�'I���W��F^$��`+�`�Cf6C!�A�!^?���\=����l���㨕B6��p�^���Jo_Z�����@��8��G��c��z��E��o����x��B&����޸x�n5���ǒ�6@5_�����y�ϯ�=�P���lv+x|���ao��{�T��J��	7��C,�1����h8�h��O��v�o�G?�S�͛x9}	\�T�Z�F���@�I�=�w��﫯d��7*[����`Baq��G#��-|������֓'��N���ͣW�'�92G9������rs4�#�Q4`��B+�U�#2c��:���X^2��A��S�����.���t\_�Pi
s�T�7T���\!��"v�F����Mf�՜!V9Ζ���* �s���by^B˫:,Ɏ�j�ȓX>�����\"����dLR�9a����b�����"!�����,@�n������fr�`+x{6s�(�}��T�
&%)cΰ�)���^dp!���("1��p��iFk]��L�x�}r��U�b.�r�aa��9z�f3F�K�-+[GP���{>����4�?u���	�8"�!FwB���{yj��3�)}Ǡ�G���a�'��/Ip˰�)����1��X��q�5��(�S�����
��N]��D!����l�a@&p��M�Yي%���'�,T���CK9�鴣`K�Ϋ�Kȗ
�{�^{�Z�}����|��QW�d
WH�1E�����l_�z�2�F���S�T�`��q-�ǟ=F{@��P��l'3�P��Q�$�FN*[��~nB�J�m�X����/gmyݔC���o����@���;����
���#�X�+�a�}�ޭ,�ȶ�$�f�W���ZP;�������s�1��Y݉|�h����M9d�-,&.����*BB�bl��fv�(�"d1���Ο)��2��>�v��0^F<4r��jﾵ�S�i�:{�}��yLS<��&�:"�{O�sЁ�^B����s��w%�R��O��p���������|�7l��O���a�w��] �\�1F6��L�`Kb�0Na4��<����ZN���:��"��?�3��d\d�ʸu�:���`KT�y�"����1v�q����ǟ(ж�}I0�4^��N��̌�\(Z,(3��:�^lo+P�&;�SX.�X-�(��᠇V��9��[�!Ν��t���O^���g�m�(�i���`�cEL?�}��)�S��/�����_ȲL��rV�!MK:���u���C�ba�ʂ�����Zݎ�,6�Uvn���4��X�S�Ȳy>e�q�ͫ��͙XZoS�3W��0ac�[�<4�W���hA�D.�
�����}�{O�1z)��u0^+ߟ��`hOc!�jA�3�7�Ɯcv��Vm�
`�M�-k�6����2�aN��^���/Sz�b��.2-��X��-IH*"k�����[sSc���l�_��>f�K��!ǳhtNIK��cB���aƶI���vk�Y�M�8�:�7e#I�������=)ȉ`(���3W����Bs��6�Q)��k��{���~���������<���;9���Fq�:|�~qV�M���E1.�k�F(WR����Ffp�
&pX�q��t�U��᥻^lI�IDyH�bɂ���+��3#A�/�3)�͐"���xZ����є��6?W��F����*d���bdz��a�̔Jc�$*��P��m��=!i��
7!�%�2n��[טl����-���%r��mҳ=�ݾL0�}�i�����Y�ty��Z%��J［?���k����,�L�8�XM�O��*V�}4�^�Q�)��RB�E��)�b>zv�f�����)��?���y	�e��7W�C>,ܸx���_%x~���ƃ��ӏ��ݝ���h��\8D�Js�`�4�[SU]�a�a�Q��J�bo���,P����S�6@U��.`:�!boBN:����\�1Y�g��;$V%�Q�m�7!��zu�
β����3���Zw�ݑ$omm�_��?�ͻ��#)V�"�Ni���B,��7+�c«��GR�j�[xBҬ��P���+�Q.�(V�;��(�3�Sv�F>?���
��`(����0�]�x2�N�Y
�Ls�rCR�L;�w����� 0qe�h�g�ʖ��W�+���Eyc7� !M&[��E� ��k �[V��\e���T�a���oM&]I���ib��Y�p�k:�X2��*�2o��y ��H����[��\�U-��c}��^��ԩ)L�Z/@7�(x,;�/o��fS�������[��pSeIƖ���gm+�A��d�z�V�����"��ꖇ�#�)�-!k��^P=D}ƬXs�铙jltދ^��� r-�C��7{�:d�ɛ'���4ߧ6s)t�MY�f���T=�0b8F���Q�F�~A�2��X����+��,�#��+��l�`���X?�����,�V���;��޿�`Ds��%l�1��e��������IN+��FU)&'��-��s�;���!�,Ʃ������3��dePgB�_Iϖm����M1&IL��γ�������
b_�r�K��	w9��_#,�����>f���C	�{�2��s�׎E�
2Y�)Cʽ�f�i�*9�H���r.?TGS��\�FR�>��O�'������<�Lɫ�M��������&�i<bBG�TsQ�y&?���A��c��.~��h7"�K��.�g��Q��������G��V0�i^��+P-X�~��3�`e,�h~����4�9]�J���!�?=�y齯H�����v���j��;�@&�A�Qțl��;=2ڲ8<b�x���1=;�'\Һ�&T�Sx���O��Op��Yp���S�T�`#�Ghэ�$��d%�տ�k���ފ�[���M��7�NP~����ƒ�|]��޼��G�Qo��e2�i�̓�P>7M `����b�>88�����xM��H�l)
P�B�O�w]�l�R����zQT���y�۸}�.z���D[���.R���#E%/2��j7;��Ɔ��7�"$���$��d!��F�>rK�k��d�%<D��V�$8:�D�B�YO��
6a�`Ul��u��H�T��֯\:s0o�kgOH�eL���bX���R'�e��%i�YS���3�݁�!F#�[�M'��"+
BAH��)/�Ԝ�\3�gB��&��#��`c�W�0�Ӏ>{v���DHٌ���;��o�/{r�_�iUA���rQw��a�6���P~�'�Y��Ϟjb�&]^j���֤�gfGU�0�i�6� ��2MZ�l�!p��-E�(
5���ͱ��SnHDs��"
rd�k6�,��l�x8�7+0��<�"~��(UKx򬇟�����y�S�^��Y<T�6H�bb9F�3)�d�9���\4S�˪V��t$��k7���ssRj
�>��_�F1Q��_�FֺuĢ�*2a#'A�U����#VI6Ǒ���ǂ���5��Z^g�i��<�S3��3�<ësԏk��jb��̓?-fs4}�:��ku�P�:�A�6���u�֐�b�e��78\�_��eI�9��o������@g]z�C��1�P.���?8��װ��9~���0�����sc�����P,Lq����>�3��RuMc�K8{�,���G�x�׆-#ȗ��P�S8�?T넣�KK+dS_�x����J����������l�v_ 巐B�(�B1��$%v_�5���G���)��&�������Jκ��mQ������w�_z�<�H �Y��~��Y
L��k�IIX�&Vvq�J�������Add��D�d+��x���_���O+��f-�9x"%�&+5�d�b��C���~%j���q����}��I��=���ʹ �|�Lcn�A_}�j5��ag��i�je�~��M}d��Q7u4�8W))0��̌��&����g��&a��I�e ��f�1�z�c#s�'��rj]�6�YDH�ߏ�ΰL8�*4���)�7�3щ��tQq��Ó'���.<�d�2W��@c� E$�"�nտ���̟j�6��a�@�i�\SO��G�v��ӜAl,#�Ɂg�J�$h4�b��	�
��;�lZ��
h�
����4x��ph�%�+�㎽���AT���LT�R�b�a026+��4�����
��}MI�т�	X��Q�.5|��8�g�K�11k��Q$A�O
�{b��mds��a8E���Q�.�p�pG����&۞2��ۖY����.Y�=􇝓`��2�v�1B�x�im���*^�:'�������M�hF^�=���ynΣ��'�9��O&��Ϭ )�X,�4o[�$ G���|�\��9�2�9:�*�N5~B8�������B�t���Z�h��s�=M�术�dd��b��ugS���Z�JTˮ1{�Dh�6����1�j��O�\)�4|����f�@����O2߈��㠼��K�LȊcE�4�%"���|�	e�®3im�#��k5���J�7��⪐����^�)�R:�R4�w�^ś�\�Q������J�F.g8�9��_�����~��QoͰ�|Zm�j!�Q[f������҅e�p�/�p��i���س�`��n\ܼ�퀑[��Z;x���3`ڄ�6�Ԅ��Cg����n|�;{mt�����{�F��4��,��m�.�������&ݑH$3�m�5	����_a�%���9j�k������_\gӈD�l��f��:n���?��}���;�h2���m6�G�!�C=N:q$� I29�xb�a%H�&��b�z��XѓQ9Q�-DU��dZ\�'}T+�W�8د���*hu)���6�=2b"//.8r����+�@�mZV���u���a�6{G.���B�	g�<�T�Rqk���Ӂ�|��t(�5;�G�-��F���-P�Ҁ��}�0�m�Z�P�ʑF�`;�Y���9ִ/�K�I�p��u�y�Y�,�����v_3�w��k-�9���{y`6Nȩ��    IDAT�V��b5�˄��+�Ҟ������KQ�r���j��F}��B9��3�Mi6Z#�՜������-�c�DY��Pw�5.P�f�1�
�t":�S	���ȓ�p�*,�O������4��.�DBܜhfpfX�R�LH��6�� ���ɰ�vc��ֱt��8/�Z��Ң*�Z�.X�=Y*�)������
��n�F����(���v�]�o�λ���+��zT�_��3ԛ$EV�H��gB�a�� �L��&Vp��H�L�~�ʖ�o&'������),ͤaLT�a�r�]��|�h=K�̄�k�IKl��fy8⡑H�3���ͱ�3�Cc='�;SDK�8�*�c��#�8Km�FJ-!���/�����\�$��]bC;�����:�#�����901#��#�*n3P낤D�Yg��@��O�����F$jQ�|�E�J��I��p�l.�Biaw�?ŵO���#�͋�{�]���kh֎q��/�b����]�˦���3XZ�ãǇ��p 8@ǿ��
Rt;[�����hZACyyi���[gO]�v�z��?�?���|�I\Cj�3Ȑ=�I�������C��T�.���1Zݱ�����Y:�15���_��?���2[�t����E�B&�1���`�,���UT�C*y?��"�b�3�����|w�o�§ׯ��ľ	3v�e�����-�/J���$Fr"l+��:O&�k���C��1G"Bք�C��a�B��w1dY}v�T)t�C��7l�Fo�����:�-`mek+��`�6QGR/��-��$�ep�s �HN��A�^S�^�Y�����<���y�'
�R&�e��d�g�11	#�sX\X6��8�kg\%���U�)�� �Q$'Q��;�D�68BR���}��UP�\�*��g�̵dD���%�&�dc�6�`@Z���Lh�$
`�Z�{h܆A$0!	V�Pj6Q�P,�hy���D����
�d/��C�P|�|Č]�s�Vu��j���of�牨��Oށ1�=�9*�%�eF�R<Dy�jL�Vv�	3�%��:(	uj�}��Oa�6����QG<�aW��Sg6���"�N�ݖ�ǯ��kdr0�9��RO�/E��1����饅<�zs���i<y��O~�+�\�D��A�Ȁ3�3a�C�ƈ	I@�|8C��F�Ĺ��X�	�����.jmۜi�3�M�-���i�F]^^A�k#p#@��\w��xҶS���);�P�rs�d'�_�3Kz�I�dւ-��C�"2��"��4�`E��+�혼(Y�S���M pd�ۄ��^-_�a�O�v�E �MZ�d�x�Ѿ��0B��S���$�7�jҒg�e�lk�ǛE.�觐�NQ�ϰ�T��g���ɵ���;F��a�o㻯��ݷ/"㏱����6��3�Z���[WQ.U���n��AnnS���Jή�~@���b�`�x�����^F�o�O�8��>��9~~��x���K�����ut�t����r�g�l�ɳ=��{�;nc4��
ʺ	w�L0�`�R��3�U1�.-�w������8�pE��(�_�N�02f�A��$H�D��ĳ	z�Ϸ_���>�:ԓ�=�Ze�\���Ԇrs�I�0zL��_��E��h�U\>�w�쭐��kfo���h�B��\1B�*D���8�`�����i����UA	�u�(hAUE�w<sE��,-�H=Y/�HD"�C-[?�=����_��AѨ|�`����-��W�q�*gV;�J%�8�#d��q	�d<3[&k����ܜ�ѥR��q~YA��k�cs󞈵�~�/j���F���9�e�d%Q�J�NN,"C�pl�R�b�8�
����`�Z������)��/^c��K��U�#�GC���O��
� O�D���7��% q2������<��c��]�'��4,�� Tu��8�$��I�d��$d�)eL�Y>����X�ݞ#�X�e��V�pg0�b6�p�C�Do�6��C���aԫ#&qo�Srw��Y�//�գ��e�hL�a���*�U ����V�����m�Y?B!Jae����,�b�ϕpp<ƿ��k8�qv�ƚx��������1�,E-�\Y!U��
/�r��\y��1>��}��<����Y�FT�"�n$��e�����р�z�
&�T��`�?�JB`\P�s��K�7�k- "%/�b#;%4Ω�	M�EV��i=3O���7��d�ˢ`�u�yig�����Hp4���q�V��`˯1زZֹF�����'�'ҫ���̟ϓ~�\w1[e�|c�G4�"LM�X	�/ȕM�k���&u%_����4^�����5S���n���s�/�qjyQd����:@y�,F���8����aWk��w�6[�u���d�g0xz���c��z��d����{�[w��է�r�5,�Q�uĤ�>���g�q��.�n�1�He)��(r��KMf(�K�z�<���k��Z�.1k*��I��~���2K9�$�R}Y9��WAI6�϶_�Ͽį>�����4=d���N�#��	:�Q��m������[(�2��u�b���;g�M�
��0-V6�R�H	6"_��gZ��p�ƃ'�E��Vs��Q.V������~6�j=�XJ6V	�S�0�=|�;w�����wr���_qR�yT�
�"��y%�|퐕����PvO`;c�ud�r����ER����w��	r��$#��D�GF��:oc~:��	�K�f��3Y�%��NDT2cJm��<��6�t����5�5:�q�矐�N��(GJX���,՜�{�3�Yf��Ȍ�L�'�o�=�^��;�)�7��M�(�#�*�I�Z�HC(19�U�yM��}�
�U��d��B�Ct긱-�ذb6E C�7&�B5�Ij�0��Pv�L�ȑ�4�ߩa�m�xt��X�8�F�=�&*����l��L_նX�T��"[:B��ٳ)�C�W"�����8sz�Q����qp�� 6���O*њ���c�[&�#��*�\��I}c��Ks�;�_=�~}�7�-���y��흟W�U	c>�W'�H��Ԟ������`U'jc��$0Y`k�Z�k_�3��ҧJ��L#튴�8�75�}z�f|�f��b��V�6{���Ϛ��I�ı���D��e�`�������<�4�*tN�/�C�:���SxѾ�F
�q� �"��i�;��$2F'��8�b6@5�`s)�Q��X  �
����$���{j5TOkT��z���E4�{��cU��Fśg7����ճ/���l{����û��v��k�� ����������
�6.��+X_��Q�V�-��^�>{��;C��4�L�|s$�v;�~rA�9��)|�7��wߓ��$�m9��jr��{^=�5]rb�.��S|�i��b�����[x�l��|Et	�JZ=	,0�v��2X����U_�Ys�՜�z���5x�������(�@�[n�0Pp%�.G����R��ўf<G���.��J�

�y4[cܺ��nK#>�..<ΒI:oaQA?Q�QO8�%��B��Ǐ����[�g���8�W�p!*�S�<++�r���>��4n4K����� ż��~�F�L*rqqQ�H�g2hӰ���
�r�~�3�VOQ�76�ȃ@Pdh�P�0T��(�vɱ�	:���Q�g~g�h�y0��4��9�řc^��;=V}�l�J�m��in�d��|%D4���	/S���8�C
A���L���Z�����<I�h�b"�8�&�e�����������U�f���A����e��`�k�t��L&i�:�J~xX��b�>h@���l�����/��t��6�Q[��KW������=88�\���٥�|`*I�$I���픎M6��ʶT
����|>F���׮^@*[Ə�������T��L�
�	;�KV����}l�/3(9�l=w��B���e%����ḕE��mP�`d�jy)�Z�I|�l���߬+�cw(��LLnI�cK&1�����V��99��
Wv�rl�Yc���Y�b�����E���)��t9�竲UM(שK�z�0�����L� Kق��5[�ܒ��)�w�ѧD܂���fsERk����6�<��%�\3���r>;�`½`��5�t�>�<S�S�/D�\�by1B>���"�-9K���>=F�zJ����"֖p|@���5����\���oE��v�����[q�Qe����x������j$�8�y���{�/ �c�ع��UC_��?}��^n����z��f���￉0 Z�l=�������Oo����8����'47f���p��J�X,�̦��u�"��Cu�&<������#*�����ht&�.���*�qS0�s��%$��9J.�0鰫T�X�������9{\��Q�+��Pd�A�(CEB`�9�SD>�Qb���t��3]`:D*�D4��-�۝���n��":���$���P)Ve��>�2O/-��N��*��:�iB�������*~�aH�d��a~
pC����Ņ%7�3�0�Py��L:�66#TX��MJ%���U�j3{O�dY�9�&��w9�A��!G}q7��CL�!�଍���.I*ķu(Q���~� �B��	Lԟ�l/M����˔�s�..�X޼�t3"9����C60F;h���������qlÑ�d�c^�I0M��N�B�F^�ϙY]A{�!�l,EcBd��]*PE��Ƣ������nS����,z���&߃��l|eP�`0�d�����i�A0E�����3�)�h��� ܷ�~˫+��Ĝ,d��H�����;j�(9��D�o�k�R.��勨>�t�o�}Q��緞a{8�����d$�c�]	8Q���t*
�1*��R�|��������JYD�
�mw�FnvK�	�Fs�\�>�-l-S��U?[D�m]�1�O�bW�����߭�5m���E_���8�A���,D$��Q{Y�Z	�̑!͑�W�7ڇ�ny}�e#?J��{�`��cλ9`��L\Ʈi*�[�_��>٫���u�J?���ČCdH	$�d~�ӈ枑��$��)9�#��D^��:���D#��T-�L�`��J��%�Ì��CJ����O�P�VrX^1��N�w��9����;�뗿=�v���$��+������t��a�N�v:[ �lV����W��t{/D�������;������	���f(�H�b,UB��w�@>�8�?�:�o�P^@��������8���Џ���(�y�qt��fE�1�g��y贚h��j֐I�Q.e��͍�������K���Sl�P��cϰw@�,3WF�?;�)��Pd?_��m�
�d9��2�v$i�^��Ó�|7{�iVG�)�$!��
|T�D ��C�c��5�^o�[_�G�e}ƌ͈��;w�<*�9sk���E��w�꯲�-iw���nbkk˄}TEQ�F�d�<�� {�Y�˗��(��4����(5�E��l#7֚s�X��X]]>	�S��IH�!#_��U`eR��rO�Uf�"d04(�q�F�/��(�/̘b�鐥��?9��7W����Y+%#	��v��tGh�X!���L�)9�rOr諗�����d�c_��g����脄���3W�X`��4yA|��ST�d�xH��(�'	1�&cj��g��(9Ba??�O>�3�x�/.a>i%OF�:���@� ��#L�&�f�Tð�l8D��$D��7�xC�?�X(#�t�:ݶD48�� ��>+A��?l$�n��b��׮^F��s�VW��so�z���[u%���1Iꕣ?YΤ҃7��2F)�h��JAz�*P=�b�\{G#\���f����r�9P���Y�����	�7+��UU��U��m�Q�uaH�)�im;�cc�����-'�vd�d#�������D���d'�C~��v���c)H1kJ�j��ю����Z;;=���(Y�rH������v��N�B��d(-r"{	�$8YDC�B�%8���.I*`�ܚ5�OP�IH���Y,Us��K��=�����b��\sK�2�uǘ�*�*���nl\����lg��B�q��d�:O(����nw�حu�l�iH��f�&���i�R�)����%E�Z��s��D~�t,� ��S���9�Z+�����^( �o�Z�a�ɠ�+�3t��!k�bGs(���(v}"fa��g|rY,̗��</;��h�&	P���"n��ţg5ĩ(��h�EYO�S�1���޹�Eۄ�����AjFR� ���F��n����uk�OۀR�J�|}"�cB+�`�͇YbF1�'���C�pn�5T�%�V�p�� �`K2S�XC���A�4�Ӻ�|��c\�q���uC��Ɉ84�e$@2��6��L@��a�¾�	Jp�Ɗ��#%	7�|/�˥}�Z_��\E?{���ŚTU�z�F��Ϭ\B<��87�.w&�vDmd���j�^5�Y����
��a�,��EƤA�ɨF��A�?B��GC�26�z�eLů��c���Il�Ȥ��������a`�<������	1�>'�����^ҁ�ޏ���d�D�XU�������$8a�V������7sIh����ɐ��cY���f�/	ǩ1�=�B�L۠X:=B���|.��W�
9!�Ą/��ѷ���v���?�ҩ�����n[����=��y����v�ɵ{����h����SUKd�{3��'
��4��W&�=E�.��^̔dK!��Ratl�"S��D��$�9�G�r��ݾ�ȋ���;�?lg8�J&z�{]�e"�j�?�h9A�@�|^�7���J&�ƀ��d�n3"N��¦{�\�$^r���([1����-&la�v���FL���ɽ�*�3
ȸ@�����	ّɥ�`��FI{�	/�-�V���������p�kƙp{�m�x�Y��q�J9_h�o�+��P*�qpp�s�큕5���Xaܝ��Ҽe��D��>}�ʷ$�μ^��/�~��Hݯ�zx~�����=�;�J��.&�
�o\���3K�=��Ǡ�'����{��!}5mN��N-��l6��C|�����'a�/�>?��4rDMa�f޼ro~�<�i�^Ms��T��PU .�Of�H�;/�A?��3 F����x����f�z��~ܗ��+�Jշ����J��<��ND�P#�h";�9�F��H'v��B�k�ˌ5S[̇
��d�%	>�Z�=�+9Ax�Yd���o���M��)G�(��8�<VW64[�`+ȶo=?n<	����ɵ�%3x�ʤф�ؗ Gz¨� �Y� ~&�
�D(�Nkf�H�i1��!I��tc�VVdƤ���`͡Ul�����3��6\��>���T_ɳ�%�a#��x08�v*�R�&���1����Ì#K�Lf0Ѡ��";?��`�F���x��{�T��U5�^f��9Z�Ɏ5�=����ʍ���桫t�pe�=�[P�!e$H��Ȕ��q��Tc�'�]BK���&B��Lf�JV��|ҍ�����+G&�0����F��6e)�x3�\H�L�qAz �fs� ��_]�?�K.�G�Us�^��`6h�U-%��Uc���]|��������Ο_B��Ƈ�F�;�zs��]���BN�"�us��.�)�4�v<9�D+�fD)�c5��Ս8l����L3H�2(�bH�#�;{�"*�r�9���_��a3��^c��ZI�M����$���d>�<�����c~�\wR)�W�"��{�_��������|ȄS�ޭW%�b�'\��.~��VI{��[c�'j{v_����-� �"BĪSA[3�6>���kN�WL��aG��y:ak��Zt��Q�Đ���WeQ�hP�f����9�!O�V�����Y�,�4��?��ܼr�[ly����1�6�Cn��h���Gxv�D�7F��Ro��iʥa:����
֖r�+%
>�b���EԎ�8�Qku�|8�|%@>;F�?�G�^��<��Z�xV[La��Y=�f=�>~������1��	G<�fj    IDAT���b֯��h����(��ʢ3�����襤��⠉�㶂Y}<�2�]���J2$L�e=�Dd�L�����z�i�U���cu^)Dyp��Ii>�I��WV�U2S,�x�}肭�F���PXE�;{A�ӄ�	�H��/�>S۲ט������e�)5�Y�ҽ��q��"�:1��ef�Ԭ��A�}%�s��2s �Q�u�/TP��P����O�*/I1�Ad��Lt�]��*�D+A~N��s&6��5Slnt�w"�el�'����3�	�"��`�eyV���*&��$��u�KZ��1"-��Ĩ4��ıE���q�����u�������ͨ њV�eei�#[����N����kZV$*ڝY���I@?���1�r�$(U�c
�yX���"�������pt�ɨ� �G.������[o����E�y K��&�`���r������~��5q�E�?{�;w��8V�=n���m�;sx���z��`��l[�lY�2�2�R�Q�6�+������2���)��`��gp���د����v�Zl��$��!b[�T2�7� 7p� �"!�m�&i�D�$Bٳ�_H:�؅�`l�W�B	�Uʼ���L�ss-,�ϙn1OGj�9Gͳm�L(x�Ls;I��9�*�h�ڐ.���$���p��O�G���h����
IKY��$	��?��K�cR�&ɫ��4?Ϥ�r��R�������z�z�:+x�.-�iԔ��ڑ��� �եU,�-���>}��&ض�O��A�����g�Umb��Sp�;�co���If4�tQ��2�ǩ�Ν-�P�)�M��8����ė�����3|xg�o�c:���}Q���d� ��dD�� �{�~��U���0�&h �>�G39��P�!Ȑq��	2Q����=`簋��.���'���U�F�T��KOؗ���}�R�R�9�^�mHB���lK�9z]���I�'9A=�Μ=�r%/�_���������cDr���H68s���-�`IN&�lms1s�)в�`��{�e�e��3�#��{�h�4=m9PO�#����C�e�1J<��I�����0��[����|�$�Z߈��f}���Y_gfC���W�i�;i����c=2VmdD�%&�D���>��bJc���$���\`� W�b�����+;i\0F�ˠ����$Gk��@x�R�n�HU���K&cUB���ǪU��F̬7�$cg\�'O8bp[�?��k=C�V93��̭�B�d�'����eP\���}'��P%�4#�<e���&��B�@0�1*�"���w�����:tŢ>��L��R���l��M�&��C\	�h ������wO��������Ol���pӕ�#K��t$I�M���G���T/��4樍�I���0��qT��/vT��2�D�`��!gŝ��˞��x_�/�*���f���]�<I���6	nI�d��i{�l4/�5�����i
M���8�PQu��t��Ś�$9	U���Enū܀�Nzɚ�8��n�E樣�5�z$Cr:�e����K�s� �$|D���0�;'��%Ϯw��Τ?����=1�e�HT��M���Z2��<�I�P)��>��Ά=�2i� ��Q)���/��ܷ&ضO��^��ϩ���q��9��=�^�����}t{}�[C	���r���p��67K(WCm<���8(������G������?����%1�PX�sY]e۬^��=�9�3��/Q�q�Xl�0_�E+!�2{]#��PV��la6��=V�����4;$���$�g���,1��,��Q��tkٿN�أ#�;�p��8��qKQZ�@��`�6
5tO[В`{�ܺ�3�����٩��/�I�A�.����8���ӂ��ջ�f3T������;wo	6c5HC�7
:�>ӄ ��#�Sʐ�Ŭ\iL��D�(#�m͌
������Ã�+���R�;���V�&��"�lv�'^���8MǠ�/+$&P#mt���)N�����zU�}l�)AE=c��L���<P�Bf���Y��/H�
K����o�r9"��. �W�`�+�?��HM�Ȕ����%�I��0c�OU������"fdE
E��
�� %N�3WO��]�̜/� ?�*7.���c.������'�u2���Eш`71��e��j�Z.�w~�]�-.��5���|U� 8{��~O{�Ӷ9�ilP"LVU��t�v��bua�`{�8�/޿�f���(D��F�~$3�'�J�1�`KB!	S����m>"ҕB����}����I���EĔ1���#�[��I���Y�X���t�8��,�N�|�_�޷���bK,�w;?�(��\�I0�{*%��"5T���V��zc/�yCW�]�)�9Vpl��v��Hޫ�V$;J�:��ݍCʜ@._�qc?B���3�Y�9IB,�Zk��j6I��J��B�a�P񀐰Ia�w])V@�Z^�c�x�`\.��Ő�j&�Q҅�Eݧ�<�|��ߞ`�|�_��G����'5ۨ�cLGqVj����3��b������w�F�`q����2�����Q��X���o �M����������k��ٍt�9��Yvh�r�򰜌�(�C`���b���;.�|�(،��}7B<�Y���l�x�c������a���4eR}N�b�p�p��0��#�>��#���?�U��'��<c�:�)�{�o�?�a����r� ���H�@�Io���k25�������Ff/�U63jT�b�=w7���
6�*�T�<�͕�������۪�`;�9��d�,d�e�7���2�0�X�V'��ܔ<�%��C�����[ll�a�LT����Ɍ'bi��ş�z�v����u��櫆�-�&�e��ʨ%�h�X"��j���W�-a)4�#u��5�$R�k$��q�ȥ��/3*T	6�5N��m�j�=��fM���l�����|���S;q���_�����h�����0�T#.QL3���<��{ٟK�GV���J�
��������|��P���RNN�X$=��>�b<l`8�!�P̧�j�/����ͳ�L�~:��Ң֦z��!��9w�߳ic��Ƶʭ���$(�у�pzm����� ~|�F�YQ���^��L�fB�yIs�L�TT.UaN�`�-�J�$�Rk��?{GYx�yY���-��xb뛣?�ؓ`kd��~6�2����S�duN8��dM�l�493�lc5�Zk��"D�ڈ�b<(�!��L��!�h���QG�P�ZM�;!{
}�x��^��|r�9q�툤����[#�q�۾���􃵇`���0�$*\k	��*:���$[�D9�}�����/�"��$�@OK�q<B1��Z�圊a`���� u��<=w���^��`���E-xm�����/uokYv��{n���ŋ>�����L��T�(�U�쑇��O�Úؓ��˪*ðQeY�J)�)��d23��̈�����}{α��}_P6��I���@D��{��{������x $�����3�@?�6���Q�n?<������
�M;8>�ds�c�m�E���v�l��If��=+�gVi��xnv8.ٿ��ڋ��fY�R��Z��8{���mU�� `�:%J��X|�҅ù��� ���'��3ze�T�TT��@�xѶ����ԃYFw"t�"%�g&W��Td�@�A��{')���w�Du���!<�y/�^/�Ι�7m�r�5��;��?�L�VH�aDܗ"������cak�1#ڝ��z-����>��S��FK�-��U+ IW�b�)&2N;�j[΁V�R�f�}D�G��+�{�:,�y����M�p�<FUɩ�c�'���9|w8���9�.��6?r�A��������Nb��P�@<Qֵ
�M�̊dh�k"�U*@��橏d�Jhp���x]���pd(�糆0�=K���T�nL�йf�^7���3RF�^� �� �5�cU��F�$���u�?8�E�
*�7<�d\�`>���	�'#�q��"x�NT�
S7���m9?�Z� �w��z�����u����B�sC�����J��$MN��땦V��5����]���k
�g�f���돆�ޏ?��C�:�1��@<<V�Qe��ljd�LH�%sk֋��b���D�����u��=�{�2[%h����T��.���k�蒒��W�H�U�8gb_4V�q=��������V}Q"V|�=<Y�mDd��B*�(CP5�T��0!�BN��Z�1�9��V�P�Aw�t�"5|l�Pǐ�'�x��
aoݧ�û�]���~����u ����{y_�*��kU>ȍjŊ9=ݺ�[�N굲e&;��e�Q�?�����^(N}GI�Wlǃ{��|t��Y�R<���M�q,,[���b���|e��߶��Zju�̏��+Wv�l���v��v�Z�������I����w���}[�Vn�m�#3���B��rQ��uW��q.I8�i���D�E�����3 �:i@�1$�4O�����Tkh�%틍q��j̿�C���kG�oD�7[ͦ�[����*/juT��J,x����fUޅ�v�n9���a��_�;w��>��Gn �@�����˗/��
�yp=��X����Ū�t���Gr��z��O��+�'�-��� �L2u<=���n���=�c `d���m��
Ҝ% �SR�Q��;@�<#�'�M;II�0����0�`{
;y���;䷲�p� x���9�=��Y���A<Y4���;A1D8��m4�wԍ8N. �$ '��Hk�b���d>O���80�5AK�B�o���Q�:� ��>��>h��	R����qzB��$��V2�#0㑏� 7 ����k�_����F��Fl�lb�bj[[�
�g/������ݎ>�0������)΍�^��$���ܲ��4`�'>�����z뜝O���؞?/����9�c/����/�U� ���
yi�&�#�<p$˭�@b������NժMҚ��O�)��I�Ve��`o#mɽ#�Ft�d�^[	Wl)qݫ<XC�y|����m�އ=����<�H<9�LR;$j��<C���#z���:��4( WLi�N����b��I�&�s:��7������[�\�Be��#�Xm��>����U����Y�X��3)V������(���qO�w\o)�`�h�$Qܓ_1��<J��[���nm�{[����׾B�=%���:؞������y:+P�ALfꍢsi�Բ���RÖInO�ݱ/�޳�#`����f]�D���6:�^��m�ٝ�u����ڴR�g�o~d��~*Z~��e��Ś��Id<�5X��}�|j'�#����5"˹�9�	n,��#ӉMfSUf��D#��km�ջ�dP�ĎL�#e�\���l DX8��O5̢f�Q�m�_�X���
T����srK{�Ջ�sf�5Z7��Gݲ�~��C��!9I�[|��E���8�d��qcl�Z+F�y�6���4l<��P[�6�%�(z�T�@��i�=�r�5�A ��C��	i�(�LAͻR9V��>*B�H[�P��1p,�u7���,^	S��5�������e��^���ƅQ$�w$�����3��#�Qe��85ƹ�.�d�9:m.�A%��j�(�m6�T	����;`m��\@�3u)�w&�A�Lծ[�sK�9@{�G��-]͖r��X��#�%+��͞F�tg�D������Yi�gg�I<��B���X�n��kL�33�N �=}�tdY��c��S�m5W`}����{��Á�Ȍ�eh1��]�%��L�Xy��5փK����u�F��L�+�����o���=-�;o����o��=y�ľ��i{{�$��t��"��JR��*��u��@9
��[��5�=ϫ������Ԭ�a+|�i�P�26%d�h�RU��6�d�*��1܂��L�r�$¶�?"q�=����]��Z����������[X�[�Q�zCH	�0���m }�矙��^/LD�Z�w���-���\!�'��]����}A얚1(s|�
�4��V�i5|�wx9��}D�86�Y-x/i�`|��5k̈k�j�v66l;�Γ���K�u��/��WSَ?�WӮ��|�`�%�ꖯ&6���+�[V�$6�N$N�bo"�ۇ��A��� ������d�F�Z޹�작�ǟ<����&P荔`��7��8��Ru0gA��-cg���*[���Y�Y��NG��[�v��I�=}�Dd��\^��V��Z����÷U�
��ң��8X\���Rsqާ2��K�f�TV���l"�2���2
��PS{��+���	�~x�<xly�Y�2���MU��*O[[;�l�\m�A^=�t�`������ٝ;w|4�� 8�?�*�B��k#?V��Eo�E+����+�A�m"����®\�`/�Qb��s�'YS��?*.'�9�ĩ�N�i(i�������}*ώ}Ii�]��r}��t2�����s�L����Y�U����B%q+-���믬�/��p���	^��&$w	в*���+ �m<�K��;s�P����O����[��y�� &p� j�Yc7$�}�x�~I	��������۔�5�%�0,b���j��rl��uz]���;v���%�[�#U���K��^+�T�~"�x��0�[�k׮Z�:��W�v�LUJn��5���������
��h���dHJL��Va$���͒ժ�����k������tm2���F�K=[�س��=_��`�8��=��C�A^��2��%�}$��yPu� �T�s�ˇt�KY�n"��p!�8a�-�Yй&�E�G#g&"�ÂF����w�w�����~�\�B) ?q��U�.�9_%Ù{,��!E<���X���rКƈ�ڏ�`�$J4ė�Q�6t~r�@�R�:��U��ش:�~�����}�K#�Gw�ǋ����*�4�Cz�3��=�~�X���Fs�i��en��S{��؞<�K�Y�j�+R��s���pM\tb�����r���'�-�N+���
�B�
N3�Y�.qciTs�Fd=���H�`��k���];�ߓ��+�^Qvp��Ƴ�z<�}���S{z8��ܵB�ci�H }J�J��X����w���S�[p[0�7��=���nZ���-��el�>4F�T���y����;��ɾ�yo�B�\LN`�͍��ٖ�l_4�S��m4l<��O���fαb����h��2jQ��tN��J�`��BV�na���Q��T�]�l.�����a��*|}LE)�+�.��jB5�u��̼�z�B8���r�:B��g�|<����v��q��2�8��{r�RE��d�|oV4���E���W^���W�%y���^>P�_t����{]^�{��V��x+d֨�CD�)(H��_H�aMjlT���C�����G#��He ��P}B�A13�d��gC[�'���pa�&8@g�U��ʯ��_��6
�aw����c����g� �=M��s_\$����^}�+�о���mm$��`����?��u��W����������h_ܾi�*�l%��-ld�m��Z�a֪#l��f�n�ڝ��ju;%��Ǐ��S2��#���;1&�
0�� SqGQ!a��:�	�
#61�
�Q��
w���B�{�1��$�5!e��v�2�J�J)���G����T�Z�U��,�s�$�AŻL��P���_c� ����^|��A(
XD����|��pj��r�9B�POg�cP�k_�f�_�W�V�y� Om�:K��\�d�3��D��èf�bgpAc���z��U�_9�Տ�o��K"W���_[��Y��o'�{^�V��~�� px2�g{#{��������˶������	nO�"����r,"�*��r�Z�ܱ|U��<�    IDAT�V}	�c � R�����v�{b�Nf�=����N�LG�kg{K�,�@M�d,Hz��ڏ?�o�NVj�X��V ��f���:8��jA>�Pҥ�����>�
�h�%�?G�xriB���]�t�vH��-{�	�-�f�
��W^�3gvmskG�y��ؒ��~�kNL#L�o~�Y�ѣ"`�˒�m� ��-O��p�
�!Yα�}$��|N�`+X����K���f�Οݖ6q����4����S��E|�����J���"U�����Xc�Y��_����Q%����ݩE�Z8
�9Vm�vdR4!©�u���lY�7���o�b�h5�|!ש�p��c��I+8�+w��C`�1����� �)�KhK��V�N�Cu���aM;C�UQH*�?V2(w&O^�\��y��j�δ	�9����
�Ȗ�c���1:UǠ��8�`{�ʥ`DP��NO��x�N?�^��	��/�l�|���8]�xޒ�oo�޴Kܼ����7���j�/߰����͟��= 9@ƿz���ВK���A)����5�Ӭ��ݪ��F���Ǚ}��c{�`�`L	R_��$�.9���E�_9Ĺn�^�=D$��0R�-�U�&�Lx�5�_��($N9Ly@���_���f������ �"�Ҩ�be�ɨjjX]�|�F����h}��WR4�	���I��뾻�#낵��LN���"��X�ƹ�3�D�e9�Q�GA�#$����5�\Q��̂��F�(�7	�z�jG�D(��.<�j�v��X�\�v�����y�Kl����ǷV�ūX"M�����6�0�mu& �6����@��ş��2����}th?��Ͳ�O!5�"�F������,3�-=��e���O�`���u��U�� y���Uc�u:m��mZ�-t8�P'��@��bJN\��Ӷ�[V^���}r8�����}z�ЖŎ�xG�T��2-pA���UQ�3V����Ϝ E�����4���Ha	W���m�%#M�\"���G{�N�̀	9�6�z�k��E�
��?�o����[��3g�ѣ�� +4F<�X�Z�u��5c��>OSӽY9��,�K��}7�F� ��$`���j0����~�6�5*�h�pfӑ�b����OpA��ak��6(N�jؘ
���@�̕ۊ'^�r�D�T�T����F�Z�L_T�H~pRp�~���e��T���8ʡ��
F��Sqg�?�ONap��%wTb}�c�Q,T�B u�Z����""��Q��������S�<ز�U٢%�&����9 �lw-O�\�c=����]x�%a��n��k�snW�DUպ*��d,�(�Ub/|`k�ʩ�U�Q.���6?�s�꯽�������Q|��]8����U�%fj�@T@,��Ԫ���&^Z�f�ٶ5k1�*JAj�j:��$�����`m��%��E��^osmD�}WАZ�[M�����0��G��c���Z�l�
� t92oi;��g=뜩�����:ЫlX`�K)ʡd�Ϣ^-k���o�����A��-bU ��&�RD؜#�>r�	FU/���l�+}zR���A��a���a����j�e��/ElJ.���U�ɞ���G�W�Y���foKn��|��[7�~iz�y��_|r3����F���Sߖ��[MC�N;:|b���%�붱+�\�LrI�N�f�����5{�`ǣ��34Uk"p0^�c�t>����6�qߚ@f�2��m�j����-Z�<Fs�%w��7��HV����Y���ut�˙�6Z��w޴s���̓Qn?�����v0�leM�����[�%��3k��R��@[�
���!��4UOҐ���d�7�׉�#��:��@
�A�G�_X�d�@�U���z{����l��Œ��:��?U���W^Q���o}�4zA5�s�2�m�nI��X�LrEU-AWjTA�C��X��3a�3�D��<#���^�G�RiAؐ�[ � ���s��H+�l�6&�ScL^�EF�8t�`�k3���
� ���c�!��*��[�$��?A˟#��C�ÍĬ�h�|1S��ć��*Gl�&��DBX��5j�{�c"ܛp�r��Y��a���ձ��>�i�"����x`B?�]�HP�z���8��`��T	Da6�2M���rGah�%�p'V,�����4S�(��4�7޼fݍ�F�@a����=g��Ԏ�to��e��0<Z��U�sZ+W�\���?#��o�#�����;9i[����% �y �*��h0�S��@�
��0q{N&ؖ!;%������*x�E��,��- x!P���6r���y����7����L�Q�|�?PU�,�j��Qg�]�
܏U#���A��t��X�*ac���$t!��`m��TnE��`�B�G�-k����ـ�iv6�ђ�F(Ys��n�%U|��#+[�,|�J�S��%�6�7�����ѯ�4(�-&��v����0=F	[�<\�x�l��U��h��s�m*�/�������?+d�u�$�u��O�A��Jn����%��ڝ��:T2��{|B�^��4��z�}{�����3���lA_�U ��y��L�J�����ƶYַ��P��ika�ΖͣT� 8? c%�P1��D˧^.���}K��}�׮ٕKg���&ne�f�����G6^��
Y�\��	�����d�Q��D�� �-K={�6�d�S6pYTp�p�[�gFP�|B���sV�֌�Y�O>��#Y㱨���)��"�Hp���0�7��M��cV���9��g��cG �L�K���V��ܱ$ih��dG2#?
�lcfK���XD
���"��۽��"˒��^��[��.��1�9����Bҗ"v��6D�Ħ`9������	��Ke�1�q�9�~11e��Lj���]���-���99m Y�9���� Ea�W�����R�f"@,+8���S�:Yə��&��"O�4c�T���{��
%Q i�P��D�х�ܥ +7��[�E��0����{�+LЗr��;ć`+Y�׉Qȉ-W2 ���T@�mlO�H��iao�$������Aᨌ��@ɞ����e�I��4�΅7._�d�Oo*�~��oت����oڣ�TL?	�U����h!�E��Y�!�l{�V���t�z�ht���ܲ��h���M{��`���t�a���1����i����\iI�����~:�C��ƺ���5�9�`�Xɬ'�rjf�Ps�p_�2_0����-��'��Q���r�!7���ɬ3���(�#*|��fz>
�����U��Xʼ/ݟ�XBW0�e��8ER_�B#'�׫�m��5X|�����)���Y�[9L&�ؓbyZ���ZU�8~�۱��r��o�K��o����ӿ%ld��������喇����de��R��P��I)�zy!�t�����塵:���z��/ �4~�cзg�G��|bO�m�Um�*؄QHt�ಒU�u*�ݸ�ko�ֶ��Mf��I�;��aj�ζ�3�y����.��fqa�N�#�\w�%K��vJ���s�l6�p0����~��-{~0��
-b�B5�s� ��Ct��}a䩳a����	�O�	)2Kzu�k�sA�z8�	�ͦ]�tY���Z�~���5�鐩�U6�6E�:�sV��%}%�t���T��٭3
��n���o�b�fD(P^j[R�Eﵮ�-=�,����E:�����M٢�iխ�,	2����~4$0��(b����
H[�!px��`R�X����^I�M2�� Sͫb1��]1�!1a�(2�U�h5B^Q�_��T�۬F2�{$��S*��X����,fK2���'5Wf��3pQq�#V���X����ߐ\�s�x�u�xU^�<�#�;:b��K��_d���	�$�`E(���\@�	�d��s�;1jq`��A�IBE�\���f��W.)�\wv�֖p$&��h�+��W"v�C�R�z��=}������;����������S�{��ҙ@j[
��b8�`K�P.'
�H5�m��A56��͞%�knl�pZ����L����V�X��<��bj���g����"��hA8¯�G����g-���E�Uu����B%K"�6�V� �]V`D�#�l�2�@��`˺��n���~~ݐ�bam��@�M.�Ar�$/�Q=~'�N���^h���v�'V���5�c��&$��z�H��3�v����	�T��Ld�Y,���^����6z�5���`A���_�ǯ,��}�/���?\"����Ǚ����E�@}fa��B3��RC��I�o��K���>�
�Dޯ��4�0:3��#����j6]�m$���28؜��j̿���׮��W�6�=�<��d<������ϭֹl��"H��#��ΨsSa�=P�k��V)�v�®m�Z� 1����#��h�V��$�R^��|X��\���A�0��0	]-AP���+Z�1Jf�Q�QM��!I��lԤu,����7ok>����|ލ��ܹs��uF$ �K����x�@��ٰ��}��Y[��t��W�Ҽe�P;�J���F�hC��^g��ph�΃m�G�()���g��&:�@��$"���+rS�@5�Y�F���Q�`+��P�r�}�g:�ь��W���TL_�C�,r���;�3I��<!��7%���� Ʋd9�������K��1�2�8�!,����0S�=����#q�V�Aj�P��çw�Oy�分+k�!<֕*�����@^/[A�Ҧ�<�j�N���B����f��#[,-]-m���A������^ѭ���Z��%������ߚ�%�U"ָ�Rro�Ү���=��3+�3����W,����_���i_�3fO�O�-O��`�I��U��Wr����m�)�h�n�f�����wU�.[���ٓ�<[��� �dv=������{��~�<o����s=��DbU�U���P�g'k'���	9ױ�����/��R.��Fr��`�%����b�������)ϙɬ1�;��:�0� y@�,�Oy��!'��l#�JN����:�>��q��h �VD�<��9���j�G���\��Ҳo4���u�1������~y������|��P�V�:��rwґ�>�@M�vcSڥ��AvRs[LS;:Xؠ?a��Q�N�`�N]��7�ط;�6��9K�i�Vn>�&3�����[���W�VM�G:�x��c{�dh��e[��M��0��.���ۨ��2���[�3\��UHX{����'?��C+�:6�ZV�Ïv8&
fÄ���2X�-N�N�ߠ"��(ܸ���K�)�`Q�I
:P�pgϞ�Ku�~p��`8MU͙à�������s��Z�E�.Mb��l������l<:	PfA�6+���#����pEF?ڡX`d��#���MM����a�ڱt ���������ł� y�;�͂~0*�<�W`�}k�����Fuy:���E�H,����� W����&F��P�e��Xt��t�"�B��
b��]
��J�9bU˕*�
D�2.�H��HG<]�����`;1������< &R7���c�ut�ۉ)28/��Y�d&�sX3��v�\ki6��߂��7P ���嫾�R�dO�p���������]�~Mp�+q�\`��t�F�_��?9	l�~��[v��Ƕ�޳��'_ў�W��6�w��rr����=K����x e��*}���+�٪o�Hls�c�fɚ�����qj?������V��JA[�U��s�"-	��1��gx1�c�%���\�
w�YN���ˤ"�<�_̓�\�!��.�b���ps��K�b%�"nKh �%=�3�NX�~>��D��X�a��u��u/�P��`���z�gP[�J=O�b �ńcG��{�eN�/�X��^�f����X�ʦ1������f�r�k������������=9�蟭�
�����!=ە̓LZZ�x��bӅJ��c��Ԏ�����ck6Sk4綽�R�doj����l��Jn+��bw6�Z�h��`g��v�\�Z���-�bП���-����8�a��3���:A�7�
-f��3>���;v�Y��H�̤��"��Y2/��<��Z�;B;|o�$B:T*�H84�9��\-���^$���0���'��	]��A��� )F'�7���՘f���2߰G��|`�I_U������͒�W�9s�h�2�L��g�C�7� �$��4��=�?؝�ԏ�X��;�x֯M)���g%��� 7��TUO��`�����+`@G#j$�#ʦW��s1�cͽG!W^W�� {��!i�g�1�y����U����~o�
�&o]gNG��� �G��ǜ���	�5	I4�K��O��������`K���Я���8��G�� �-�,�Y��:����<��[��������oKj�Y�/ǍD-\'������qT�	�1�2�J���g6߱o��W�ٟ֬|�;v|���V`�.�|h���X��B� UoB0�t곲J9�v�j�.T^�>1�?}l'M[%�_� M斑���l�9��Gg�~XÁ<Gf�D�Z��_opHՓk*MO�H����E���e-�:$�"���B����������)e��-XW�!/ֱ�[ĶS4B q��e�a�Qg;�Jљ�p3��W���sv�s�sq��d$�<b�a�X�F�I	k�?����[&�����K]��l���Pٲ[��*U)m9�\��o����Ue����.��9L���pi'�T��>&�3
���6�e��R*qPN��L�32����j5 G�b�ԫv<H��_����RK�`;�	*�2�_��/�.J)�TZH��Vm�r���%���/'�E\��ݪf��g��K;�u�E��J����6�5P�l#~�A|"`S��̘��ժ/��>�3������������'���[b�GZ]��v�თ�i�k���ҕ�bs���SM&�y!|Tj�lѕ�����r>V�����'F�6���Xݬ��jF`���% �!�뺱6�(�*�׏�~Tp	���A�|Q�Y�S&�����`Wܳ6s�Z%F����"�؍"��|k�F��
9z��W�T�T{
��S�I;����̟C�Q�`t�����������d���%���Nm�ꅬ��.�v�*���b�^!�g�L�u�1��3B��^+s��@y��Qa0k++6��4�U_�K���/�g�W�v�i�5�B��O�B¼Z�X�<��S!jwe�,9l����[����7^�q ��@U���aa'''
��N��ЦOH_���k���g6޳���;Vm��O���v���ȋ,��[� �N��XBz�a�r	q�[�<��ulw'	0�f�xϞT,-uѨz�������σ�F���lc@�ǲ�I���$�ZX|���L�U_=h"�z���X�]�@��Yk� _�ڄ��D�S�9��fR�������"+�X}�ޢ\���H�D�`뭰Pه��X�ƹ�l�ѫ��9������u?Z��{:�*b�+3˱g��[��oS�r��oY��#�j<�Z���w޽�˪f_�=��������?S�]ev�_��pa���WTw�ҦK浨֪>�� 6��9�/�%ib�v�ڭ�Z�`N�Tb��`�an��M��3�=K�����Җlr�5lC�g
���z[���w["" ��I�k�����V��P�P�,��;�K����6��m��E����#A�_a@l�@�ID�����jc2qD�O��>{�`|'Ɉ=�������f�>s�����}�(���~��j�9E6�j�F0�$
@v��v6���g�������f����u�XR�Te(�ʖ`Ke��S��X�3g��t�uiJc��
.@ޏr�������U`��QbGB$�ŠƤ`B���`Io�W�    IDAT�D��
T��+jS��^��>��mG0<	r���BN(�S��p}�LƘC#A��6 �ཐp �>}�\,��@�� �D՜�QA 8l#��^k`wƤ�=�I�d�J5�1@��|�ة5�2ZF ���W��:#5�#׈��b#���U��g���\��C���bHu=������|�*�3�ۖr���ٽ��
�|O��I�tgK�C����w�`�s�����5�u�?��7vt��DGI(�}$�)�� 6r�sB�dPP���f�j� 0f�6,�-��~n�g��{��<�7O2�Z�D/k�х6ld�G�\*�p?_���9��;6���g��z���kM��D"�y	.0��S�T�F���U9<<��>�:�i�z�9�2�A�����=pZ�`�9)�Ft��	��>N�z��}��������1��w�w�j��ǉ�}�^L��zT�Z���b�����K�m0�\�}��m����4[��+ش�`����"���A��д���5KɄ�n80rY�t��Ҫ5k�uZ���K�������s�w�o�ꆈN'4�Ԏhe���G}[-�A�����O��j�r���Mt9aQ@�M�uˬ��&N��Q�Anp�9�����n�{(E��
Y��~�K-�vy�Ƞ��T_洚q�%o�y:FT��R|$f��H�7Tt�/^~U�맟�tvk8�y]4�����s��s����D�9ن��ܙ�
�����٨�͎�KJ!�U!޴MY�1?A���~��p�.�y��c�$�>%�oa�R��kT�����"T�Ő�(��P�d��������=[��xf0�%�����93��K��E�i�O#�S�K�s�3t��A@���~����a�Ղ���b$ N�8�{^���?�L�S�f�{Z:��,P����aU	k?�@မ�����ޞ��N�/��'��5�ly~w�?A��?��W��B�?FC����)H��/��"#�"H��������{���~�w����e�Zw�$y��2_�T�!+���Ņ�K�0,޺��=�G?��o���:u��?����iOl����3$�R��RT*���lY":��b���j[��Y5�������ݾ77�nZ�ְ�L����sx|p��`����9�8���C���/
��G��)9�PO������cqF�q�Lœ@�>�[�$+��'s� @��`�0Fa�u��ɬ_䙐�g�T�gA��s���26����X�эs�����gm��ݙNu�u����=�hX��&_��
�l�-Ux��� ׌`KeA�ʶS�}�*����<���{ 'R�In'c��/�0AU��1Ė�",:t�Cu�b\΀J��VJ(Mͭ^g�$�n�4��ᄊ1N�����4k�k�H�yL�a1Z�!������sV�T�Z�H�i>dCc."��r�rԋ��I��8�}nG#�r�bU=_�>�H�x�����I_C\� �8\��U#*|}���9�B�ς&kS��ʫoسg����u`	޽l�/0"x�W�/A|�\�f+��\�[+W���=�����U�;�ڡ>^�,A=�kyFeְZ��DF����Ҝ�om����l��-����j՘�c���P�E��$T���DR�&�&��щ?��r� ��/ʭ?9�L�j'���O�;�>�Ku�^	�Zfv2xu�׳A�6�Gx{4tK�j�H1 $elA!6w����Сj$�5��P�7+9>�"�8��{ذ���#(n���1�j�Q)�p�]��4�J.�Kg�=���=�y�KvC�mG�NN�φV*�#8ё~m�����땢ƅx=d4y=`�W_���@�6j	��r�y�[�TbE����~h�W_{��������ճv���������@�.>OB>�m��Z9��M��b�P�ehk\�������-/.d��l�޻ew�#'p?Kab�t��+�,U��eHR"�II���bc���d	7#�W"!ًATb'�*1�6�fJ���g%Β��8�Cr�}����ע�8��ƀ�gh4�(:�S�F��g+�r؃�G����k��&�j��.��բ���aooO��Q$OP(�<�)��?�9
f��:(�T9�^K)��hb�UŐ��V���7;��Lg�۝έw���fD�~���`�����`1>�������4���l4�m:�-���6��Ќi���qI�G���L�	�����2�WƆL��T �����X
yQ����Hb�Jj�ɉ�[�t��ڠ���C��{:X��l" ���ryl
m4���B*���*��O�ݶ� Z<�s�U��X���BV0P	�*й�\C$�E#:H���D���-y��UkO0�g����=�\�Z�X��!�\�xή\��jW"��JL� �f��ݵ�~�#��届�h�S�c���_�Ě2��v�z��F�������SBx��B��p��C�x:*'i#�]��{@a,�����q�}� �a�bY
X^ҷ�y���0lJzQ��n�CS3wh᠈� f��H���" �"�À@�f3��:8��*�8�7}b~3�
���[�X���"���+��e������0YAgP�&����s���� �1�?�?x"����!�*ImUk\�:{l�-�ELבKd��Au�%�aCK��Wǖ.-O=c-�,Rf���o���v�5]?\��ˣ��>��:\��Ϩ7^��R����@�{���G�����������NN�A�m69QM����"hy��j�R���W�NR`�:m���
啵z�&���w������m�zM�?��`�XL����'��5�N^�T#��z�
00�^H�9D{�$�99�t����?m
*}��V��T֑���=SO!��8�b/TO�Ǽ���Պ����@#�N����=1����G���pc��߱JV-s%1)~gDs�o�����N�}�t)g��s(z����*VQ�lYۜe�)�c	��J�`ۮ5l����ݷ�~�d����ۓ/������X�MK�2c�s�0�LSU�n��,S�\��1	620�f�Ԝ�>�m@� 3zm�|i3tY!,dd�.W��]rhn�fѶ7f��dxd�<��F�*��]�O	�f�bU�(�k�#19� �����xH���nf2Q8���֝���͇6]���rŦ���tQ�����<��1��E�ߘ���\㴲�T<�B8�a\[�ѡ͊����sd�9`*����Rb����!�r�-�F^�K�6_�f���c���M���B�#�Y��Fް���Q�*A�K���ӯհ�����>ǉ����_Y,�p|OAʐ��!�#6B"����ܨʂ����%�~�r��ޗq"$3gUN!�2v��OЂ�a��mHD��T"�>a��b\�� �;����0Z]�����xy�3{*M�0߫��X�޻�wX�IP����7s89���׀zW|���_�B���v�d�[�ל�J���KW�lQ`Jӡ�k�X��T�R�ש�^����V��m7n\W �7Ѵ�đ������H�R��	�������=�����ڎ����v҇�H��cC2Z���V��v��-��rj�݊u[ʐf 9f��C�<��/�6����Qt]���]�-������<C��2�p�V=��O�}W��������h���j`&�L��\s�#�Ą���,��9EI��D!
)��U��G��[1<�8�� ύ������{�e�mA�B?7
{����woߨg�>��[�A�"Lf ���"�"Bʞ�x�� ��/���0J��H!l����שlw:��o�y�+_�`;>������=Kg�E��x��p�ԻX%���&SU���8Ԡ�3.�^.������RD� �`eaK+����/ Y�؏Iٖә�Kfv��ɭ^�[���x x��ّ+�|��7ZƸ�xoe8~έ?8��ڹs�b�B����u��������'G�cZRW�P�90JB����;m #�j�j��&���LR�.!��JW�UVb�m�U3������v��-�4#��/x�<�nG�v���:�Rq",�
�%h"�Ѳ��޻�9L��K���$�/7�Rݰ�#F�A=�����-kw��r���Y�s"G���/�&�71'w]A"����Ke�#�d����W~��-CV�{�ڈ�Kz����{�^�D_#A�=i�(8��U���SՃMl�yzF$R�+ t�^�k�Ȧ�qv��j�0[�PS���z��G<��<�HO� =A0��C�s�|�@RT�k H�ߥ>�<���|�d��bƀ(@��������f�n��,�����,)L�}�#~�`%c�����ݯ�#�W�+��gP)!1aJ��X����!�P�l�=�Ԯ��mg/l+�Wl>��G?��1�7�1Lk�ϋ���f��ܶzT>���mk�i5���5{�|j}��N��6�0��G����^S��lyQ�1[�l���d�,�|_x���[�&��L�X�uiB��_Z$�9l���e/�A
 B�ާA)�ޥ�$/�\�ڑ��y���ft�bb���IR2h'�������yO7B�T�Pp�Ǌ^�Ԗ�PW�,z-~�N��3G��5<�z��d��3�Y�>k��I}Z�5T�8�(؆���o����_�`;=�{�?8�Y�����S;ҿ5+U����P}<D��d�1腘K:��C`2* U�d=�@0ue�mУ��Rj��銾����3kTgV-d�?�9<ˋ6��`�@g��\B�#+��|,���g�h*c�a2�to��<ٳ� ��$�R**#�;$�㐹�/�/!K�2MX��DN��{�gt5�S0�,�^h�ݶz�!��ٴ�w(��s]F-ݍ�z�[-v�P���U��Lv߶�����\!1[��-�v6�TٲjeG��Y�BxU���;i�vZ5��X*3ň�R)3$ý�e�(���pZ���,vv�7�/�m���fCB��Z'ArQȯt��� Ar��Ug����\�vz�=�Z�$X��SP��$%�&��KQ��#�@�����\�'O�ĒY�-�xIBR>��,�����O�%	P���N�*~�đ�����E<�4�ɜ�l$n�q*Z��au"ǉ�������MF��ex�-E�by�W� Y�-�k�u?�^�5[ޗ�J0���ǵ 1ar�JE��3���M��������+W�l�\���[ߵ��Ħ�5d91d^?S���U��x��eY�FICЪ�mo���Aj�`i���=�/Y�v�X��Y;*P,�w�,�YA%�l�<6m��!���b=2�DX��U�����Ց*��Z�D����*U�/�t�\�z��V�T��q�`�s�$�Z\�Ο�u����#@�g	�o�������j�l�x��C+�{�^Ism�
����;s�8V򲲎L}�FQ4$�d1at���:���nT)LX��p��E�\��Un�;����y�Kl���t������,�;R�/N"1vSc3]I
��x:���[z�E�F@j����꒢��C`d�񥚕�[��Irv��S*�ls#��NjMQ��t���pn���la�y$��U�U��̶w��Lm:����b�b
��õdG'c{��=y�\3Ĝ}�X����y8�=�zE����bpǉp1�ez��@E�p�yBH��{���.�7� ���g���(�R�+�x^ockC�(�m�ӕĭ9&�R��ۧl�~��eT_�f��ٮ�la}���M�-Ǌ��mH��l�~w���P�B�����R��z�3uV~�lL6i��S/��`e7�w�g�3���RP���ٷ��`>K��dQc,QQ���<�޷��ҏ�ʃU�j:��2��D�D���˼GE�$�}�l��~�p2�I�q���PF^C�T3v9w4� ����R�	���m����������	cT����
���0YpC��r�^�Wȅ(~QM-m8x.�x�kWR�:����s�e�R��T���~�W_�����ZE��`�����`�3�"枸�~p$B��Z��.�6<~d��~ƶv;���-{�u0�C��̓B[��@r���-gV���Ɍ.�:%�h׭ݪ�s[��w������̞�W,�nل~8s1��9Sٲ�X�be)����YnK8q��c�/A�������'��ȭRP�	6ҏ$zb'W�G_e"c�2�$R���ɍ��B��W̰�z$)� �[��cm���/���$�U9=A��T�z�K^8%Ϝ`*r ��0��>W1Fc�,"��^ˮޅ��*���<�1<���j�P�7[贇`+�����7�|�KU�����ç���j�J���bn�'�è������P�3�	$	*6zQ��l��w�B�B�	�%���G����g�"����K%��F�n/�Vk$�Zh�l���~�Rqp( 7�|㙳;���h6xo���6��QdϞ�ٳ��b�����~��&<0g����M�}�E��*,�͗�����T��
D�Ytڛ�|�О?�w/����������-��N�m�=�F?X���/�>q�n��}q��6s�[`�e�T��T6Q��ա:�yb�M��w�Q涒�%g �W�A���/���^;p1 �vL,��$XQR�V�I�����XK�y�ah
�H��C��՝8�csRޓ��G����г')��>�E/��^�eBH���Y(�^r�E��L_g#����P����6��Fk�v9��e�DT����θ��%b�{=���{B�uQ�`'�V��RU��!�魈 Z��ǫ4c.�bW��^�']Ml<�9�o�-͎lQc�!xLɹ/��޼j׮_��ft�`�Kң�02����Ib7
*�S������vrx׮_�h��7쏿�W��1��:�S�J��VX(�B�B��V/X��qa�V"�^����jf�̬�3�я���my�g'�(�"�~�E[�!~9<Jo�?|d��y*�ٿ1�bR1�-�rx�Tf�T��������}^#�Y��L�V�G01�b������5�-��H|lY����kFQ��i!N�n`K��.��^.ō x''�)���D"KB[����v�=\�֠0�ďJ5$�}�&W�V����qKȋ�WĹ_WwSV�n�uT���_��olII~;��UkB��5q{)���z^�z�k_�`���?���t5��<b������Ȉ L���{�g��[c�g0Z��x��n�8��_6���%��%�ڀ-�:��-�;��/�R�Qh�,?�B:�n�fۛ���,|��Z�1�����m�j�����s�n���&��+�/��* ���`��ߗQ����SU��f�K�!�W�D����Ρ�e�I >��"�ܯ�/��8L�*ؙ�K��������T\Sq��ͭ�x�����Joon�GAy���84~�����?����8�t��ͤ�U+�5�@M o7z&@�(������n���}��=z����-�|�/&s`1x+�g��6�*���iK$}�vZTZ$	NHsWe��:�ټ�sӳu��,�#����'��T�\����#T�@ty�7���(���.F��a�Pc�NN\2l{G�����I���~��9 �%%��
��az�Q_���˛tА p� �* �5��@�$we��T<	��{b����Q��i:�l9�l5�4�oK�uH�Tě8��=6����ץ �����܃{������Z������+/�|޷������+v�ʶ��7�<A/����CW��Rby�ąS��XF��������/R+�m��"Me����[v�O��ɨ��v�`I2���~	��W�"�zz]���F/Vu�Yb�,���G��u�Z�Jƣ�MP��6�3\��jKV��P�6a[�@]I�FU�r��*2�By���տa�9�"B���1[Y N}��(#wb+�P�`�^.0;����(�����e�    IDAT8�V�,�"˚�O�at���9��iD�@���gl=A-�E�N��Q��P���	�`�m�l����Ƶ7�|��>($��	�Kv4���`*� ���n��l:a��e� x�Ɛ]
6����8��
��\�o5O��Bu(�!�:*�s��V��6������ll�~`�:�M�N��[�6um��L����H���G�d�M��:k��� ��,������N��]�'*m��Z�_T��LE*-7h�����@��sx�,6!s����w��IZm|3�=���������������ST�:A
�ҥKlggW�������&CU^2���oݲ��﹬�lŨz`6�-I��ݰ<iZ��q�58��@�rq��4��[��uͼ��o�D&b��D�&N�����C?�~ �ϕ�D��`U ��/Bw�9e��A�<�"\����d�0�A�	�q�qxp_�_���za]�2r5��<���}���H?�Dj��o:! �\.=Q��3{���Dq��a|���W�)���p<r	I�����INt@�2�u�`�q](��A��J%�}� 6@ɿz���r5�HRH�ѯ��f>�����˱z��t`��P$� sG̒��r7nܰ�W_*��L��S�"��U������P)rxVo����'����'�����zm���[g_��|ް)����&�+�ǰ�C���(%9P�*����ZU�q%�Q���۰ái����
R
-�-pȚZ��2�<W ��OrØ�dH�l9�sUp�q��Y�Q���g���D�-�-Y�浔��`��n�G�c�T?�odYc���5(� Zͦ�����Ǹ��'�L-��"��%[�4<_)�'��ޕF��s�&I�ѵ���MErL�f��%I���.���%��	�����[=�^E�U~.�{�����Ұf����}٨���	�*׌&2D1Ё��Ƈo��%�lo�����j��@F�<�s�ݪ��/�Z\Y��Jeh���r�����'4�]�b8�ق��t,H6)4�D��ק�(d�m�4+r����ҙu��̤!<�/l<�[	vZ��b�J�ة5��q�����nY�ճ��M&�����_���yO�l�e0O`��q=**�J�̢ -]-��{�r��?�3���{��Ⱦ�d�Ξ۶�rd�[mU�$��e�{牌2ƤJjp[������Φ]�pN#@lbƅ��`��]��������}d�>v�~ym��}�6I6-)v�LƷ�����2�u���a�L#��ҡ��rY����@J�`��C3jY�^-fF��"���e�@a�!4G4��_dL�l^w�i��׉��r�-��ĕuf@�w
s�u�iĈ 0$� �\���h��쎏�l0�#�L�Cz�Ԉ�d�{��{-�P��>B����D 񶂣T�y���G�J�gX��^gF$�� �_W�NbA _F 6S�U靺r�ˋ I���T��IJ�eɚ"j1����X�6˙#瞎CoiG�wn�� �K���mwT��FV"p�/�̣.g���?�����C���v�e��ݻ�����+v嵞}��߳w�m�Lc7AymnE�~�(2_�Z�b���YͭE�V�kb�&�?/k��ߵ�~�Ҥ�=��PS����	B���BM�����C�$�x�Ցk�A���Z���:�BL<���tlc�e]��y])|	>��b
"����$A�NILy����U���z�����Q�4�|�kEBNU�jy�p����g��b���k�f%_���[�0��(ơD&�����'D�%a�7<�U�k�x�Ǔ�޶��lA\Ԣ���w�~����H��J����F���&�6_L�]�����Ǝ��h?#4T������S��Ð�6�T����"K�E�M@-�v�Z��M�G6���]��C����3;�uxb��P�C�0/�-EI�!�h��X��é=�;��޳��?>a�����>R`I����d2b��e��b%�ƫ��k��b�L���s��g�j3�<U/y�����ⱂm��t�-������ �`^�↍�bn{6L�~l���pg�
�\;V,n�:�{R�b���a�3�U �Md"^��+Eyh��
�ed���$���ѧ���2u�-x��zCd`{�qr�`1����o	�5���:����sU�I�;�
�%�#}S!0�ɝH6�Fmze͆����NX�#H/4�ZW�^���0k?@�1Kƞ�� ��Ҡ� �G	� �g�l�h�7:�p��W� ����\�D�q�g.��,��,�S��*�!4��c�͹�H��g���`�ҩ����.c6�7�<�Sx�1�M�bckS�X�ޜ;G����=��\8L��>e)W����]����Դo}�;��.�Ŏ�Ǿ�4C\`��T�H|�dV�fV���Jj�d�џn�%&r�U�j�c�����=;�t,M:6�F�=̽���M �D���W��>��vd���S�E=G�&���aݩ�;�g����1��h�/*B���Bb'Ғ4�Z�*R�n1ⷷ�w�ێ�v�>V;!���:y/z� 1�Ai��P��������%k�2m&��}�P	�K���(i�	�?>
�{�+�Vα��-�-1�� ��>��f��{D����~z���__��_�?~e�\�Ç����`�?�'���P'�T}�����>J���F,})':%$� `�;K��؋�c�"fY����h��'��]dTa!z_1�4 ǘM6Z�^����+�Z���X�������/�n0�](lI^ck�{��ר�ы=�(�0��@�Ǻ������XAI�{��
0 ��l0��Pb3I�W�Ԫ�ҭn�zu���{�W�������3v˜�bZ�U��ސ�
U�U�%�C�V���~���=~�!4�ZV@9ٲ��|ݶl�"�%)����1����#�T	�y���`~�4/t�T�hS��E�X蟒�/pb|�|_��������N�䕠��*|��n�k �0�C�3]����Z, a�H�jv\��C��HO�?�b�!�����T�F���Mܝ�_�L�~F�T�̣j��`���y��W��Ș�.�}#8z%��#p�Q^�0��$�t�.X�0vL�@B@EK� ����[i�`+/��q�RkP��
��5Be�����FW	�ܯB����x�X���g��fQ	,|N�U�������kg/5�/��o��ܣ���A�l�I	�E[�4h��`�mf�Rn�v�z-k��Vn6����~��c�7,/y�%c��H��sD�g�A��y�ǕL�,�cn̮$0������XDvm<�i���Q�����b�]D��&�J%T�fl	������y07)��O��ԫvꜼ�3[H�A�$ [׌w�b^G�!�p1��Q���� ē��$[�j�ŭ$�xZ�G��=� #
�[�s�y_��֞T���E�r�7�V�H��`�=�Rۧo���y�?����lA��\&B#�(�r,%�ܸZ!t=a˶r����m����?��þ���k�"���4�4W�YX��U*.m�?�A��5�;�۴+�q�i�x���`lK 7���6�,O��(�/)( J�ϊ��ha�=�{���Eǜ0�N�3`���l�� ���h��m�Fx�lf`���ARp+�}a|��(��ٞ]��+?��xa��e{�6�%TJ!ؖK�ol�$��$|Z�<��ѡ��k�:6�.�������]�!�⤂l�%2l���4{����d���fϝ�Y���gϾ���{����B�������aA����4B)�^T BM�;U�}-w�qO�Xe�GɈF`g�@a.(�4�B��}X�-�!g$�
�z�I�y&V�Ι3�#
�s��VWBL�R�pJ�u�ݫXaB.'�q�as�H9Mmx�w([�G;i�9OV�����Կ'��!��鷡|��^�}���a`�15Q�	�|�E�0`h��H2JZr�`+)r}Y�������:t�Z�^�u)Hai���^q�{� N�.8��r"��IZbR�۽�(Z�ط�߹h�^�)�޻��٬fh�g,�[�$r�F��
�i��.X���R>U��L#��v�J�������}�zb#C��y�����j���p&��菷,
r���l��`�~DYJu={�턙Z'/e�&Be�r�+��\V ���M���Rϑe�хoX���Z�2b��`hds��f(��}�zJ�p�
,d�b9!��力u#�s�ڋb% O��#V�Jf?PT����1;[�b����/�D�$:�`bt��p�k;b�ly)E�]�Q=Z[�l�OT��\�B�mw?������7��<������s������zbWds%S��h@v(O~�[��H^��?�� ْlI�(��p�n��f�ǚo����|���s;~i�/P�U��=����~��k����KA�q��[�{f5��F���#�6��l
�(Q�$ifv�FE�x�=���e�A�k�62����aw0��*�`L��E'�L]J?�u��y�jLl�k���e�c�z�j/=�e7n\��`d��޷�,�ě٠?��틉��0G���p�O/�E�;
��n;y��=�� �dq�-�F��G����`�𣳑E��̝��6Z�h�zޞ~�����ު߰{�����Gn.�	Y6��]��gW�\�j��|�-�?�:=�v���Éݿ���~x��~R���\�q|>�2�=����8��\�`f��N�����V�PE�S�/wz���$�x��K�A���\�]���#Q#H�j�ReF���墔��sA�X�4Q.�Uo�c�hR�� @�S�0Ǒf�?��\sg��5���8�֥*�r��!J�P�8����bBw')�H���! �g��
�]�+�dҸ�٩>���Qu�3QA�k6��9ZC`,l���ji�y�I���࢛���w�0	#=�%vrKrq��E*�C��q�	{�[����s�
Q��2ש�v蒔�&����C̵m��6�ۋ/]�'�ޱ��ڷ��w�� �mv)����Է�f�V��6�Y�����ʹ�U�k֪����V���џ�>��~�V�-����#㾤}�	�5\
���<A��%�����Fp%㞱�=Y�
[PI��W��t}k���}�~D4k��t��vw��������W��[̵go)iJs�<���%��<�s6<ɞ���(��i�_�u�Lу� ��Gos�8K��yz�l3%��b'���M'�C\����������I�1���xo�ZH+9���zS�-�wjh#�㥍�&�����Z�W�%�h;]�+�yY������%� �2���׹ϩ��k�T�la�3�^.sѦ3��R'rP�0RPJL�d�<��%��M�wvd'G��_-칛���s5�v�a��X�(�'�r���ߛ�N��ÞCp?V���������V(���9����u�r�S�OS�x&�:�P�,�|�:l�Ԓ�AB	�>�R���F�`��S�Q���3O?f����Ù�m=mw���{l�Y������r�R��vw�T������v���z�������{��J�{��:�N2M	y��+awR��m08�ٸ%Gj��f���4m$�W���gk=	z8T��� <��5�fnV��\W*C	~��9�g�_'<Iu2��h`�w�7�z�Jh0�i0\KF*�W����aμ�z���}FP�=��5j5��L�yThX����ɸ�>_��U$�G�W^�WB�+�=��
�I0r��F5�.v����/����J����wɓ\��ֱ���P&�*������� �=�%&3ȼ��p)�)�w��UY�]��J�YYUY29@fs�,�������&B����Y�>�n]�Ǟl�_�o���f
����b�\�D���#U��e�\�[�<�z�@��F�=�W��4����P��5��2Ke�HQ$�p�b}�(���֮����}K�G[�4Y�I�E(W�h�w������($ԻLm�h#��m@eI��9��-�^W�%�l�>/p�Kz�.���e0zr�Dh{�(���4�d��`����T�jMb����!Vu���5$bn�'�YflK87y�8':��s�IG\Z�ް��&c�R\��agk�8�Hd���,?Fީ�?x�����8�9�B{�G���dr���Ei�? w��P3dzv����N؍���!9x?rR�3�(�h;4g�}\zN�2�'��� �z��N��:>���}I~���孱|r�>mu��Y<�@����\ۙ`�"��Z"L�K�pj�q��� ��?z�Y6|��0�!���ޠ��
ST��|�T�J ��+��Cw��
ykԋ���={��E������ݹ��n�y �r�b���}]ӌ����T�����n��?Y�MvvұG����e�����Ӵ\q�
���lK/mz��Ҷ���[ڸ����Z>;�j9#r��N�]x���^,`Q�C�q�l���3�J�XC�A3A���X�;Q�͹��7�8JpUrrs����d��?C��W'�`�!������<���_D�af;3S��y�#���䙤�D�`+Ͻ���mR�A@����؅�]�z�����ݮ#��j�����\��j}��SHT��d��"�$ssAk|�x9.�l��j� ���e��Τ]�C�26�5�>�B����b,:$�ϻB���(�������˗܊.��`�$r�z�wY:9=�}���T���b�dv��m{���v���}�߶�w �ԭ��2>7�ȏ-�b[S��FTAТ+�䐉��m�7�$��J=o��=;l���oܳ���`�80�d0q�Z�T����Κ|�N
�毒̹����:�w��s�s�I�\b"�H�:Q�^)�t蔽0��	p�
6�?HĻn�m�^w;���`�>P+&���5((���!��珱����}~�d4�iG�3����T�En���?�\[��F�ux�{�$�ѣ��)$'%�$�>��ﯜs�x[9�7B&��9۝Z��+�^x6�I���1��B�m�������o�Rd.�ӝY�3��<2s��d�Bb�9�J
6���~.�6�1{y���xZ�;�!�2h�~���"D�J��eb�|6��{�cW.ڭ���N�yݩ�{t|bC��H��C+�D�>�?�Y�D�K8��ЫE7f�ݫi�p��������N-W�h�x
d�>M�c�%�8�a�!���y���s{I�0͢j�����o^���/X�s��_._��۷�$غF,U)���7#7�5�"�e�XY1�?2
R��������v|r�Uؔ�ٖ�,�ٱŪn��'�*�����f���V�����׊V�#ߖ�:D�\A*�S>_�rի]Դ3e鵻�;c+0J]�	B\o��Hd��H��A��$�v���������9'�`3����!����^n֪���@�s����{�~@��Ęa���G�ZS�sDߘ�.�T�������n�3&P]�xI�-��1 >��Ր:���Y���~����F	���cu�d2~�9$������>>��>�iJ��a_����JCY��hb�j]�?D�C*ps{��O�g>�II9�7-bL^��ؓZ.zZ'�'12HJj�������G��'_}��.�+_������a�	ab��$e���i!k�:�^lk��mղ֬�k/ɜ��U�B�a������k'ݪ��UL�%��ytL r��ry�ۍ�5��=�_��\��d���Ԭ+���6D��绯�5b�Z��TeZ3�iO���O00��`���xe�Ιu%Jk(#B����,JW�2O#>J*��.3��6���U�äN0S�M�FɖRo�\����'���\26Ic>⌤y{΄��y_�_������DX��/Ir�@�x��ʺf���y�sϫU�j���3�����0���׽�6��dP���Z��ffa�RيU)�=�����7�3#��)3�@EI��bӠ7T��3��*�s����g�����ՌtZO�އ�ۓׯ��/ܴ�bdg�Gd�    IDAT:�����c��ﰸ���`k�{>U��՚ɜ�+Ws�����{vt<���]�B�"1�q�2˂K0.&�Q{Q�����*Y±����(�i$���瞹jOݼf�Ή�F�&�� ut|*�*�O���p7�.��=��������N�G�ְ��C{���t�)xi/��G]�\v�t���2����Y1?�|v =���̊���a��2H	I*�ԃ��>A�x�jT��B4:��K@K����"��H���x	��刯W*u$ -%/nc�z�e'A����d�LU��F���C>��^U��H��^ӡ���a�MA{���CBA-'I�1ZCB�u"��~��oi�rU�'(��T�d��u� �Cu)z�\d�Թ�s˺���Z'RL�TA@�k!4���W69�}o�:Id`*������q/���O?i�z�%k�+��`c�#b�Yh�l�`K��{ i�/��K�v�&	:g؋/_��K�P�.�Jf9c �@��e`��L��Zw���k�0rye�RN0r�Y�j� �(R�}�Ck
��|N�VN^\7+
Ff?�y6�m���V���=['��$�r�7I�?(9��x�� '0�����ʄ�K5ҷ�>p�[���B޴�HTY_)�r���GPM� ~޿��f��~�"�v �%���j�@
��P����r:�b��眓�*��h��	T�+���m^�5A
O�������L�A�լm�Ӯ��V+l�����O���3�L�g#�ϡ��EW�{����٠������,D,�E�����*���ŭ$9�,9��k�����Y	G�?�N$��6nF@�re^�TrV�ߚ_Z���>x�-�x�i�<q����:]--�ݳ���U2�'�?�>"��J��e7"�mWȔ�6Y�^����m��՛[&�P�;�����{���P��T�Y�gs! ���bd�[���^��^�i�.�0Զ����*�KzN�.�p��E{��v�+Z�n��|�C������<�w�}w]-E��L�r�=����e9�ҝ�9�ul>=�lvh��Y}�W`BP�4�f:(��$Xj��7Pd�l('��SV��*}�X�'�xV6� e�i���G0�����D�N�Ƽ�4v#7��S�w33���\��g4�ﱳ����s��Чù�9�F"e1Id�a̡�ߩP�9�|ͧV+�TY������M��R
�i�P,XPdR�xW�$'�W��D{`�.i��0Z0>���-�H�4��b����zP\��u������S7�O~�%!+>҃���3�+p
��0}��dȞ,�������}��ߴ��I^<�"x"�`�����
9�T*�u��V)8Ajk�j�ZΖ��u�����;A����F�T�gTqy�jR:S�H�W8a9�օ'"Y���5%؆*�fo6T�"���|�%��'�qF�%�#��bQޗ�'rY�t�
�YPͲ�"Qd,(*K�����;��R�-e.^��V�N��U�D�+��l����N�B�-���E΋���@���p�+��C�&����!By��Y��ǰ���S�mV�
��`%oUj$9,Q~a֟�l�������A�U����GK����@=[.nΖ��΂�!���Ol��W:I�SPN=ي�����x@4RlI�[X�E/�v��U�̤Vl2��K�|zv&z���k�e&}��7pX��kY�jٜe�-�n���Z�B�0�7�|��{��Fӂ-�5@���j�or������bkE��h�z�p[E����g���?���{gvxԶѠb������2yl��,ɽ�m�l	�R�� <4Z^n8%{x���bs�W"3l���`kp*�Z�F�#��ZY��w5/�5Ո�{̀���Os��B��;�83	���@@R]Jڿꇖ}�_�;�00\T��*8LRE��-��e]�=�V�{/h]U�����O���O�!��&�zK�-�]d�wy�( o�ê�W���#0&@tҔ��;�Y�\��c�G�T0�QD?� �=�L��&�q�z恨�A(����O D����g-*;,��q�>��� ?3�X.���瞲�|�Sb��:�ږ�U,93�$3$l}mx��*k>�'��!��׾m/޺b��/��-��9ۺ�'$�Ɏ� �Α�:Ѝ�����F�E�ʖ9[����?��?z�`�-s�h���60�m΍#��_�`,d	��o�����(�#���x0r�F(GZ�QHzB&F�ؠ�DD��q�=ͭ�7	W;;F�Xw���Re��UYs]��=Qt�T%̜'[P%\�Ua�7p�x 7�6G4Bl�q�'I�n���8��M�����b�Ϣ�K���
`��3�9�����+!�x����K��y����:ؖ��^y��͏Aj��_99<�7�v.����:+���[�p:�E��C4�7w����9�<>�D�ٿP�Nլ̭ɤ��M�gd�<	X�Q-��v�vje�N����D�g�H#T#�nGR�����c ��=k�l���p�h{HN���]��Ձg�o�����Ƈ�X�$�?��l�	&�S!!S��
~������CPf�l��sl�?e�~ˎ�{6��ûG��%W��C��ꎲ�ݝ���\���6#��&iiNEҴ����w��@��
��<r��+*�G�Q��xpd;;{��ǥړ�����	"�\�C����e��8�@�>��$]�w�U��K�P��@��^�M�T�|�O�h�~R�P���=�}3*UHH�&HMϭ�_��H�0z� 3_��H��MTD���UQ����;��q�9��!)�g�`�� H�� ����Dz���$�B�ѻ�Z���G��c�)*� j�=��H�B$�HrK,8cya-���	<�#���g��������5P�"�^҂��6S��(���d>���q��M�6�ܱO~�q�x�d�m��'iD�.�ٱ��� �����z��f�*�5�f��Y)�dcٶ�kb#/sy����lǋ�z����� �$[F�$.�DY(Δt����+Hg�ܔDG6adB�hs]s=F^Z��!�t���G���6�=C+�k��){$�/��1Ҙ8/��BV�/����R�'�ɮȞ<6��C���VhNR�ڄ�Q`��К�n��<o$�R�Ӽ{HW�:����8�I3>���i�s`/X9_�w�M��"�`d���b��_y�����Z�2���>M:OlÙ����額;���L
J�EE������\�v)H��z^y����y�H�T�Y@�=6��:�+S�1��i�@N�`pz|b���JŹ��U��g,���Y������aϦӊ]ػl;��m5r����/�o?��|�'�XTl0^Ʉ(B�M$�yI�k�@0����n�.Ҥ���/|�g��T��^�/��g�����Ά6����Y�;E�4_���3^�ۖ�~�b��|	x�*�˗�Z�ݳ�|���:��[vݳ-�,�%(���l�pxh�yך[Y{�OY1�����T9t�9��$X��<�?،.l�p�y��`˦�p�U�a���$\v/Gp"��<.`&e勥��IG���B�F�uD*��vD�����xD����\bL&B��z�N�
(4޻��Qlr�&`_HC�QQ�j}F�M5"�->gf����d����� �b�,c��ق ��� �J)���d���I{��2���c���N�e����u6f�\L��@��3����?c�ۍT�;�N�&�R�r�����m�'f���=!���Znvd���M۾��?�ӿ�`;��h��X�1��1�t�W�1�Қ������YcܼR,Xs��m�2Œ=:���^�m�іͬ�e�O`�'Q���l�wR�D14�z��?��
�DFk���FN�6X��F�5q
t��JF�M�_�iU��³V�@�⚞��4��VCҤV.FJ�D$q��uOq�3潎��%g���V�c��Ո#��7�7�m�OEZ��۰	'��P2Ȥ����EG H�G�Ȑ�Re+"W���-�����S��O�֛�?ǯ_(���l����h�~u������uzx�.��΀(�g���WbJ�:��?P�{u���$/O��F0ܬ9����G�dZ<���*��|h���(8��0�,���Y��T�����.^��+/>��Y�T��m?|���pܱ��+�,m{+o{�V,9	���{���m6/Zo8�r�d���&Ӿ�>9�=ࢃ�g�FV?�WK���j����l��-f�v������i�}m!����ڝ� Q��}�	׮^���-�taWD(Fo���AW�\[��i۾�Ϳ�~�oFl�-+�Ի"�p8�g=���2}���S{���ը���#m��ɘ���p��7�`9'�8d�^�<px�J/�: &����zpR��8���
j���x
	���S��Y��6�����lyX�av>�a�����uR?�{�^�a�$���"jC>CK0`�+UA�$��u��咍�r[��7���u��σx����%�K��""Zp^���4R�a�DyŢ'-��l�Ȑa�tڶ��a��I�� 	����5"ؾ��O��VC���a-x��{0e�@�^���E->'{���<󬝝<����~���[cwi�����5�K��X�~����H`��} ��3xn͆��5�ڌ�3�Ƞ�+U[�l�k\b��G���jQ2��E�umm�����h;�ƥ@��	��rYc8�ra(*vn��"�7��L�)��>l�o'�ƚӍ����u7� A `l��^�Yߥ�E9����V"��׮�b){k3z���)�&��A����?�C�9��B�p��G�"%>�?�?�)֪
�Td��$�x|���p���^��-�E-���O��"0�ǋ �`{�ï�'�_����j-����ye�EV"ܯL��<��[���"娠����dt�SC%���d>�)
7S<pS���:����4�d4�j)g���F#)0y�+/]�$f�ȡ=���}����dֵz�i����޷�cf�v�RnZ����5�6��dC����Gv��r�X�0���y�ơ�@;N79US���һXT���0�p	>� ,X&3�W^�b��+��O�yώN��lܰ;w���*؆v/=&�N��t���*����D׶R�k�0c����X�!#��;V,�X�@��Nkn�'V)S}���37�ۅ�;vvr�ୂ�E�����v�+.X�J�:�J�
�C@���N��O=Rشk�X2Q�n���E6.�.Vl>��~�bS��@Y��J�иKb�9Ni��gF�H�F��Z=�N��8Tc,	�
G3����x�)�H��`�.l�6�Wū*6��RHj��J0��BA��=f$��Db�p����v���<QI���.��ʥ��n���c��'� ͈�3�<c/���Z.�J���O����Ѡo�N[���Lz���^<��svzxǦ����_�e��?�������Z�L(�e�x�z� D�f[y�UWV.έZXY���E����n�XmhΖ�v8۳e~��٬`X�&�ک��.�O��u��qi� g*k��Q2�� �ڮ��		��Y$=T����O��j���^[������XFI��ֶ�Iz�h$S�p>�,�R1�	Y�gރ���8�$y�����}�j
R����M
(����!�#�D���xl�E �Hh��8|��P�K�ت#T$B�}JX�XQ�w���s�{�mۮ����'���d�:w�{��_�����E���Ӷuzl���&Y�3�M%P!�KzםU�bh�B�uiC
^�X��df��26� ���M����1�Q�,�Z�p�����8����q�A|1]J"ϖ3��*Y������b�;x���������};>���$�V(Y�^��+lK\Tx��p���b&�F|��Y'����C��Hp	)ewS�m�L.`�bab�ܺ`_���ۻܳ{�Vo>f���aK}%Rz�X,h�h�ٻxUd�~�1���&l�m{�w�o��r�=b���lZ��4����ss U9�M���涻]��;>������h(�P�Rj1fX���(6B�A�	S��n��k4h9Ӻ!��=s=#����\�GE����*V��TEG�{ ^���R�Y��1_;2��z�:\R*�u��601��4�7��8�^>�*PQRy@���� @y��J7 Ii\J9��v��"�[:�J�}>l��S.^�믠�;�.�t�X��Z�"q��3�}��:���Ǔ������3� �I�1���!�8��14ر:XAR�l�I���=c�ᙵ�~j��³v����?���}on�p=h����Bx��Hg��E��ӊ�V�2NE6��VU���l����Go�`�k�eY~�c��Y� �eqFH�0G����u��s4���@=Ҥ	�+�=`�VYr� GU�W$*B0R0������T̎RQR�ˮ��d�~�իW����p�2�ŵ&�ܜ�� )�jZ�ީ��D1�~���j�$A*z�alA��vm������B(��dA-�X{)G��
Uh��E��^��+Hye�	�:���
.H�mc�X�FͶjuۭ5�r�ŏg�m���g��7���;��Y����'9�LQ�qat�r�'����`'`���+��`��ߛ�'n6?�8lۈ�,�߃���C	��wxHљ|e�u�WE��m�p��(Ӟ�j=�`���l��z=2:��N`iԪV�1I���p +�-cw�� x�?����Ön�N����H��_+K�4��M��k���U�n��\,_�w޹o��d���$� �ԕ+�lo��m�]����|�f��̬X*��۷���߷A������`��-_��(�j�U�V2��/�=Cv���o4j������8+;��x��?�����O� }��
Z�j$��a%��������L����w�Z��Z�>|����<V���*������POwcH_�/���!/���p��O(��6䁜�����%}.�Ъb�L�|䳽��+eEu�x�8�:mUҳ�lO��d!��㚭{�I�k�����R�Z����I�k&�D,�J���v��M��n&x����4�Rg�ReQݒ������\�#lf�x�9N�}����nڍ�.ڟ�v�ݹ�:���Ҩl��DT[���Z���3�X1���-��1g���������~��}� U��zN&P�BH��yVf���r�k�g��
4�E,\8EP��X���%��D
�$�Q������y���bһEj��Ju)��&��/_��`K'�#���;!*ؤY���s��h|m��0��H�xz�J�  �^���<6�ɑ K)0���/N�N�H
��gҾ���Y�g7=! +�O��D��qA�B�N(M"\�<Rx`R��$hA���E�ݩ6��­'?��m����m4m���eK��)z�4���J�]3�@��I/vI�q���g�����jex���CF�̩%�A杤�"#�4+�+����.�L�02X���[��סU�XV6w�^U��m�vm�t�)X)e�R��iUT{���l:�rf�W[�=$�r�J��d����!�{$�Ƥ �,V��ˬ:��/<a���/(�޾wj���}��#k��ww.b�K�_������֎2���Gm�8���Lʕ���ӷ��?��MF��8��,�+'#y:�=[����t��/��p��v��%��`�a��Y/��"�%}SH-!���ȃ�g��3����+Y�9��=	ED��6�~2R�Ҏ ��׉@���Qo+��l�>��Mx�{�^1o̨��Ɩԃy�$�ϓcp�Yt<;�8�`/'��{|��É�Z�쉨ڣ2�ʛ�3t|>���8��D��DTR������N�Q(�������|�){���P��v�u��I��n�"����
��4��X�{�����p���W����l_��w��{{�?�ш(��N.�i<�SG��t@B�RC�Ń-޸�f�bEt�wjV�V���;ڲѼ��V��le9�|��eg�?�~%q+W��m�4T\���V-0A\\�N��휏{;XU[�8%��    IDATlK�U�%�U�K�O�%1�i�PP���u���x��'jeŽ'Ъ���j���K�3�K *`БXo�I&��	n"'�=I$��oP����3%^��~�}�׈��=������O�A����m���C�w�/������������!�R��ʭ?������8���U[7��xb�mD*�ƫ[�՗	<�s�2�h�t�px!���Zmv$�Y��q�*
OGƀt�7zk�}��,ln(��Tl,$�4'��u;=����0i%d���Z��d�� >��<W��Q��� }c�]���[G6v]���,����1�p>�F�YJ�T�@��F�Ez���.:�3=��?�i���bo����'w-_ܳ�c\Z�]zI�!Q{��x��1�O����`��C0cS����{�	V�a�>t�ƪ�Kz�lRz����袸�ӿ�Y�b�sp2r�&w��M@���Nm ��F6�ڨ�7�+6�/2���|'�i�X���C�n��/��D�;���F�4���L[�fx�VP_x@ż	}yO��sw��s+�S|&���
�8f�Dx�α�-?$Aʟ�p���
e�G�4y� �1<�#I��Q��_z������ 2@Ϳ������a�J�� B���ޅ��l_}�U�t邳��: �R��x"�y���{��!	-\��=�\��O>i��[���=��{�ƞ}�kk>4;>f�-,_�ʏI�����Y	BT�����-����n����d�V��\����D�m���l'��%M(�"mW�"xl7���@�� �b�"��i.hj=[�v�^��QiCh?��B[��/�����I�zD%��iT�hl�;'�q0��p�ji�e��F2�I9�}��8��������z��H�%n��j"#�<��ZGIfQC\i*@�*dá3��>b�������{���>K�b������(9��}��RNe�%T�}Q��}�֋727m쇿�_�=�����MN�p��h`��xd�g�T�Rk��\n�ግQR�P.!Hq� ��L�������9�������b�2�;�()��.�I�Z�t.ъA�%e��<n.vQr�(����O�E�Hv�bG����C���2<@�YF�lR*�P(*�0R�p/�Вʑ^g��حtyO���~�מ��k_��~����OX�~��������߶jK�����]�v�._�*&2��p�U`b�i�n�siw�ܱ�wokJ� �̹���[)�z��1��=��9ؚ�g�"D���A�z�X���$����r�����5Â��lV�Q�������rBVW�"h+���N�Mil(��h
�M�ʂ�8�\6�\�蟁���2k��S��8\b'��97__-��ٕ�&�/�-�1l7�_��I,�H`�q��`�����*����r�rh1����>�Ip>��W/ۭ[���Wo:�PR��nL�dڳvK}�`�:�=���7�.��>�'onٕkM����5ۿC�.*آ����m.�d#�+I!�6���uIƂ�/^�+�;��y+T*
���#��bY�[��l�t�}π@�l�L��sOAJ���D��(�2��� ���a�,�y}!B�^��YP����R����g"۱��$%�	�T��	jgY�ӜF��4�`�N���c���V�y�3��E�S�T\<F���Ť�s�w$|$
��,��{64�#و ��\�כ��:�>J���Q�wmA����P>1�����*��^�ĭ'>��v�z��`t��t�R�;=���)�$��#�,� '����㹪\�@�����F0��9���S	��<�٨:$U����~tx��Y�geHh�p�NwwFq��@��[d#a.��.إ�%�L����?�N��j��1���GOփ�̚cZl�9�փ��Jy��݉G�O�����Vg�;��I���_�������3�o=f��[����B�� ���(ؒW�<����c���ޏLJ+o�����'?;[�8#T�9d��I����r��)к�'9�k�{�	�w��R�A Q|m��`��.�mT��9S��U&f��rT�#�ǡ�2�	H7`����A/�`=6!&PY�"�%�[��&�M�=�u KyT�!	���2`ۀqׯ�`<�;B����6�uV!��x�
h\�/�oSB���>:pI���f\S�����2SJ��4�! ��6�����r9���k|��k"�*XG
����H	x�p���x=�8	�O>��]�-۰��=�TӮ\�����؃;t{3�-�.�E&�R�so������lw;o[��5�̧.����+������[�T�䍖��g+�doep��ٺی��	��hp]�n�
�ĕ�bLAo;��]�����S�%��<>��TV-�'l�H����&�f�Tt�>��6�H�2yֆ\f��Ba��H�����ۙ} ��V�(��Ԏq��+\����IK��F�2놿�ِ	�u��M�@J�^��G9�"����LF��\�j�,�Q)+�
F�6�_��T������{��^ٮF�7���g�
z���E��,�\�|�]y�B�O�=�d'S�2�w�jV�����2��
���0�+��R��SE�(���)k��_b�֪e�P��T�}exP0	s�R��% 8땀K%G{֭zA����\��I��e@7@��3I::�B��#׏�K��M�b���D�K�Z�>f�����~�>i������o~���o��|��DCP��U?5��z�j;;{v��'4������Ml�����Oj�����slK�dZ����-�@Jc[NJq�6�g�n���M���g2�ؠ��4����ͪ�*A7ؾ��ϿR�!�,xe�i|���L�}Y��&6n(&�(�g��^Id�4���T#�J΀�O$i/'���^���d�W��*����ϣG����g�`{�5Hh�־�ㄈDB���Ä?#o���C�:��N������
iI��E���nؕ+W�`v��uL�tq��0��!G�%�!�$�Ik	~��]�ݭ��zwl�]o����P�*��uK,�at��F�,��
�%�8+�g�v�bE�{������,�.^�U϶�Y��?~`m�%2p���*ۜ��ng?���F��+���wiu�|G0DmGU���x�$^�� �|�S$J�����`��ኄ�Q�d�a]��T�,�����L�Tek�y���k����\��n��:z��z�Ȑ��l#*�H�z�N����y�D��G�k���h�Jv$� ��H	��;�oL�wh#'���Z�-0r�\��[$��>�`��<�YY��q�h�+Z�T�ח�5�lג� ��fC���Rd��d��H�p
��X3�s]єI�&t�r!��?�Q�H֭�9բ#��,D@�g+���y��m4�Eh �oѦ���j[V)"������w߳^�c�{M��Se��鰣��N�W�Ju$w�dF@�;����R�7	t�hE�~�7^�/��/����kv������Ö�ޣ!���1S�L��;�,�a2��z�J?�ʒEL�}��m���fX]�g��0V���+�))��JvX`��Ѭ�#7���=��&����L�f0��Q�� rN�ʋ����}S{bЯ��$��	G��4��0|�����9��Q�-�s^����Z��G
X��So��a���u�%�?>O�u �0և���g=gl��?�É�_�Pr����q����&�e�!8�A�;)�	����<	�3ͬnb�ƾ�^smw������U-����̴r8���eL({ѻ6�[��X����d_���;���۬�+Y��h]�m�|Q��°�(k����k�V��,�l�[-eD�wi������62�-0r�l#ز^8�Q_�0lS 	IN�(8a�t��DB�� �)9�0Q�����f�(78�Q�����$����n��A����U!�6`��s�
|��*8۵	A 9i+إћh��gդB�L���#�^���B$0��:r",_�o��#��ZF9J�<��qŉQ�ne�A*`d�Sm<z��[T�?Q>h����Z�;�VظE�v�vrJO��z���"�����n��X��K��aF6�t:��l"d��X���+"��Q`����Y��u�Zp�N'�nW\a�s�q"vc�?tj�*g�BM
8�h��2u�R���ۥ�<zt,����KV)׭���E�Df����l�4�Ch�)�������a$������^��L#�����������Z3+V.���-Ic* CH@x!O�v���6간3���Q���ټo������?���̴���tf�z�Ǘ�H�eNX�sl�|�GHE:���O��>Ġ$��_6�*�oI�8�Q[h�:r}���7k@M1��g��9�'^�����Q�T��Cʑ�'#�zP�U;st��Հ�t l@���UU��
���7�r���D�bIT2�^���U�f������A��҈�)�x%���60�g���j���.;�c�E�y��^�Y��U��y)IAлpyϫe�h�}�N�NG�����ؤ9�JX�g�wl4<���}��+��K���}��S[�M9�2�ĥ(I
��J��=��Z^X����?x�l���U�M�s�eo���F�f�-����}fl4�k^����,[�3�7@Z�i�FmͰ�Q�W=�#�>�ʍ��Fף���[19����]��Q�V�� u:�����(=�X�u"���S�ae�ceD��O��c=�\�
Ɠ�Wṃ�<J3����zžY��	78qFFu�8^�Ϧ�5�B�(��)��Q�y��(ʹ�b$�^c�� ��a��\�~�02�}�ot��,��bg���;>G�������"0.�L�, �	Y�o~W�X�׳��Ve�e�6�S�!�<���sF&s�􇏎��+Za�J�����g#�d���oc���F�x����|$դRaa�[%�~�f�B��ΔM�껖ɢ�۷ã-`���t� *iA㈓T^�������p�멪o��CD�L�LX���;/�o��?����w�����s�P0=�+���$� ��{A��^kj�˞�Ѩ��q���~�އ��9]�j���)��|<�2��$T���%��d��R2b0��ϗ���on�8hT�=�e�p���ܵՆ��:P���+`�Ș7�r�0C�{��}�zM�Б��s7�1A��"��{V�K#k�L
r�=�z���F�^UG��A�P:̸�
"���A&*��ێJ_�-cA����h����#~-��&�4Sc��Z�6�%����7n��������!�	ctz=�Zp�l��O��$&�._�բg����ŗ�٧>������}�?�ˈ`:AH��Dv1��"�e3V�Q�ac8�Ra�Q z���V�y������FF�b�k؈���(�ȠPH��%�Xfm��ו`J�"��_Eb
r��õ�FKDgEJ�6!�8�)Ur�9��m��9����IIP&'�To4^�F %���TǺV�9[F!C�����s�ƺu$$�?�����0��7�Xk�}�3�XS�Ұ�"��ux|����^�����y3��T�I������`�9��W�ã��{��4���7�v���iuu�o5��Rv�voر�l��2�f��y2<h�>8��a�s 㱬��)N���l3r���Z\�:f�3k�;��-Z~���0�m��K�Q]W�T�3���c97�H糡��Y{��5��W�F���%�ە�/ٽ����P�V0[6�C���r䉓 `�q����ɉ�N��5K��`bvS�󂫎�W�����oپ���4�3_����퍍�"�7�O�V����v��%�5��k咕�%��;�l��4j?x���B�Eչ\��`�'��-\e��RI�%�Y����m"��W�-k2���D��1	�c^6��f;�w�ԝ�����w�ff�բ��Kso��(-��1�U��{��\��ѯ�k�y?�Y�a��D��B2�^n�A&��"��w#�����!?�	Iǵ��C���@���`=���Q�ǡHG����E<7�(D-���^��]��$ؒ@��#'H.j��HRСF�+ނx��ǭT����[�����?�˯۷�u��H����l��U��b~���G����WV֬a�9�Jɬ\Z�ҩՋ
��b�Gb#G����`��y���{���6� ޻���WC�=��#=N0���A�
GpX�|��պ/�:Qe�y�G��Lĥ�ϱ�&��uD��{�[�K�/U�!�ļ *�g����\ģ���.)�${3�r��{W0sI�����:��5����N�^Y�I�;�E���6ׄ��-9�ە��n=}%������`�:��[�e�� �L���,�Js�+�<<��pj�,�U�%˗���mnC[,GR&���V)l2���i�n��7��5�L�&8W��T��(;(f_�9��FîF��*s����9�H�%�2���5
@
z����.�ј�/m0�`����g��Y��O�!�+����b���`_']Z�/��ac��S�nf|2S_���������_�o~���o�e��>8�Vg�`�C�er�Z���.J&�B��R�R���ٱ��m�5궿�o��޷����#R�����wEbZ%��P��N����Б�s@��ҁ�س1�ϴi�*H�Q��I�#�eH>4;�������p2�+ض��R�oR��+�~�s���A(i�F`T��F9>l���DB�M��_M=ڀ�";"�D��DD�)X��)��рK���$'���' ���� =���3F�/��	���$�����.�H������]�7~�OFV��NT=�F�����ao1�R\X��={�ً��7������{�޷�aӉ�.3T�3+P8�kr�( q��iT�l��i�`[�l��#O��l�o�fp1�)MM0c{n�N:�\w�	k@3�)�ֵM���$���,jT�Z)IO����9������]��V�`ez�\ͦڛ<?A�X�H�J+Y	O�2&�����ґ���KK�I5��H����Er%�֫'���/�$�������������	�o����Q%�'�l�hg���S%�H&��rTbmla#k��<�����l?~����[���A�4)�h���-�9+�J�-���<9l[�����=}6�p�X���Ҳ�ѠC�9Z������f24�Jեls���y�Q��� �1F�SI4.�VdF�p )ʵD�2���Z����z_�&�Ž=�T����ӴF%�q愻��G�|'�j��h��߼6�FHc:S@�X�a�h!�"�h�����%���G��/����_���?�Y��k�{v��F���M)恷�H&�2�D�-��v�:�n�k���F0��۽����xBSTo���є�6��H�'A�Q��ro�G��؜mȹ��)����z6י��s`	�\xo5L"h�&1�5��^s���A�8_�0UT$*+@'���|�S�B久L�yY�W|�P�Y��#�l�F9t�(��k3	�j|z�I�%����*A�h�"Z'I��4z�:���-�'w���K����3�և_�ܢ������#y��U�"%N�B~�mr<B��F��,��lbׯ^�Bvb��=��%{���7�o���Y�p��3`޹�i%��A�K��X��|f�V��l���C���z�����:�f��Fe�lWF/�>�(�Ě��A.��R�$D��1rNx`)W�tA&,��>#Ye���+e��:�O$� Q�F�¦rL[*U��'�.���`K���fo)ˣ��g�\H*R��Y�m�!�5�u���v"�z��na0�e P*�/k?t$,q׬��^G�`@;��2����ȩgQv����vw��+W�|�*��ß��:��w�-W�N�vt�Q�)款-��Z#��6���u<�I@^��*լ�T�<d��ee������=:��Y��I�hV���
6�b��L�}yV^�kZ�Q��j(8�n    IDATn�։ժ>����=-����PV���� �����m�0H�-���#�N��2�����C`;�����P�2����;I�1G6Y��c����`_���տ��=xԵJ튵Z;:�h�`����-}�����.r
�'`k���c;:8Qe�:j�l
���f@#0���[JHHL���D2�<%}�f�މ�5�y�6Pl^�6.��u6���4�L�X$�t�Gp���G��7�B(H�\�6���Ħ%Y����8Tx\T����U-p�f��^�_P
�FFε�]T�q8�w��Z�:z�8�f5�%��p$$|�P���5+6����.ir+����ꩴ���G(��YY��̛O=�q�K����I�h�Wط=L�|n|&`}���+�,��|r`��z�n<�g��_�+{���V�^�芤=1-Y��1[ %�go��}�!��[����fѫ�j~l5g�����vY�� �1t#�iq�:0��Q"�i���ɍ��t�`�}.�]*�������F���'���W�bk)*E��$����.H�������[�"��h�f���SA��$S)�ʍ�:�m$����Jӥ#���P���Ík� *��ss��
�I/@~�I�QD�jM�Ý�r�����h�V�v�ĵǞ���i�e�s���������m��Lr�i�����ܚ{%���6�m2��0D�6�����m��.�Vo�c	xi%ڠ@�㕝vv��Igdg��ʳ\Q6~(")�M1[�������e[��<�Z��4��.\�S ���"&02Cp%��F�C%��v��{�:]#�џj�*M��0Yb�vEc����Ŋ<�FcP`2Y���h��D1��|�%�Wev˶����엿�)��_��=h[�~U~��GT��<ز�Պ��y_����+A&����&T��zvvڶ�IONE��W)d�ʕK���v�����|+�[�<�e��lÄ���k�F������O�	M���=*j~�I`��a��Q����uhs�b�5G�B���x���~����1ؚ��s[�A/z`�k�`D�8�t!&vz�>��*���B
HC�� Չ���S#U�X���!b#IQ1D�)sUo��M�!� y:��%�Į�������uϞz�i�E>nAT�x*[�m��*ZF��Ү=�����k�Y���]�����o���������ک���4��^2��Z��%� YŌ���m�kDA�V�*�bD��T�T���k?�/62���V�?$����0�����1N}�f���
7�6�sor�����ծ�ߘ����>��r"�2fw�V��������/�ҨKRR1�5��عc[��_��T��L#�	�i1����hڡ쭤D�����϶Eb=�"�F�\B�:��<�����Yμ�`���q� #�~�5�}k"�lC�"*ۭr����?���u�s���~�����/�~��o5��ǌ�Y�2���7S�u#���<(� B],[�PR��t��9�R�ʎApAt3�5i%�>��mw��O�*Tl���8�A�@e�����׊��U��p�9���kiF�,5H�?��h��A���J�cziy��R)���f6���C)d�dS��&ػL�*�<D!�Du- @gȲ�S8?���ǿd_��쯿���m�z�:ݹ��ŀ���d�d�[��.�����l>+ry:��t4�Ng`3���w�c��̃� :�8�w��t�h��9xe��d肙���,)��VT�1��X�b�1.��;�x?ڙ��0sT�����t����mR|"ea��i4!*M�%x.�^
�i�gS�BզQ;���C[�3���#ٹ�N�8�p��,k�+��
yN>��O].� 1MU� D��o�Q�=!���<�4) QY:k�Rkፔ,�E�fl��T����*?*�p�}�'Hm1����O
��]*&�ܳG��s��q_�R���d.��eWC;x���?�m�������{V,\�^?�ZH�I����3�V���Z]Z!?�62$*��v�V����;:IԂ�m��kc�ir@��g�<�j��Q�=�l#Iad) X��`DNWħ�{ ��gL���ֲ>#�r.K�m"ݗi�3�o��'z��#1U+g�2�-�%$`,��'���y�pY�<��
bi-�|��$�n�}�w��( &R{;�z��87���Y�����x_�F\k��1$�T'"uK�9U�0��g�U��o>q�F�q���ggo���{�����]�t�V��(k����a�@9u� �|{6���m�a˚M'=:u���g���$���U,Kv_�[4����Pҏ�m��[�<0x�#z�(ݣ5<���
���Ԅ��+wB�E�L��x���4�"IQE0��h�@���0YX��0ˠ�ڵ�d)��N&H�$�F
2皰�YJ�0ز�m��k?��h8H�#+��O��W�s���}�[g�6j��=<�^�Ì>��&x��v�1���!����h]e+��`y�͆]�>d���琏Ô��j�����d�׎`+����O�������D!CNp��:�e�6�R�IM
�MN�e���s��\�
@ٌ����`SN ��t��*%���L�@��T�D��=v�8x�3��<���<D��	I������S�Viu�3�H?v<k����	q�*���p{��@��C�:)Z-�HO6+r�� 2~oQn��'�����5�<Tf1j�k�fByM�3�|�w����	�W�������ף'$g|�H�"�⵸�E�	�C�J��}�>��v��=���忶�~w�J�+��
 \oTҀ��8��ʏ[��,X��d�jުż��b޹�T�=<����MW{6����eq#�έ���f���g����i�3��@����E�c$J	D����賒���$W�����z�iD�׉�DO�U0�	<�0cOG
����B�c] ���Ґ�G�\���k��O�v����AL{0A��(�C1J\�!Grf����k�k���@�����Vv�%���E�Vs����-���$�k�-��g�Y.[�T�f�a�J�v��c/����w�cl�����o�h6<���-��/�xV�G����Yf5�m�免�};9jiCoU)�����3�Vk`�A�f˜Fsc�m�U�H���z��Ck����y䲡�?v5]H��C��*Z�s*#�u#��� �8�s�8��*����_��Ҹ�P��b�q6W�\��Ճm;<�Y�?���D�SU˜s8�,%QA�r��M�ĺz¹'A�0c5�A�z:�rqd��{��W?y˾�7���߶�X�7֘�\�sm��m����yl�r��=��	��g,t'�����G�\��a����We�B��k������U�'k�;\vz�/r�s�9F6H>^1�!�Y�g�C�P�V�����X�/��q?ct�0���H)��R�y@� 3�af����{T���Ò��u�-��`KdM�R��]eIa*}���n��ҐL����M�Lt2��qۋ>'��WoԳL>k�^��ݦ�1�����fpp1	��B��HB�G�|�V��4��a�T]p�2uo�lC����^Y��|����s�n�V�}����K�=Z0��O�
$i�WG��kM����$�m�s�S{�����=����k�;0���'-�G���]�ŘAȬ\�$U*0���V�b���5����^�-s�-SrQ��W�0q��d9��~ib������& /��x� �\��O#���JOIS(��^(�K������I�'��r�uQ���ɏ��5EƓ�+qb߈���	����EX��I�$KΗ���4�@�BAA�N�+PQO&9��xE��/N�QB� u~�kI������:&ؒ`����JY�Iu����<��`[��[��Z���˗_���s�cl~����;ov��X�T��nX��cO���E��KV�`?��ao`���U�Z�����9�{3�s�OZm;>��lU��h*Y��֮�i�h�&*�?Aىe@���S,��RK�]��p\�;,)׎FUL6��m����[��s���gi6X�P�bDne�R�2��=z8a��h��1M�XH�3ym0D$l!c�zI���"��Fb擸�D�lj�����?���������C��l�޿�o��T#=h��ۆmo���K{
�
b��QƆ�a�j��#P���-I�E�@�� Tơ�����%4��)�P���%��{���K��[v��J�V� `7��\z����:��p�oF���V��Z�!Y����H~	�~6�&k3��xo�C�t���m�] )�e#�F3U�T|��Ҝe*J�\^���HpcA��H���kN�`+F)s��E�n��L2�B9NH�a[��tX U�s$�
��0�t��a���HGT�A.8�-©*��J"��ȈX MI������<M�G��cBӸ{���x뒂���?Q��/�l����F��C��(�o�*�Kc��EDƉ�����U��\o������[��
W-Wڵ�rn�9f�����E�H(���'�m�-#�F%���`��$�`-!Eg�W���u�g���E��	9g�I[��`�Xg�H��=�D%�5X�\74���ϽJl(|za7�`+Q�lA��
J=i�	�@p�#�V�d'�J �kWUn̴��0ж��4�D�f�T����9ZO*�:s=���� �?S��6��/_~�cl��u��[�vۗ��u�Ά9{��6�$Q�sY���{�ﴬ�yd{۰R�V.�d�>/����Yg`gݡ��]-�Zs�z��9�2w^ffR�b�#��Ř����W�V� ;T���EhC�@��cBP-�ߝHN�z1C�6$��3��.+i0ͅd:����N[s��2c8� �R;�B��T�.���:*4�����BD��esU�������w�g��~���P�j؝�G����Oa#;a�Q�r�$򘵲��RU�y�t����
�Q7�$<N���<h�!�&����D����'&�� 3'y�蕽�c��x��~�'�n[���l���`�=B��A
_��R)U�^͞�p�����6��$�F��$'�ȩ�r�A8�u���0����8<'x~-�l!�������#��vꛉ�{1�R��dCz#?��PřX��Aߡ΢'Kwb$a����H�R���U���۝���8�T1'���u�$#	υ����ɱ��?����P=l,&�p�c@��Z�/>A�Ǯl���׽�}��������G�Zn����P*�r����9"5Y��8�`����-�d�(Y��V�J՜�Je{pж��os�l�\�`a�����պ�;6%�鐗^ 2�3��EJS�y�tk�E���	���t> }��nC�+f���@ ��@T+=�`�}�>�z7���_���p@c����3';���'�g�-��`�uS�6	p���r�kz��[7ӱ�����XS��MÃ(Z�ټ#"�b� ��Ԋ�� ����>��$a
��8�`{��Տg���ty�����C	�#�W߹l���?�����
%��̩��e�����;����?cU���(��V�8Y�^wh'xa�[6]�����j�y�f���FV�-�����{eM��]�\u�;ߞ��m��`I�%KF")�iɒb$�؉d�%GS�%��$��$�%��"�T$��Hv7�M�po���p�=c��֔��~vU5#�L+h���3U���>{��^ko�jwa�-�0��ǡ6��l70�����&c��M`(l�-%�H�n֑�4�۩[�S�Q6����f��7���s�%f
ޣUPY ���V�J)2�8I�ɨ3y��*�p�a��L4[�<���W?g�l�𚝞aN߰���4�G�1[F��ӊÄT�Tl�<���G/I�x���`�C'�G�����`�v������ܗ�Q8/A�����1R�|T�a0��|=,��l�(��
!�4	m3��RO*nNs�!�3�&J>��"��`ȿ��i�ܝ�V?G&�i��?�̩��nH���d�ƈJ��O'vrT۱A�z\�R��V�
�(р��a�HXV( �	�]R�ZWG��~��P��g+�����$k� � #�%����h"Yн]{���~Xg>*o�-����`��<�����#��F�:t��/_h���/�g?��=��y�g�ۿ�o��#+��4=���b,�8�-���T�l���r%�F�ի�흖U[e�.�v��k�n<���M�w��:=�yΦK7��a�����]P(Zˉ����fzV=Ȅ@ĹE"H�\�i��V7���0�9������\)���%�)��2�'�&R�z��WC�݉�����@�@�;�w�Ԟ�ڳk���z�
��Q�1=3�&l%>���F{G���j��g�ו5���D���@OR������*yg�ZS2���e��VQe+��\��vgt���O\��zo������;y��[��Ɨ�M�v��C��ܲb������`�bæ�:���7�V+��<���LZ���{b��+�{x�����<��`R���`��m8Om>Zn9�FynO]޶g��X�&6���/+�F����"#c�s�T�R�c4�3�e����^@�B�l юnoi�aNU����c��E�=�u	X��ٴ�lyx�Ն�*�����K��{����l��G߶�.��=�?uQ��Ƕ^m��]����!i`��s��7�P�`��B1�Jl�g=�pCI��i%������+��o�G��k>������g�3���V���X �	LE�@�<�S'��7��(�,�؀&W6i+G��*�=�P�	�d�As�a���A�F���6��(�3�^l2�<�G2��cҰ�7%A�����yR礍�jZ�('�Dr%-�ԛ�{a̠*�Q/ڒBT�
0�u���Z��P��K��!�s�=��ӫ�?�ix�d�öڝU���٬r�]�{0^�����v��a�����#/�����?�_}d���Sr+6���$�0�B),��m��e�l����e�dRa��;��ݛ�6[�)ؖjU��s�s�y�tb�u3����HP �J��j2O��<�[ +1GkT�1;/��M��ֳ�\��-׸��v��zDE�sϊ�aJF��AB�x��ܚ�k���K��N��T���d-jK���D�rB��l�zX�W{O0�Ն�{2���)���ؓJO]�7�f�hPa�(V(�j*bp *e]��[
.��V��SO=w���������{���{���o��n}
���R�*[6�7�;jX6�Z�p��JQ�i��PD&��l�������?h���j(X&����ڵw������9�,6+8�o9'`ά����Ŗ=���U
�-3*ޅ=|��1���Y�q�j�4�gC�2#���,����3mJ̱!�8��E��&�dw!�!�ͨ�]�&4}b�D��a��'!z��6;�Y�lCI�^(�>�����1���}p�b��g)f��L��N��>;8/z�QQ��iĊ���2���ӻ�<���5���o|CU���)`G`����{��j3z�|&����D J�t�E�I�9܏4J �n��Q.U+3Ozb+�Sa�kK0�I�.�sUis
X=6����,T��8�X��d>6���6���<	�ʧ� O��}���������b$�Z��mD4�*�5T������{oA�M0"�')�-k���Ȭ5�%��Ǐl�$��-K�e#�u�u�i�ucm#�?�n���U�����}�+m>m��?n[2�ǳX��R�ǼW�%�F�����j��F&ؾ�ޱM�6���k����L�a#1j8�z�p���)4b��mh{����=��O,ީ'��Spq-������(�9s�D	����m�oA�M�w���gU���B�N��$$��sy(��� f���K�.�IDOJ�3�M@�Ţ'Y��'�b��D��f�     IDATȀ��8Z�J@Α��=	kK�3#���ν��)JA���\*	� ��l;[��O>���f�ч2�޼�;�����?W��HD�T�f�ʮ��e����l3�ws9�j�m���쇙��\�$��jan���X�T���{��{vwdGݜeV�!�	+2��ﲡL��fϪEg%ss	h@�Z�b��ڬj�H�̓��Ix9�!#K����d���I'�L1_����`s���;7��6��5���fK�֩!� ��|1�\�E<1�����h7�#���9�ti�>����h�[�62��wm�ܗ6y�����=�D@^���0��
S�c|()��Y9�[�R,;�����n�d���;��{���! nN��Fի�+�F�2����w�f��I��P-J#+�I��5�8,��l_7x@�c-�K����Ub�D'"ɐ2��g=_]��i��70O$�<�E��k-(l�3�~�]�;�Uީ����x�
��{���%*�D�3A�����1�4ju��ED����s�{H\��C@R�/��8��1��g��cZO8�p����"��k$(� ?�Ѱ��r<��-�3����rv���}���/ۿ���o�~c�&Y[֜��|�y/� !@޿�V�Wl6G'}n�vɶk6!�a2⒃yt��k��ڃ�]{�����-�b��cBΣ������j�dF9�|i=ǬsI}[�${Q�Eb�6��%KU����0\� <�g0�u�Hr4��=�l:[���=0�gӄ����a��~/�=�XWkQߛ ���v{��L��ua�璜�`+Y�j�ծȇU�N2�X�Ғ�.yK��>ap="�g����Q`9�8��v��ȋ��[*o��V�G/1bAU��l������]z≏�k4~(���7���0����l�X"���UsM[�/jh��m���W,�V�����li��@:0m��n����lo�c���Nz3{��#{��=:��dY�_���l@��rKk��V/ͭ^%��W�Y9���6{%�M�w{�?H�&��Ӊ>����P���󞘋� ���h�=����;�pFE�ʐ�l���'Ć��=^����3+��X�4�V}b��?�����=x8���l�'��rb��Z�Y}>�:B�@�Q���bz�ꫥBA6�� �T@��'yq�{�z��p�H��ݻ��J"6LxFT�H5F��/�|�r�'ʶO�O2�!��k�$C��͆S�JF/	�5�Ц�g��&�Uu��u���G�6��(���D��>^��x%���*?�ֽB^�a{���Kq�f.��"g!��둵oX�	{�R�^.n2�����5H�Q��� ���6٨��~��=XT��ц����y�&��
���`��fN �ܴ/d��c! x�ٓ
������?o�7����g�텗��|�K
��a�}�!��]n�V�i�<��jռ�m٘_X�U�B�D���5wv��~O0�`Ԓ����8yc�'��.�*�d����ӺJ�b�$ z>d�Y�?/�	�I�j�L���T���K���n���3ㄨ�A�:����ҳ��&�e�U�%���DK^�1�H�$�؂�+q�(6eJ�F3��>��֑nk�}3���c����IYi�K��&�}/��_�KR@�%���eʝ���tq��Y1�a4�J���l�M�zW�~��l����/M���ϣ�C���k6vYhڼ�g��$��,j���	�BJ���IW�S<-����j%�A6�Ѵ`7��;7ۃ����Uc���7y��"�p� �C+Yf�n=,��wl6�S��(-�%��n�bٲ��~�JE�� k��;�����q&I�֥j���F�TA�E���5z˱Ѱ1l�������w���v�����_���2�Kvt<�n+�-I�)!z+3O��3�F�-2�x�	�jz��`q�)Ң����� ƠZT��0s@ir�&<���T"��#k��+Ǩ����4��C�ޣ���FO&f��D�p�s1P%QJF��y�T�i����B�xR*����zČ�y����<U=�J"��˨X���]��&�\�;�f< I�b�]�cuX�+��D)�sm^���_�sT��BI�Bي �1�d����n>f�9��Ϗc�kR�>�=H+l�����`d�#F�X��N�^z�%��gvv��=�ܶ=��s�����%�H�e�^�2}pX�#�L�P)/�Y7k7��g�jeN���}}�j�Ζ���=�q������x
6&��oe����Q�t��D/��T���DTp�h���|Dk2��A@��Խo���1g����Ŕ$A:#�֬-��$o����$Z��K=���y*�ޫ"O����=���ʖ-�Eb*��C��c���)�}_ �z�#�����fR��Z=�����-�4����%k���`|ދ�$w���m'���h�Q8�,"�n5[���}�Žz������)=ۃ�_�[ó��7�޵���n�2�e�nKf�0{�n�rѶټd�oٱ�5Z��H`�<]��N��CY^�A[X9�y����Ɲ���h��-sq�1E��~�&����t$�w��Eт�Mg�7UHX����Ê�ۃ�x2���r6�$�62l�&����#ƒ����}<���#��H�y�@��%�[m�S�)�s�ٶZS�����v�\Ǿ��o����E;>��:��T�|�Wo���X�v�a��$֤���$��CK;z&����/4z�C��wj��v_����xV@�G6�$(�-�2���\6q���QA�Ҧ�%�k�����ί��s�4ʤ�x��N�e��̢*�<.�	��'�W`��4��+tؽ
_ ��
:0�	R=��$��d�QQ����%�]G/u\Re�x��Q��~�*+����*�R��T"�3�[���ͽ������O�KF���&�3�Y��k��3��w65�6Z��^���Z�VF�-ݷ�_ص�
�����p԰��g�y�-7�BH��
y���U+sAѥm+W�����T��j�{���ڻ�4-WٱZЬ�9��¦<����`�|'��s:�)S�o��
�T\I�궦j�u"�#l ޲�5�}DI�y�&���7VPi�J��l8^-S�%1�+����|��g���]��?H�Jb�j�(�V]�
n�W�yqR�)I����b,͟{�[�.Gc��>Ϛ��L��(<jU��L�`\�FC�h����{��Mk�ǢHJ��R�n5ZR�z�駟k�Z߃�����K	�''�}����o��Z6~l��D�?�bU�QՆ�-۹�Dl�^ɌG��ØDYd`���rE����N���KRq0Zw4�����;����ĺ̐�4��,�V�#-�Yq����*��U�Y1�V�>�L(�,����.���L�BȼUma̜��\J�8�L���{�D�R���qasTo,���$�/U"0LCC�4�1�45������o��ު��ѷ��ti�Q�����eyβ��NͲ�,l�[X1ɻ�2�F�����J��o>j"BF���HJ�3�L�^~W�0��YتV64Y��'7:��/�A�9N��y�B���ƈ,	�������`i�ȲU���/�^s��W�k�V� #��٤lP���4G}���X��J�yh�J!�,���1�("[�tD���W�
z
R f������7Ru�H@��JW��U�y���4���nx����*^z�I��,�.]^/��s5���I�`��ooTՑ����	)IoH�r������>����>��y��}�f7ߝ�hP��Ӂ�{P4�0z��*�.��[*�6K�U��Q�Պ'��Q��)y�v�Ў�U˕�l��I��l2_:�d���S�4[j�`4��#18�MW3�����������6�D�Z�V(�'�.Ѐ����V�	�(A��n�ϒHE��MS�kQ.����",����J~&�}�T�7H��3�������|���zt�J���[��h[E�����$x@"s��g�(��|2i���#�����l	�+���6r۝���sO<�l��>�P����۽��<uoW��c���U�]��;항�o�r�1��l���o|ӌhY����w# Yl\|l:�z�b����C;<��G'�/d�%V)4�	�q���fӱ��\���5�=HP�sV���g�!O�5���% ��MGsY뱙�8���U��
6�����Mlɲ� j��,$c�Է�������E=:�~R������~��޶:U��_��^�&Ӫ'������`;�;]?>��D͟{��n
�莦2��#K��a���g�X"̐�J64yY�"� o! /9�4����0C��R����>R@F��4�������?�&�1𳎫�(���v�WKlC�7�	�/*1U�	�c����'��T��Ca&�U9ɡ�s�֏���4��u,)�C�3�ov��x�� Y���u�z^�>���/�-A�TN� �j�'�; �P���A��֦���67|S�{J"ݜ�k��'����"����"��p�oI1K�<���_c�Zg��[�>�_�`��Ծ��W���f�n���˝�k������R�k�0g�:s�S��ђ��r)�V�ݩJ�������C��f�۹�`���p*�����ɥ�Qm�8%�f�	�Tĺ�I�U�g	���.���^̥/|_�á}�W���p�F��L'(��#㇜��$�=[��Lz��u�xP�{�I�b$�2_�8[jC]��T�^��"���S�'�H�A���F��a+VK�<��� �������K�s��h�T��j�c�>��DPc��}�s�T�(lm7ۈZ�>}��3J������·�۟Zd�-˺"9i�:v�-ذ׶y����r�e������.�Wt��sX�<�3m^@���(;<��{7�h��\�l���W�� :[N�¹���تp#}f��`�}��s���Y������1�ˈG��M,gk�+Nl������6#�X�<�tbh '6i2w}�}L�L����Ɋ���vN�j~�`�[����V�n���+
��e�F���b&�Ġ�HE�7�jH� D��R J����!_���?B�~m6^�[���(B�H���a�� +���!D
e�#�^��u���\���P?k���ɰU�W��kv3؋��(����C�~��J�R�f�Ǎ@�5��ڗT���{�Z'2v� ��L��}R�J�][6:�dB;9��ؚi�06#��o�������xp	��Q�6�]s�2��`I;�׋1�hYh��u�ds3����I�+�g�Y����s�"q��U��"#�x^j?>磊|*�����Xvf�?۱g�ٲBeb�|�M����h	�?:����
s�0gI�h1�c�'*ضEkT1#��Y�f�b�z�^{�={�^�F�]+��l��L�`=[�NF$��z!&�j���^i��iL�FP�*��O$���xL���W*s&!^�&��ܚ��
���WJp��t��&$�cW4c��o )k�_����汒(L Sj�e4��3�m)��ł3��~�3]�	��W��(�J�Y1�&Tg����;Y	&� 3�J@ӳ�ݤt�q< E�ݐ��J6�����Q�r$�t.z�����ɓ/>�����PV����/������5��hxh����fGg���,Wڵb�i���T1�% O�l�1#�	,`�`"�bk;w���ЎN�v��}
X� �E\�[6�?[T�T��SWwl���Z>�y�޴��X�:4�}w(��-m�l����:;3��Ͱa�'=��Pi��S�&9���h�i�z�����{���IU��g�.��^�"�7�l�������
���{fG'��;6/la���z]�!i)��X5(�hϬ�#�W�Ie)TfT�%X�& \f�bs�!ɋX�i�M��w0W�[�������;!̓�?����ಒ��	�h-ȷ��a����E �=DJ�{�?�Opu��;�z��/��2�YJ��7���H��>˴a�,;��x_�d����|!����q�;L�~�-Q�
Ip30h[���I���h�x�P?�����^+�yTȫi}?-��!4D)�{��!����49��C�P}$|�?�K���5��	� 0 ��z��*?�����~���պ�����7n�����(�26G��F��)\��Y{�d�&d��5�Ek��֪@��;�麽��M��+��)�f˜/0�и"JU'�qB���^��5*3�l3�M�8rn\���k�'q��1l��#. ���Fi��<)���EH�yo�ٳH�a�#��]򞩪Ŵ����2�&�8���x�&g.!�VB���K}o	�h�`��~��^��0|#�`��O�T�J�9������G�{2G<�y-I7ܟs�(RQ�%ըYd�����@��n�O?r��G���N>���d���;��ϳ1��}I��?�;>1��j�/nY��6j�E��.0B��)��TR��L�;�h��F�a�l6���3��&�����O��)o��@d�"�gnfO=�g�V�ZD��vv��w5���o��j�拜�I��t����j�I&��, ܉�����<q;�m(dV�kK.O��q�	������Hk��=�Z�lQ�B��v��k��9�ޮ�����m������p���u���C���q׳��*F-��q2Ip��3)�A[�35��~�ަ�5|4��o G�y�5�ে)	DU�=� �@ڏ�c/�\Ώkͦ�ۓޯ��6
�s:v��{TmM:9��v"���DkR�Qljlt@O{���:��ͅ�Z�$�OyXxj�t�1V���X���]$<�=��~�$ܵ$���5d��LlbU��|%� ;'���k�d�Q�8V~�[%Ӝg�V��L6x~WjV�T�PI(h�vDTHQ���Eʛ'�ձ91(�Z�@�.�2���x��؞y�n�Wl��[�oۍk�,��QW�8C+��*��M|d���o�]��^�
��UKk׊֬B�)Z��ܴk��ۍ;]�O[��n۔i�Q��Ζg���J� A�8�g�|&�\����Q�ds��T`�n	R$�HvG���2�r?�d�g�L���,*�7Wn��I�� 	�p<߄��漞ǜ^Ľ�3�>
�9�o�Db���L��������l�����8&HR<����/���vb�c%��;�?�Jٶ[M������c����c>��+u+�+B2��DL��Bf-L6�i�W\�X��E�L .X�R�V���.���z����y�C�g�A�{}�{t�V6~��pxh�bݎ��v������s�JՎ5�;R� 
@������&v2Xs��<�C0�9ΰ��X�i���#o��"�)��[ع�]<_����ڸ�[��M�{��r&�Xɱ�"���|�j�+�t��7�.V���i���
\s�����J���(�q�aN��v�=2e���#�_�~��Q�$o������'?oW/��O����W^�r骍26��U[�/�2������|�u6����!���xy8�� ��`��8Pj�g*$-� ���T��u�i�R��j�v�W6Ti�?=+g�'��x"��pT�꺲FԦ

�w���=`e�f����rQ�$l���X��qlb�&M`��R�0���S�j�8Y9�_�G-6{b���B��08_B��[��y0��5�^/�Fө�
�Ғs-[�]d�4��F���S��3IQ,�g	����g�0$���*��k��G�V�0b�)pDEIK���z�%N$|Zs�J=�RU�9ϛ^o�T�ְF�)v/��r9�v�l�Ϸ�T������*���v��]��6y��<�O�"� m#cᲰ���ꭹ�jE�D���������wg`�]{hk[��bg�6�X����Gc�T]����*�5���@9�x����4a'3�#��-���J�/���E�#G�[ίp�	H�,)O%�9�K��=���_���I��/�H�I�B�Q"�T�g#�ٓX�p�<z��ad�o�m$��;�zS����|ʜ����i�C��T�uq�YK�-�    IDAT���'����W.X�E��>��dn���?�b�%]�J�N��N�fY�j����EkX��hRS{B�4��l�M%qi�v~gw|i���/\����F�,����?���B6E;x_����٭{�2<�W�V�����K�D僠2����@O�;���lH��e��<z|f�B�Z� �~)�2#[�a~�hV-��T�+,�b�f�D�0�If�L��|U1��4�z���C6O�;6V0]���,Շ*"ppG�C�bU�p�\]
����Ԓ5&�5�h��^�o����'>vEf��Wm8h�o�έ;)��S	�y+Q9��E�01����;ҩ��x}s�AU�W��%[��I��9�a"�����Ksy<�d�>������P�����I"���*��'��׃�}gyS�F��o���%�+�A��C|��������C>�� b��Io7�4Uˆ�_RY%�`��rµ�$#¹G�W���"3ة≪��$�AM�'p@�>�58?7!G�֡<�7��q����Ծ@@3��:<�B%�g�,2^��^Uo����AЏf�Q�,��EH�2��`�5�0<=�L�L�I����
uT�V����<'�xz��v��v+V+l�5�j!�����}{�ݼuU{��p�gk�F�q%9N�^�Y���zcf���ꥼm�֨�bYZgk��{���}��}˖[V�f�70��$#T�$�����v�7, C�5*T�_9�'s{��@�H�6ѐ$�𹒥4S��x���% O$��{R䞰T��$�b�!������X���9$N�#x0B�6��"X2�Aŭc�MD��Ti�ľ�g^��ჵ�ǢF�="�"�ll��G.��KO_�NӘ�Yqn�gG6�r��pf��>��ӱ�;�ȷl��Ԗ�N�1����R�i�BM>��l�U�9k��Y�,ըcD����w�3.\}}3v}/��/e�'��������ߛϺ6�`8����vt6�����<L�m����5�%C@ �9z�Gݮ���+%'�� �l��h4��b�p,N�ި�� �a�f�[�Eπ�F�A�\j[�\�&;��͊��o�D�g��0T���xB��]03��sj>��WQEG�&�f�0sU�$��tqB����-�Y骚bM�~n�9�_����~䇞��oݴW_�n�\;�ɴn�E�2`�����ͦl�lzTD��3����}_�ydĉW�Y��y���ƻ�.�SO6���2i����u�( ��hC"���:�(F!��U�+[m�e��$��s��iS��= ΀;���HTű��#]���������'#���BU	}ĪWa���fLK�;�*[3}I�V�7)Uy#N�^���7ZJ@ $I�"�6!d*��+��D_4`y�˦��6n�����y*i�v�ё52*�'t��� �:+&>Ji6X,�ef�R�&��L'V+;�聇dk�DB󞥞ɴ�����OB�i�A�Q�L&"�fG��sԐ�U�jU.��^ն��_<T�Os��7o٭[e�f;���H��Ge[,"LC���
�Q64�d�֬m���%�ʹ��B}�޼~lߺ��f��Y�%����-��W�$J@��De{5���H!��.�p]B��J��ֆaE�)12FNB_��p��,�u��<!�NdCÿ|-?4�ӜsXF�����WO�CYJf���E{&�m)c%�� ���-^_|���LQ�����غ�إ�}�'쥧�-7��P'���زEE��*���m;eL�t���PP,D/��P�l�F������Tޚ�m]�.��V�e{��?�ĥ'������l��G�[�\{����G糾=>�ٻw�6^T�7��E������ٲNˮ��jlf��t��?��Űkg@�3�3�rp!^�(�$��u X@}�Y��X3���Tʌb<�{���+� *D|Ӡg���"�V�&�f@�Ǽ��*y)�67����O�BX;٘iS��Zb܅�����i=���h�f�nL���ڧ?yՎO��xj��r���
��#���xn�̉_d�[F����B�gT�)���6&w�A��|�Ϧ6şW���@x��nb�ݕ��(z�z�Te�|�O��F�,�Sa����KE\��
��>3Y���7����IN<�	*n�Xd�8!�B���5����GC�)X�|�D�;`4�x&"#���t��⵸&��k�r����Z߲V�hy��cZ�v@˼��Ʈ�F�Gbn3h1>��Ь�H���K��6���ٙ")���^0�^�y�ȗr��p_"��vѻcJ}p�x�Z���3��܇R�h��1K�.]��1.X�v���
����ŌE���v'����ح�5�ζm��L��i�Gu����C�� #�RF�`n�J�v:�2�,��j[��k��}`o�8�y�sۊU|�A<葻�+�{�y��ҕ4R�d@���8W�X�h,��S��ׯW����'�J�6dUيU�=��i�D�֎�^|V�㊊���pD+�,U���k���!�l���^
�NI����y<C�_�܃A}�8&}d�ut��)�a1?��\nُ~���JȈ��F�����t8�-;�N��wo۷�߶r�����T�֑q���3�Ʊ\���HZ9���+#�v�!�����~��KO�������o��;wn�O����ѩ]�}h�Y������A1�QP����v;u��jh>NRa���Ãǖ�UT�2���m�A4��:5A�Mn:��ɑ-�Sk�k��iX69��Z�M}4&�����#l��傊ȯ�`���N"�d3v��iGe;_��$�M�dM6'���aG��Q0r��	Vskֺ�+������vE(���;g�����L���U0�0t�����RI��!��Ռ`[�|��щ����4��,�p���(�T�s�����76"eʉ ���|3��@�T�U���ryD~N�=��\�� ��%%�b��˭Tk���M#�o��T"�QpIl�Hlb�6��@c~{���׋MD?cx>)�hsJ�G�N��B΂��LNL�q}e[R�1$�2;Α�-�BG	b��+�HW�-�����H�jA����416�6W6q���0vNX�\6w7�`��D<��i�8q����֮?��]�2�H�+�l:��t���US�B�rrz���\[��yvw��ē;��P�"��Y��)1~�߳o�r�޿U�ѨcG'��.7��[��D�`��N�f�:Vks�W��m�a"S�欁�sy۾�־���M�J]��$���Wu� �A�QٲFCv5�I��d$-�Q͊۰1��zNB�1����vz��R���&���������A��@��x�]�+�x�սO��0P f�VCjKD�)�����:���'�i�����H�{i���
�NP蓌��ʹ�=u�l?��/�Nsh�eO	�Ã[��7�s������q�g��yÎ��Y�������
�:]%+S������k�����lIu����?��K�`�?8�x��[���A�����}xl'����(��sd����U�W
K��u��j���"@���Ç��m8�T��w��e1=��Q=���?���0n5*
�˴BQo�+Vc�����<SU�e�dg "�Z����n_��B%�y�β6�<�0�d�_1%�0�:U���R�6�m���AED�l�����y���Y6Y�ÇT�M�w�v����XcF�r�$�d��#s��k4���Nsx|����:ؐ�;A�Q��[����?>Z��D������66��K����l�QS-�
����d����R�/�����ס�������C�9���6}mՃ��%��N
b��]ְ�D�=:U1�������=�I���ͺt����%R��� �Fn�^�X.����F�L�O�7�9`ŨL���`��	/�xԀ b���\T1�����Xޕ��9�����t�_�b�g���Q ΍g��TG��P�� �~�)S��3HO���_%W�U�f�ud2{�/P"�ȋϬ�.��.2�9�+(��V��ν����ݸJְn�.�8�K���-�5�,4T+�u�%k�8n��m��;�ƍc�΍G6Z6l�#Ѯ&w2�p̫{��u�z�I%���_��ҹ'>�������E}U����J���*!n8:���}B���7�=%�|�c�3jm$�$�ꥧ	~WJo�^��S�h��{3_=㔌��HN<�����z�A#تm ����USì�\�ȫ�Za���;f��>kۭ�e�C�w��ݼs`S���㾝�j�'?�qkv�v��#��+7l�똕�Y��blC�d_Сgc��UK�D��T�Ћ��t.����'/?��}e�	�z���������c;8��p2���5/�8YUwa����v��rm������<>�ÓSO)+�6��/�''/H����dؠd:�V�x'��w���lUm<�˩f��#؆ 7���£�BH�:86���C�IA,�'�
��s��D���d��ƭ�*A~+X(=�^8tHe�����g>�	;>�ogg]��M�h9���]�׬Zk�d�=od�l1��|"��l�����!N
Cab�����Q�"��Pǳ��0�±�|lK©=:��ב�G0�����Nl^Q�ש�ub>3����cW�L�t.�z3�x��6e^?`_fN�$�b�/����{�;5N|�?�
��DS�yg��&�ql�ke�y�ղ���xj�	��f.�Sp����D�d�G�k᠓���g�	^t9���5jx�:��w�6X	VIR�zA'�cH<�����n0�RaD.m�$$Pr16���c��ýzw�U�8� M�tu�@���f����m��`9+Ɉ�,DO xvim�Q��w�o�6U�������v��_߷��U�۰�؍��2�\�׹�jyk7qEBeQz��)I����VS�v�h؛��7���~�p7�l#���MlZ�߾r�j��]spF�u�5��'����� �Jk��$�����d4#�q]���^O�nZ��!�}��5��h�8�!��@[d���"�ߥ^�&����U�]��rˡݜ�J��;�Aք�ʔ�s��]����vi�l���ݺ}�n�;����깉��'��瞿�v���e;V,W�hVٶ	��^� �5z����z�:��+�.���<��|_��a�c��Ϋo��<<=�ó�z�G�=�M���Q�-�4jv~��
���Ʃ��D����w��{t�c:<���2�+�C� �xl�sa����gMr��ڪ���G�;뉀��,�����Uj��y��G�d�C�r��R��b�RU�|���~<P�R%��6[]�P����x #����)�;?�	�
Ҽ{����9�R�e���6�f����$Z�Fu>�i6�f�G�U鏸g�H]	��P� ?J���q1����� ��c!Q�\~e�F&��%��<cPEAfrpl�W���N5��T��5������Դ�YEH:@P��#��'I�A�X,i�����:�/U�:N�](Bl�ZM��זs|��yM�^�5��B�z$'�$H����S�-��ɰ�H��g�X�NΎ��jX�Yw�C��=U���\���9�`E�ec�9�k��ؿ`If�g�����n�����3����6���3�H0��P)����uI�8g*jm�02���~O�^"�U�-�s%:�z��^͘ 0����d�3�	֪�$��Y��Cq.�P,�ԇ�l�N'6���杞�����7*vzִ!�I6l�� �Ê^�So ȧ��.�4ɬ-U��N�ꭖ�U���C{��#��۶�׬�� p'E.�"��rέ�.���P 'ı~ث�;��9H`89J�5�|�=��l���-7���Je	���BJ���GeK����� P�������Hz�[��!SzO�gq���E�'�61r�aOb��-�$L���4���[O�L)U9�Y��
�=�d�T��Z����mO_������~�v��I�8����>��gmgo�^y�-����Vj>cխ����dC�_�^������V�5��iv4��p���Ͻ����}l��e�ڵw޿s���g����mo(�d`Ye?���ɉ�_j��Wʶ��c�JAY=�zgg={�w����H3�#P	=��`	��W��=d#=6�o;�r��
�i�<���26���˦����鄝��?:��Ebf�s��Ye=X.�MG�06%��W��^����ԫ����0U�G�˿������M�5��=���QO�i�<.7��ԯ�E87�;A�k[�4%S�.]����dx�d��z���5~����%���6J�|�ɬE�KUGvL��k�%���$'�gz����TWz<d%)�y�2T6/.��b���7��( �,)�uH�q�!'�d%>�1���r�qҋƄ@NR6.���ԍ�� =Ɂ�H�6�t,T�kC�\�Ԟ����y���I#֌�'s����;�V�9*�����-�|$��:�M$4�=�SJ8$&��Y���AJ��'�� VF���,蕖}#�.4��}��$;r��'y�����G��}
B(!5�[��P��[��3��I�n��׾vho�U��Ӧ�quG���}Jr6S�-��Ts�锬�`/�;U�jg{����u��׆����٭�#�X-�U�\�x��	=flc4�
]}�ZS{B��׎{ɚ��$�alM��I/=>������z-:šX�P�����Ǔ�~9_G!�$Pz��ю�3ޏ{����Hld��ȝi��v�5�ٽ���I&�v�Q;����)Tx�$}��) �֩U��M(Z�vxҷ�df��;�*�m���G�۶�~�%{����k��cY�-+��(���ﵛ�7Bnf֨���(J�ZU0Ix�vv��H�����O=���/�-'����_>>9��ǽ#;<;���c;�(Gә����2w���Jo�����zxri�V�r��ݺ��޼F��̪���B�P'A���1D��6!.�t4�iַ|�	��K�-��J���^��R���l4f5n������Y�7�nwh3�B�̰�r+5*���urR�IT��'���/^��*�.�����j?����l���e���T�$3������Њ����/����S��}X�XM�"�<�>��`�@� u�a^G"強o�k�e�M�W�Z6���G־��o*�f��a�"Hb<䚱�WU�*I�-��?".i�F�띎�Fy�`O�[V$nE,�%�5OE��������I�$�@�Q�3��'c��ԧK���))��w�!y�z��7W5��}��ZD�yo���:�P'ËV���	�k4��#T�"%K�.��Ӹ�C��.���F���}���n�ד�M ��*΢WT��͉S�l,�����B��5��9�lvb��4�������}�ώ�ڵ���[6T�{�돭��[���uN,�V;g4��$�Cɸ��4�Q_j����gg�����C{��Ȳe�W+���-ʫ��E��U��R�fO[pP���8�-WC�ƍ
6��N��	�!�%T#�d�a�x��9
�OV�(o븎;�Ʊ����N|:Ml���I����G�(R��c.������?�^�ӳ�D��Y��.E���n��:}.�+��9�`n�,W��'���{���:�}����?�)q ���u��ll5˕����jŊ *���m%v$��*������ٳV�e;[�~�٧�~��&ؾ��w���/��!Hu�?����N�lFe#҅o�A����2u3��gV���ZiZ�?��w�A[�W������ ��3te(������X~��\R�Y"�1B��ŧ�0Z6=���.b��I/�=<�bS��
SY�L0ɴ�� +�١��L���d@��n��#����>����~�����Ye7-g}+,��$>@
k;yiB2�%�@Y~l���^��]A%)81����\c��?��T1ͺ��%)0!���b���4�XՇ^o����$��u� �#%1ZD���Ge&q���H^�5p��*9I��l��d�ڬ�ڮ5�<��;[��<��q�5����8	3H���l��U>    IDAT�N��s�F��_����?@�T��znO�X�1o9�-�XU����J��9�mP�f�y/U�J�(�^�����Fl�u����?�l�5�2�
�7ߵ_+�Y�������3��
�Q˜:cYf�Y_�����r�����{#�ҟ��o7l0ڲ��$#5D�'V�a<�B���D���N�$��R~)_h��jQ�6�d\�W����LV��(s�T���/���<iT���bk#?����>�<��R��'ҡT����m������/���Y%k˥�c�d�f��hK"N&�\c�}3��^�6��t(	(�C��D�^J�8�3B&1gE���jR��H�u��p�˽��%G��M�|Q���%s�5+�v��];����Xy2�Fnd��h�����J���z׾����su[�q<*Zdk>�V�!�� ]��bŶ[{�ll����?�����}l������z��]S`���Nz=M�!Ȯ��c����K�:&�6�Ǝ?k��K'W!��+Y17_Z4R!GIe&(��x|�Q���T �l2V �T٩|N��n� Ŋ��~ C�i����-랍�rx`BN�o��@wB�V�Ez���o�!�\�?[-� ����~�s��/�����M'� &@ٿ�H�AG�PJi(逝���c�%W�&0O�CQ��RI�}��8t,�@ �;t��k�UJT�x���=b�_��C�2zUi�0W�����jP�L�P��ң��rWX���q�Z6�,�!�E�Zߗ�9{Ktm���הH�����5�2�4�D(m>���k�^q���uܣY���nx٢C�h\���*W�?����l�Wv�a�*Z�mT��B�2g��^+G��X����	2�t��"x�s6Ÿ�a����<hs�Φ=�Nl6?���`8��d7��W�|dﾻe�ٞ�K��'�D��Ւ5�@�s��'V�ϭ��Q�J�lg�i�[e+V��+��p`�������L�?�]r�MΊ˪8[�[a��*!��%U����-�
7�w�OʳD��ω*�d\_smT����vX _
�2���	d�E�|* T@陜�< �x��'���{��%�)�:{r���/���͜�'�%S�#�K%���(Sݢ@�XF���X�$~�ӶZ�}�*A�;�6X�_�X1�Ye>�O<S�����(������޸c���Kuiїq[��>nT�_���.��-�۶5j;v�⥿q���/����wo�}p��wN�������0���폼�ņ(�F�=,g�a�l�G+�.�FAR��+��<�7�Q����Or�`���4몺Ն3�=��j�<dш��֠��Jh8����в�S�2�k7�v��%�v��=t����QM�zs�[�Xձ
��k��wmZG<T�&ؗ`[���~���_�i�.߷��t@!=��+�r�d"�j�y�5x`C/u]mFD��������LJb3��d#gc��MN.�9яL
GA:�����Q�*��6�c����ڔ�����V��E��A��J�s���77���W�u�HAd6z�k�sݟ��5z�v
�m���v��Q�H<b��D<x`l�1j�����>�g��#	P N���΁+H������`�	Vo�pJ>��6C8	䜬 cdj�����T�=
A�����e�Q �I�2��k������ b�A�n�;��~��n�ܵl~�Ƴ�e˱�������]t�܋��kx��lg�%9�^� ���4��;�?��{v��ٲ�c�V��K9F��'�z�6�+���v����7�F�zԵ,�V�s�#A�#��Yb\0�[()O�l�(��\y|�E8
��0���42�3��B@"yJ����T9���p֘WÛ���|,N�d��:��hE������F>����!B��^.�
�ff[ͺ��h*��ƶ,Z~���|h/^-�_���v���ݺ`_z�ͫ;��v圛5PH�na�{-�ze�M����[aQ�F}Ǯ\z�G�\����`�������7^��s�s�Uk�զNK_L�lе�hd���Ñ@���I������ҽ+8�p�����g�A�c�l������3�*%�g[L��ݕe>�N�v�Z��5�52�w��zg�������4���vnoK�\�7����2v���l4�>0�+D!���$�yl~l��%x/���\)t��	�ǿ��f�[6ߓ�v�X�ܼ"�Fz�4Ɛj\R��X�b��Kغ�{��� �8�*06���몂I��s	�?)���d���;�Y���^�*��Y��SF���a)��'z5��/ɀf���3��� ����޺�GY,z�nϺd�̓}*^�;�l����mv6���5迮#`F@&�E��BD���}�ji�In&�����GR��w�(¯a">����z$��-Ч�c�i;|�D�"R�̯D'�����d'kT��w ��O9rmgDh��߻��a���Ӽ�}�o/�ܳ;�wm<ݱ�lh����Յz�Q�v�U�'V,��fǔ����Ef`���۲jk���쏾z���U�l�=A�<��l<_�6v�G�@JR�:��VJ.]�6�N���Y����C�
d	����z�2��6���h� b(���܏��͐�\%6�M}]�Dfqc�.P�5R�A�~�0�˃(�;f�]Y��1�#�m���#�%��jW.���s����Q11�<:��Pl�d;߬��K�#�~Ξ�r��>:�?z��u�U�n_T;�<]Z�X6DZ8��Ė]}�Hs���f�\%kT����>{�ʹo~��/��|�߹���N��{A󭰋�3T��7gc;��N\.L�l�>J2G�����F��*[�e~OhH���˾.�& ��˦C��9���d�l���v�B�v�*���e��w�����������TՂ]8�cO]��^���[�?���l�|�D���wHPa4�t���$}c[��n�^.Fi��^�O��y�����n��M+��d�����"i�:;N��Z`���=�E�{67:����P@M�f�'A����L�8 ?�C�Q�y�:�sm������L�T}�C��+U}`�%�]q<���3oWu�3���C�U~D�%�C�kGf��BD"�\5� �+i�GbI�/E�4]O��<��J<���8N�qbwK�{�!�G����C��{�Z7�W�)P��#�ظ��'��{}�|�q�{��'�&���]Y�Q����O�'�-=��D(�eg�{�������ӿC�-��?�I�Ɠ�fg:��xiGGf��ڷ^ۃm�ر�ldV`�#`C��P�өɿ�\��VٖӉ�"_�s��[;m+�;���3��˷=����l�r�Z�˒�{	KXω�TE$��z]�XJ�f�~}�H@�+3G5���w�w����-�a*��e��F0�a��n8k*�tH"6��~�}V\շ�ax�3��S�@�� ��%NCb���w������h�o���5��+r`q'����C�_<��"f�y��s��KO�Ž�=~x���ݷ��Nm^���@�][�s�r�C��]��V���o�o�Y�*;�-o+�r�(䭞�Y�Y���?g��5�;{��i�):�[�ē�ԅ>�F�����o���{�z������Jk7�v��aHlCT�Ύ����1o�z`�L!�H2/�"2�%st6uԙ�2[*[J��x���&UmĪ[L����&�q�E��.]ڲ����۲�`������������
�F?���tl�Od1\���w`j^f�-���o��,9����RQ��_������V�ܴv�ge`��R��)B"^A��QيҒ*x��[R�o������z�럄��cAH��h�s�"	BA�PE�z�^�A�*�����2�y3pF��?��2�zO�d�]�lu>����0���!=1���R��vEZGR��J<6������ùJ� �F�@j��M^�������*_��ݐF@�r��6Bt�Q7���R�l��3�u�����sN:���ֽNs����6��>D�g��������q���xg!�Z���}I6�M��VbݰF\�8����a{9�lܵl�S�%�^.+�hno_ڷ^ڃ{6���-W`-��1T�{`n�n���Jmf��u+�i)�\B4�(���Ζ��;������W޶�^�
�][��%X��QU[��>"�'��VvQ���f�Dh�$��в�g�2�Ǯ����'��y�~8�����ֹ#�iW����
��$S��{����'k�E��	�*H}��!��Xz7���>�����:�{���ĈVa$������ ��u*���fs�3����~�{����߿mǧ#{�����l�,[�V��E{f��/\�v�nw۷�=��f�ڎ^��,j>g���.�o�3��I��p��Jź5j���TKm�r���|��+x��_|�j�=x���K������|��޾sf��MsH����4k��C|a4>���h����Ke��A�dN�IG+��BRߖ
`�� }�o�I-��g�4���L�)X�;��������=;::�� A�<s��F��gg���ƀ {9� �,^m�i�M��Sӆ�LU��Wy��B�(�V�g?�m�����UoZ�������C��fV��e.�Hv:�)���7>
&ZUA�t��L�o�P#�)�ġ���0<���a��N�z�� �ɾ�^�,���
�:����9�W�!`y�q��Hl&�>؟���ʊ�(Z�ASK�C�ꏖ�z�ZO=Z��S���u�^�����:���sl�l����z-�Ii�`���D��n$4���x塻7�����������;b��2���@gV&���+���*M^�������y�(20r���w	h�A|�)�β��L6�ٽ�{�;C�qcnG��67%��� ���A1?��V�*ՙ���.��,�E�� ᛫o�H��-����폿~�z��M�a�2������V��%>�I*Q&�iԇkE`EH���;��{%��d�@ϛ��O��Y\֗���h����SR�|�a�;"�vk
�9� 繓�"�%��
���W�)a��xMx���,�/i}��Zi���),�p�RPOEEM�T]�uH`FP{]c=�񙍲3M`�>͖��𠥺=�O}��������Gv���v��c�w׬޸�r��c/��ɫ��sW�0��WX�z���bC	ђ���c@�.����6�z���&Y.�]�{��ٓW��k/>���h,�����/�v�\������׮�y꽇��>��ɨ���
�~��V���T����J��\��Q_@�(����9	�K�����q��lɳD���:uyCH%���V�٨i���Ce�̨�L�ҒE�93��y��3B���� ��74�=°�}Ro����<�:�6�bޚձ��t�~����~`�܁U�&�$ �0���&җ��ȉe9�ȇ�
���a� �3���V��+%1�Ŧ
/�w�4�*�ƻ�C�^�jC�  ��>�fp39��*�w�����=ˏ�`1���j�Ĝi
:��G�&���$��6�\T�`8H������=^�)҄��r����X'��=py�C�ʇ���IkJ��\��#�����Иב��%�9%XF74��?)R2��$�_���}OI`$� �&9�	rO�v:�b69�7��݇�����n�7��Ӷ�5c�>[�v�Y�r}���Ejn�����Z�.�5E�B.HCӇ�-�-��;�\�lQs'�B]Vm���I͊����$>�Sp==я{!fvb�k�'��"�&S�v��N��H<]���2�_N�T�kJ�"q���	�s�=��<��Q��'ף\�v������W�+�XPz�@����Q��}Y�V\�9���T�S�˲-'��Nmxv�>��]����+����n\߷���������'y�c{��s{v���v��C��+,_:o�ƞ�3t����m7Z����ǮX���A�
��]�p٪���쫗��ؕO}��{�]��o��]^�����������o�����=���k�2;7vg�C�5�i u�3y���b�-n�ʈ�1|Sq �>�UcT��	�>`��ك��#_�&����	��̭���� �����'iFf�R�%�b���$V�N`m}&q�ѹɸo�!
���TN��`��o�:�K��������U�e�-���ǁ������,�뒰��� %<����~�4�`���VA+���1��5+�)��WS���2A�Y��6�K���p�r��������#Rծ+�5]9`\m���?8��6�m��ڍ�J�`Ǣ �*��@p:�P�Zl�}p�"�76����Jړ�������M��'!d�F/w�h�ae���=؄W�XC� ��e3u\l�)��)�䘻����`��\ m䞀����B�!l�c�a�����̮�m���s;<m(�N2�FO�UJC����Ǭ�t��q��EؠB�ۑ�R�m�r�^��M{����FsF}��X�Ҳzظa3�O����b$K�,����&mUVe��M�I6��4�����HV�����=�A�� �Y���GzYhwv�Cr�&9$�Mv7�U���J�އp��qo&{VM,�d#�2#o\���=�9�e?��\@&�������<�t+`�Ky��g�ҹ����|�9C�����w�|���.�ij��g�"	>�SM�Nn���Z��$�#�lF���#d��b�Qs��$6�_��jY#By1��/~��	U�J	˺�5¨���5��_{O?�D�{��v���	�z�!Ƴn޼�������Jx�s���=�`XD����X�爳@�PB%>����Խ�3LfY\�r���Z��6�~��W��;��?�x�#<8�=	+C�b��fî2�B���1�}�ܜ��9�936uq�W/#����ͣd[�b�r�p�TC�'�6*�0"u�0*$�v0���9�����<�	�[^�9aM_;BɆף^q�ô��27�+�r����^���k������x�f��d'C#_'w.�m%(]��#�c#��Ŝ�5T��	Dg��=^ߘ���x��@������`�������7\�Gw�7���Jڡ������7`�q��=�+�I��)���Zv.���+UfY+���z ���˜���}��֝����^�1�����18y���2[���%bw�~<'I>;W� �p͟�����ri��u6�j��*'F�A�jc��Q�tf�0�9���M�l;�QR���f�� �[��}o����J�YKpT�����M��Q�R*�H�<�%:��*W��nK� ^��^{W�6W���4�4���*��"�Gt�V�;�e��`K4��z� �ZI|��3�"�'�����y�'S�_&�(�M��2W�䓧��ЋT�`�m��=��}��.�_���$%h��l?!�%�0't�|޼�@9��/�RѸ�A������q���ed�Ed�3�
D�3|��:>��-�+��4���t�3<��'�E<��ӳ��h�d0�Ĉ+i*F�[�s����`m��G�p�b{kk���."\���ڕ�ߓ9[:�����s�p��{C�?���}�XLƘ�)#6So%�!�1��y�VY0��q�l=�Kz���1�S�rB���-7�zD���w��lÙD�(FMh�PSl/�S�ƊFD�.�*J�,����Cd�"��6��6�rYnS�+qu�k���$�(�M1�	V*g����x�����#�z�� ~�ڜT��g�XLC	�}�P���d����c����Z���uԨ�tf�e���i�ʴz0��g��Rs��3M����t�ꡆq;���ZY?}�fT\iɳɐy��W�0}`�=WG1�ߣ�� JI�h��*n��|�v�iy��^|�_C:�5�����ř���L�����K���x�y�NWlaA�6��^X�`)����@{��a�4׷���z�IH�h�َn�(�����?X��[�}���1`5G��E�j>�	��V���JI\��go���̾˵:�B�L���x����e��    IDATL�5d�U���k<eF�%�w��2���fj/)h�3�}J;T��`�[*��h�55s. ����>{��bՃ�γb������$�1��|m(�K̮O��c�N�����`�ݭ��6��1S�P�0{j}|��>����6"�k��ʕr��mf��

�a�\D17�Zc�^\�sϬ"�!��{{{�Lc��\A����ޭ;wqx�B�_A���ETBo2"�*��l��|�o\��ׯcww��X_����e���\��Ս���?t����w������[�ٳ�t�GLgk0��d�A�9������pAR�2E���H�K�/����D�mq[�c�Ҕ��CI����S(JI�Ef�%ͷ�Y�XX#���"����M���[�0.Bxq���o���&wG�(9�\�b�D�F��rr1�Q:�?����'�B�C�����g"��lb����5d�!���^��'��#���6������jU���`C�zٝ�&I��;�e ����ЗA��V/�B��8����'G�⥳�v����(a�2�n�-�&��'�j���$�|�9Y��X�D�?_el˚��e&����s̿Y�5g�xs7��l�������ۙ@�3M����?D�|nD(�gf��|��� ��5�ߥʟ���`4�D}b`���Y�@�I�3I�1u1�|���NO��_(���8=+�3�i�cD�2���X[e�v��f�f���%�9"���.��+�u��L?��[x��1��M�r9�zs]d2(1`ۀ�)���ٺn-���Cб�k�Y[ig��MkJ�4.�P}��0�=gA�>V�`5�Pa&���� $^��r��v�y��N��r���۪���=_�&9]��=�P! ��w�9/�N^"�Ty� 妲U,9ǹJ�
jq��_�ň2ml�f��a}��gr2��Y�Q������ν{(����F\�a���ְ�qv�����x��^|�)t�m���R�aue�bm��}���ٶZ��������{��7���ߙ�K�SPMcL�a��ZL�Ȏ��M��E���-�����Q�8���hC��Г����RB�d�f��^l�# f�!J~тI���9V녱��$5pZ;g�	hU�'�фRf	LI�v'1�M279(�g�A�ѻ*?�Hhg.�cs$U���������#B��"#�� s9��\yX�'ɼЛ b�����jI$�Ϩ��;�$��ʑ��]1��')���Xa0���'8��0��w�0����֎e3�V)`�nQ�e\�az�4ɪu�!���(�g�P'z�^Dfx�8$����8}���~��ȯ����"��3�e�).�D�+;~��=iw��gٳu�Gɵ���5���f�`CK������%/��\>�p|��yF��6�O� ��`<(��H�|��9���j��d��ޛ���<���ì�-'	ʕ9��.��P���l�mk��E��js*��ϼ���Y��|q�|�~����fW0��Ej����Ԝ-�9�����A�עā�[/U<�4�"��xE���ׅ���1$Rםm�9��qB.?2����G��Ť�L���#U���|N|I��!ٌ���Z�ބ:��Y���}��E]c"[l'W��? ����(oծʐ��Η2{�T1ʹ*QI �"�qn���X/`�Ʉ`
Baڝ��k��=�K/����m�����	z�1������pu���z�Z�����2*e���ؾz�.]��`�:;[�������_��S�{��nh��h��C0�҆���9�m��=+'�(���"O}�XY�$�@Sd�@mQ��t�9��Efq��ii R� \ �t���x���r��9i�M}8�{F%3�$��hH] ����(�-��,�4�Ee��۠<���	��P�O���|�E��G��'"�HR`���D(�kȅ�L�њ��*��hdɄ���	�E K_�P��~�Î�'���ֲ43�t���3����O�t&��%s1�6��lY�c��8{l/f��G� #0z�Q.Y��]��-3[�[�]��|)/��B6�vZ�O�ǋ�6}�đr.1�����t�2��������4�	���_��otᇴ�U*ETܱ�7����q������L��� c��z���]]s�v�no��;c����wr&B0�a���b�F#��F�7�gh4��M%sG�D����ɋ;�fpis�y�����wv�����ެ�)�g[�������(���,�F�ENA{��� ��|^��@ش�m�xۉ�m������m�{��
?���~'�S停2���(�w"��L��<��B透߫҄u��X�HM�4�h�`)]�9����>1�#�tr��d
j��Û���(7Q+��Zgen�(7A.���Z�����`�-h�����짥�L������@é�[a�Z��Q\��j/<w�'�ȡ�B�\�U\�t�kW�����F��9��ß��������L��ɨ�����ɾ�l��|�l�l3�����)f�9����m�Ԝ�I�g��DU���4K8![q��%>7Vr������Xr�2�0�'5e鄹 C$��K����@#J��|��}*+
;C�2��4��Yv�dd�� �������T�	�!���t�Aˡ�� �U��f�6�4IΟ����;�����6q@��ܘ��U,+6��W�7�t7�N�V��G�ơr(3�x�l�4� �U�H�lɿꁄ�J�ig�$R��Ren��0��aP��/T(~�vN8\D5{Ƙdo�9�.��}AGڱ���k�&�����π��7��(�[^��>m���b�l�L�Q+�����[�
3�^�0pa���
�x��˱ Q��I�$�H�yz�Lf��c����dqzV�xc4c6�٠�{��9����-�Y�T���%�i�E�K�+u�u�^����An�q���(sT#�9Ҵ�u��t��P^?m���i7������� ,;.H�0%<�x@B;�Y�*��s�Z�규�3��d���s�v@@F��-�����F�f�a�ɶ)���v��9��*������ہ\���PFUؓ��k�T	��.2�uO�Y��6��|z�A</�Z�Ѩ�x�94W�������Op��5ll���_Gn��8ʖѨ��s��V9�A���|	�[[ߺ���������#�y���Ə~���o����|0��l2���##�g+��H�=����>��@�if���M)�6����ڡ<3�a<��s�kt�Y�0$~�RX��ZʺɃ��`\���AD�y.3a��D�_:aw�<?8����u��2����t*���iLc�G\*�XfF�kζR��[_��o|��Bfqv$�nq�f�-؈QVf�-ed=�|�-����hӐ#\���Ω���;����KRFNz݉��3��~Pb�C/)D��"p����y�1p��f7y|����В6�>})��os���abkIB�Ζe,��[�+�^wg�~�;�m�=t�s������ h9b�waM�}�6="��r��,�g�>��6��/G�BO7�ӗN;��$.� ���a�3��p�n��t�$)���8<>��1����ࠌ�.	-����b�͍26�#�ԁ���2��t���ƖI��P@����KT(#�V���?���x�?@Z�p�?�#G���M$����$�����rm�0��$	1fa����s���r�ꑙ@;U��=�C���C��*υ�h�� nr�"!�R�����*o�)(i�t��:~��v�ԃ"���wS:V�V35�[�D�g��4>�Aa#�A3�7��0C�N�Է%M/� G(UJ�q��?)�W+^x~�<{E���گ0�q��M|�/�������BC�c�F[k�Rk֐Ͱ}���+t��3��ݸ�TP��>��9�����򋟿����x�^�����h�X:[� -�K���ܷ2r<!�џ���X�P��L�S2AG�֠��4�d��`����]���-CV=��l3o�|Sy6l_9'�(}��I��Ir^V���"�S(t|z�2g4\�ٺ�VԦ�eمΖ���ը�o~�
���2J�]2c�2+���Ψ��A~ND2ƍF�6O��"�0(�Уl4��z�K�'�Wu�<�^<3�
Ip�v�0��g��9wq2���_
$�;r�>��m�>r�Q��Wa����-���8[/Y�����.��@b��(�5�O'����C�����}�ˍ��2�;����,��]���l�ߒ�M�]��a��3۴�����Fҟ�9�dN�J�iY�乥+$�,����Ύ͟Н��ݛ-�z�3�T�"�Bs�s�����w�p�v'�&z�:�]�=d�cl_��ʥ"���M"����|�C\��~�a &�Է#7o�VE\.a8~��{�ٯ�Չ�/a�Xcx��C��ؿ��R��Zd�e��,2F��0O���if��%%`�]�U����%#�'�36Q�'2E�{�<��+���#.�r�}@���<�h���XbSԓ5��C	��'IG���`C]�Km8����QF�*M�"#u ��G���y�u���{m\�R9�(����#���w{��#���gq�u��޻�}����ؾz_������b�I�r�l�j뵼�(��.PE>����ooo?����~��|$�-��~���޸��wv�xҞ�t8���IA�nF��aOz�������b��b��+ڳE`��a�#p�22T��ר	)�-�::�p\ӓ4c�i�14�m�&�	urE�n�u2���f�RDeF;07 {L$�ll����UD�GG'h��`b�xP��٨�9����oJ�����.9�|�|e_�r��.
�!2����s9��f@lE�<%X���<�QD�m�86B��� E�28[�鹺��}[=!�IW3�	J[�o����w#~ް[6�vFˬ{�7�����SHz�?dji�l�K�.�L���� f�� #�0:w���~��'.�������b�e�m��������@ꢳ�LR �p���&7�k��|�O�&��t���fI�X���cr^�:g{�~,g̭�,��3�i���L=���5�2C�G'�j��ǭ;-ܺ�E����x��BX����Vj�*Ds���%K%T�Eeb�EI�j��m�!WdO����.������m#o �F҄+`�,��K}�pY��c���xf��Ԅu���e��6�\��-�|ۛ��l�K�=k�e��!xňQ���N�S��=fbZ���l����!Bѐl��� ��F.�D�grJ��O�����et�̀��F��%�KY;I(��0j9��p8�P�VEy1�Je�o�\�T�O_�;���!�+i��cϾ��߻�ݝ6��M�eI�գ��(�.�@��"���������wG�a���8�Gg���՟�z��]��d�����'�^�dH9��D	Ȋ�w����&-�-(�et��<��-�l�8�'\���ٔ�x({���2^=hѠl��&$���ї���Q#��Sx���	�>g�B%Gq �ƒ�)�\F������v.>��,������"E�t�R�<��� ���U����.�E�������-� g;Y"�
,M�gˌW���6�(����9[//�a�̖�t�0q�癘���9��#�=�JWΗ��eX3&���!-K�FϚc0��㿷Җ���4�	�=;G��4�^X[�6�Z�qY*]|,�S6��,��H� "Q�I����r}�Ƣ|c�-���밶�����j��.�-�����4i������7 X���y�2k�3�7���#9mF$V�⩜�z�ҳ��9V�Vea	Pfs,��^��V��3��pz֐��p���d���kuܸV��JV����J�y1	*� �S�^w�z�����ȕ(U�8�񳟿�7�:@�_@��*���r���J`1���U��@Z���~�	3P�t��=������0����������.��NM5;�l3о0��/aI�}A�����9U&���>��WV�4*Y(��$�+TiL��E`�y���A�Y�ֲ���,�E������5�H��L�G�DJ�1�þ�"�D�|(�`�>k�(��z_��3غ\��！ÓC\޺�z��8����]���������X�[��X��Z}�问��ի��~��wv�/��o��/���[��8E�.f���D�LL	�}�Yd���eyyB�����qr�$���u�y 5�!��z�d�*�Ij	��_&��3KE�#���������͠���e�9�ћ�� m����q<�屸�y-,�+����~�HW��H��@�eG�����W���/�Q��PȘ��\�3B���E	���@V�a���J�[ !��FhV�jC���Μǳlc��0���KuDv(''�?IgPiN_ݟ��:0�g[2s�v����Y0�^δ�fK6�Л�5� ^_r#i��"��RLN���3}$����/+�vKg�鶅��yG��6<�T����%M��a3��� ���8.:�0�k���q�n�MP�~�z���?7Ԯ1gk�Rd?3g;��q�>��^����#�J���8j�����89�a23u��b�����2������V��"���T��6�R��g��v�(�bl]]E�D�Xz�{���)�}��YY ��"�T��5ϲ��y�� )躲�3U:[@��A�V�sS\�Z�N�#����ێc�:X�����^Da�A�)���)-c?ɞQ.�3�>�l���ٌ���44�Xn^��o济FC��h'&㡰8Q>�"�h P1�Y[YE��Q�bo���]J�"�|� �U�(` <�@cEdHZ3����Ѭ��܍\�n�`��d!���^����x���U|��7P)-09;Vu�X��R^A._���?�r�ſ:�������d�D#��O~��W�>���hM�a.g;p$g���Kf�c�Hd�],�d'#��c"��I�E�=�L)��~�����x�٨��7)݄yB-0f&���|��m���ec-FR�љ��˙?+�Y�EbmE�@"ҍlVY,7�C���l�	��+��dن�^����\d��E�,��gqn�z~�W����|1Vf[��X8��9E�g3+H����(����,P@�L�,3F��/s�Ƙ�$�H��3�����l���^�/+/���C��s*��#8Ls�FG����nC��<�W ĞZ��g���6�"V&�� E����؊����2�w�]
8���K�~��/��T�h�c��\e!����X�I�U��<ӧ�U�v�˿O$ӟ��Yw,��X$R~�}��,B��Ͻ��l�JթL�tF��� �~K	4�r*�9�힜-�~N�3��N��a'��g+@~�|n�˗"\!�9��Z�*�x#t�cL�D�P���QY��*&��#�SњJ��9���~���"�������\���=��:c���X@[�����\,I!h���|���R M�"��?�*5Qf�н����,>m�s{�� �P��؞Qf��8Q�����3�5�,<���ֵn�F&s��E��L�$L��NTu$y�LεH�rQ^�S�6.d������1NOOq|�F>��ӟ�l0�h���"o���Ҏ�J	�Ҭ4ѬE�Z�ak����:����1�p���ƣ����Ϭ�k��fl����*�u:�?��z�_�����G�H�����ۯ�ݯ���Ǚ��tp2ʡ�^����a笟(��|�Ǽ��|�Gv:���D�ŏ'��Y+#unV��Yb١?4B��=ztx|N%��T��2�4g\�`i�J�	��7��WY� �0GEm��"|���ȓ|��e��xn}^�|��,�N[A)���X�b}}�RY�+���_`%�㋟Y�|.�r��Zq�|f�l;C(}d9;�H=�/�Ȓ!z��yк�G�0��g~���s ��IH�E�Ff�)�3��k��{���t�Կ�H��6���,N�P���F��F��Y�,Xz��w������Dk�er���
�>M@�$�_:�#�%    IDAT-�m$ʃ/������f��?���K;fH�x��<���0EbZ:[�Q�`�6	rl�v��F�<i \��Yf�C��{��&k���-̡�Msr:
̂�5�C$ӡ�5꤃�t��<~2Ã�%���N�gb��D�N������<�i�b����0�i{�����ڼ��9����qq*ɷ(�(Q�N［�[�w1����Ŝ�#c٭;J�?��G[a�}���9b��M�P���$���r��ٻ=��+�2���f�KE�zI!���z�b%(�-�:�>��( Ƀ�{���hW²�V�.C��s1[��x0�~|p�	F���{�(����N~V�RA�!������Om�� �Zg-k����qMZ�;g8<i��idr�q6��899�$*��S'�#��L���R���Z8��pxJ@m�ª
�+5���.��JI�f4�"�#�E�ַ��ֵ���9l����wo?:��{C<9�L�2�y��I�MjEL0t���^��D5�ɐ�@3�t;�Z��7�y�?U�W���R�!��f�h��<I%h��sj��q~���9��=&"�D���s�3Vփ#�˲>���/��"9^_�QCc���W��`��O����:m-l�"sd���r��!o4��^� <@ÿpuc�W�VD9~��lG�t�bI�`B��Y+	88�@Q�q<*�Ѣ0G�����i�Ό�`��)*V���Y�����A��	����,�Pvd�\��tЇ�?�rQN&�1���:�$e�����?_^b
�d���}L�j��.��>��0�TbZ���U@�zvɵ�,Յ�Ճ/���U`���_`%��oMI���@@�do�"4A.oԫ����,��I�kR�fp�h<=�U���qy��`ɞ:;����z�r�Ԃ����h�9�L.O	
Lp��5�����U�`R6ٸ������~���Fk+5͚�c�C��]�Y��R����M����I�@+�Yeʣӛ�۝�ӝ�����6&��U�2Ѳ-E�2�
�XrȞ+�H����kcwcR��A���霽��t�����h؜}TD�H��"b�9yZ~b��Yb5b�������֕]'��H 1�pi'yTb ��g�d��� ���ep(n�Z���n�''���:~\ȁ@�Q%L���ޛS����l�A�s(@,�{��M����ߗ�@w@�*f�\�N445�̄m���L#��-�C��AI��
,�S;M�ZD����+u�7k�gt'h��q��_�|y�o/��������O��}r�{G$�`�SĄ�	�6��FBǕ+E��G=9��b�b!LgZh���g'�O;99�h�Ӣ�n4V�Dc����4**��H|le��c���..:�S�`���:Q����bd
�������,�A�W��x��#�m}����U�m��0���5���K*Rsf�$I/s1����U�,*�9�����7X]�&wP�����3�<�I�i
*�P �'��,GR���эj���Y͒YiI�@q�`4�vQs�!3���@�Y���:*:8j/���9p�����4:H����f�h��xT���H���Y ���]�e�I�Gg̉��iJ��<�hɥ�r�v�B�;U��y��.}���,񜳺 Ԡ�e�ɱ��N+�'�HĦ/̌# ܨ��Q�8� �D') �����>|K���<����Y�^�S�y�߁����ζ��xb B�q�q	��.�	N[�:��v6q�_�`R@�?F������ؾVB�Y�Zsq�*��C��D�P�o�V�P��#F$m��LZE�&�
���ƋN;Y�'V����+�h�e��OM�@�u����P�MԲ�X��Z��^��Z��YM�)w�hw�#̘��H:\'\q�*O�4�����-n���yB��#Li��Hb�v�z��+T�e��in�81ahwZ��s�b�W���$�i2!�9�k-��ڬ`}����u�	�~���4Bo8ŀA�*hk�5�B�O�RQ �L��&��p`�{Ł�d
ڗJT
Y�w��ԑ�fT��hn����u���	�����S����ݽ�{�~��b�����1�5��h��U�a4�cF��p �؜�^J=C����u��n��j�T��{��X]�j���u#	��m��za�6:Wfb�l�E8gƆ�`���?M���H"R�Yـ|%@Ƚ u'��z�&��E]�� �Cމ�;{���5��ʝ\6R
�J�2�q��b�+����7�H�����z�B>��������-d�q R��ҏzx)%��,��;K�<��*]	ҟ��B�P�I&�lu�lÈ�J�賜�Mz���aV�N�ʭACU�_�eK�s�!X2�؏Bɗ������R�Wo��CzN��ni��r`�Kd�����z/سX��^�M;ދ�m�eC�r��z �Ǭv²�`YR�"w�z�F������T=�J�yQrw��D� 8L�)F+/�'�۲G$P*�ǅ��jG}9�|��B\��i��ǭS���y8���e&��8k��������_���v�z�f����4�a���PD�����J�ʰFa�*6$�)
�Kf:N$D�BI�g�������!Q(�^��*+Z�j#q`*g��NAb� St�B���ull�aee%rk���Ɋ��c�@��8o��&�0Z�u�y}�Nj�,�N�k�~�Ә|��M�;�l�]�9�Ұ%�����%'t�RV��"����	z�� �}��J��r1�Ri��f�ZQs�G��w�:�/S���r��J��u��rcF-�v�ԐsUBV3����Ō��R���qn�b4�j��8��/���eܼ��ݼ���G���n����O~}w���U�����p�Yڢ�k��^Y�Ypn�%OS�
N�۝S<|t��3T�%�j54�+6�AR�	��m&��π��#� ljh�r�\�������
�>I��|v���q9��h�Ԏ2��,���1%s��l��e�JU�S� ǋL��t9W�s������(_�$U�VC|�U<�,���{x�e�@t�)��r��<�=�@�eM�G�:�2��݅�$�2�"�r�<���r*sz�L�������F����?Ke��ϗ#H�n��K�_YS%���3��T�P�k����y��K�� ���ey�ʫ�X`d�ke�ý���s��$x>K�t]�{�x�t�Hڏ);�qS�~	|ʽ�	Z�9��T:�c�3Y�T�b�����K�	��P�f����1\��� [��#�u2�؜���#�'{������	Yn&�w!��5�}6���)��>n�k���*�K�e*����LF�\���O�b��t��Ҫ��Q�o4����K�	ph�g�}�A�Fa�rFK86PM<G�7�Y��D�5ә2���%{�En�U���Ge�z�Z�bI߳\��ރ����`H��yR̆����3VǤ���Ãm_{�|����5���{�n��]	+�$�@�K�14#�p���.����!N[�zr��~���ؓ΢X G5I����C��a:'+`]%}:Z��N�G�'h��8mw0Z(i�{@N��+Yi\p�Z���U�<P�NQ+P�Ш6py�n^{�?�q���;��~�$ ����g��ݟ�~��.bf��/��Ii9�3�<��N��?C�z6�������s6��&�Y�X�W�qJDR�1*����և�Ո'A�i�}8��l<dC��an�X�u*�f�C��6	���*V��LG�d<V��,�ZtaR����������k� ������aφ��e0Ҋ	eQ-��̍n�a�q�Z��hAZKF�e�*ق� �9{�c�#:[��l�@A������ۖ}ܥl�VS�%y�^�M9��>���)İe��\��\je�;��O��lA�,#0Og����"��S����9�U��r���!:�)3�v���BƜd����Y����d��]��<H,}<�ә�]/���=��%���$�:���*H�:g�*1�L��C��,[^��?W/����q?7�����J �SXVnԚ�q�L.T/1�������!N����q����1�m 59]��|���<>�B	�:�M2bnk�7Ѩ4A��q�"�}�XW����o��V�36i}��o����3�&f3�)���JC��k#h�}\����W�"g�0⊰�hx��gNB�>�Ԁl��E何��r��?(�#R�(0�]d�u�k��i������4S�c���Vy�\�(��v�aϰs��F��:��XLȩ0D96�b:��;��h_�(U�`�>x�Y�<>ii4��lQ:�c�uzj�Y�A��@��]�\!S/�Y�)UeP���b������������������0�{�?|�;���������K��p	�(��d�b�� C�	�6���(AJ��d�f3=0eߖ�R:7C�Z�ɯ��e��ۚA�	�A��eZ�A����̈s�8G2A�KC�0F��76�X̸Y��2N����_���a10s���F�ҵMn�@�a����ٌ0+q���׮Lq����'�Wϐé��)�5�Ȗ0"Yȴ+�[n�(WWn�y8ϼ�٤�[���!C��V ��eF��2�Ġ����˷N^!��P��R�e��/���������Dl��z6e�7��B�Uk��.��Ѹ��9����i��5�d?����{��p(��x��0p��+��T�����޲V�� s��^�_�K�I4q�~�c�˅�l�����*�Y@�
+�{-{�~�� ���X�ú��Lg���"�ё�)0&^!*Tqt�B��G�l�no��w�xtP�k����Y\^�q�F��@�4l�kh6�dG���E����x�|o���g-nbN;��A���;Ax��'Lgt���G�%f�%oo�8w�Yol\B�VQ&K*D�����[��@���X��;R�Vh?,�� ��/G�A��{�+*��2����ϟ���O(����lo:0R�)e�<6���q�� ���fŎɎ�Zr�����g�[�u��/<�����)&�,&���Iv�0���v�LB.���%���0�N��w���S��b���X�aց{���ɘ�
*E�@�Ȝ���n^��_<s���������=If��I�c�ׯ����}��Ȗ�҅���|)�U)`:�j@��9��z�!�mHDGK�S:5��#�8�����cڗEyuY����f�7����VV2��Z�&E@��k� V�li}��sr�t�ζ��B��(p�Ҏq��2_�\}��亖�lb�!�=�,6W#ܸ㥏qiu��2�]d	~�9�|�&�"�I��.��A����	��q�f��/�������θ��2�Þ�tH�'O3(i�%%��YF���`��H��3c��n@I� ?/3Z�gk�Fi���\�gg��.
��Yy|�R+I������'NZ��N�<^���{�|&zr�[�i�g@=;���8bڪ4L�u�TJ���m�e���,3����Eg˹v��|��M����K��g��#�]�t�A�͔�(#��������e�����NO3�u��'GU�r@TR�����Ե&nޠ-�#eT�-j�W�ה��s��'?_�#2��"e�b�&J7�eKA�Ơ#ʮ�(�v&��t���B�l�Zu�ƪ�ttd ���²j��3,"wx��C�����ZPz�%��Y0���ԿB@?%Ebp��w5��[���["?ɲ��9���A���{]t��f�{���2Ý��8�sv�^��~G���:�pL	?����P�>C�-�樔�ܺ�(.�|�G?8<��I�YFζKy?�I��r��X��j��8�C�P@�^�J����]��>������Ƒ~��~$�vg�������΃�>�7�c�<V%������(�94�0�{z��)i�3LQwӧ% J\�2�*P�Q��S�T�
�=��H�KեQ��W9�d#�H��}A�%Pē��r?��,Ȱk�#���q�8p��<"qs��M� ��(<�&cM!.�n�Z��Ic���f���nl�a�y�(�Qv��8#�:[��F&���B@�|z��a�ed�|�w+�?`����$�*#���������q؈��im٪w�r`�)lY�;7��q��H���b<�YQ_�I=+��;�@e�HB��ن��n�8�;V$< X�D����3t0S*#�2�Mz�s.��j9�`�L�PT��8��gk�v�L�z~���=���>�z�X�jX$���L���i*m�����,4����5�Ld&��4ְҔ�

������f���;�:�=*a�b��a��^,����sU�
Cą�FCrY�r��V��E`220[B�G�N,Z�G6"܆ �)O��HZ�|l�xO(vOA�ry���u#�GOb�6��@L
�pV� _g$�0YP���7����e���Y�kɜ����z�^O|n쳪lD�e�DGK�Ri9��.A[�<�V���9k�J 2�
$)�
s����= o´�ɸ�~�x�����6��[O�5G�Y�RA�_�b]S�vgݞ��z�!��	r̆9��"l���c㜮�ʪ.V%4��f?�}�{�ŏ��Ɓ�6��H��ǧ/��ǿ���N��N�=�[p�I�x2TI�D�����	ƃ�~NRn7�\h�~W�>w�e�M����$�� ��m���K��v�@#b��@|���ͅ`5i�l���Ǽ�DI�
y���]�x�jF�E ���v��8G����Δs��)gG�e�Z���d֓Ǯ7W��C�00����k�u|��>��}e�Ji��JQ^��3�WvB�%i�bC*;��oTuX6�sIҴ������#,Vt�}��9�Y��LE�k�4��x�v�5wr��8��D�����7 ��t�[�2' �z�6o�Ќ)7��o�ˡrp��x���1~%�r$�^��Z���9���tI	�� �zj��7�;[3| �cAy��|
�5>e�w.�@�����5���`'��t���b �\Ҡ�&����%Wr(x� Y6f�ZC�C�}�{�l��s����a N�>�^��}��[��8�ԯ��2���Ox�����k(���7
(�9�C�ӽ^YYQ��2Kn^���l� L�gزt�h2K%B��w�}c8&�$��e�9w�-�R�����s䣚����Q�eւ��l���֟����hc�/�?��,�vr�g<�y�d�ݫ^����$�3ߓ^���Ih ���A
�<S{L�t���^�����Dt����
��o�C�I��u)R:��� G֌�`��N6}�z]����.��3�e�k]���Y [V6�����YW�Ҍ҆S�c��F2-& ��ҕ�RG&"1����R(��J��K++Xm���/|�s��o�H?�{?g{��3����ko�?��=�L"�G�E0N���дD��g=sS�zG����3{%��dB�b���a ���e�+W9�^Pc>�����J,�2%!��K��(�Ӗe-F�z���+2F�)Z��Q�ZȊ;]Ε���tiVFd�ǅ���*�)� 	�L�V(��+�C���*�"b6�c��m� o_ZǍ+<}m���6N�ŁDJ��(�i����,��<G�T0��^.��N�v������専���Z7H�Q�E*.��Q�I�rH> �*
��t�,�̟�]b���I�I�i&�U��'a�3�Л���H�C�%�`+�:]�!����gRZ��
�K,'����rps��-�'���~���iD%���ʟ��L[KQQ�+-����$)#����ce ���g%�0O��<_��ƊԔu6�@��&�o�Y�y{���총/u�q�� �F��ρ���˱J�!NB�������Q�'��z�'1ƙU̙M�gsM�g�ެ�3����fFΖ��"z	�"S�`�v&N
v��U����8�=f@��5�1E����e�<G��,�|��B�����re]���m�|IY9�'+Grt��|@���z��������vA�=m�ns%��'b��7K�Sjz,�� �;���F���_��i�38GqV���	�Y��N�±(�i�0mTψ*�=�[�    IDATJ��"'6���n�'���'�4�D�ʬ8��VT�G��6�Ci6�Y\��c�jq��6�X<�&�Z�N�P)R����f�+���s����a�o��پ���?z���{����(`2���2՟٤'J~�j<�b��>&1��\<50E�%��6��x�ٛ�������j�`)��h�C����'�&&�ǇM�:#n���gy�R��O,��C&��6-�T|�������H��A�Md|s������q�T�:�P
�&-Wjr�\@f�á@a�B�˫븲Q���������^�����"�Ƙ����*'!(h�>�]���(dfGc:S�n9:�d�	�[Z�%�Oi�_�3��Fu�@����s`Y��gb0��vCN��2�bjrd\�ee}�� ��A{;�����y3��(O��C�<5�$�u@ԇg�c��ݟ�����Bm�i�Dٹ�r��Ξ1�'�q�����B���������2�q��j����:��� �X�<{Q�`�H��R�y҅s���
���!-�Xて�e�$U���+������'���iV�T�6�-��3ԓ&BfQ��Qwn?��v�Dh��@q�|	�8"H���U���n���*j���
%�=3[�C($o�3�J���y^>*��Z�|贉����R��2(�TYG�q��&r��ا�\	��x���-p�;1^�k0ل���4�fp����-)H4l���K��21%��8��,Gd��}Zw�b�QW6W�@^r�֯�ߨ�<'/}B	�)-�����#�z�#%El!�*���gݎ�
�=@����DG�����ϊ�9�u>�r���g:ߓVm�!J���vS�"/��V+X�ױ���?������o�H?�{?g{����_�������{x먏ք�k���!���q�W˸Ԉ�,-���a4h��n�X�i�.��~oI
��/�c�V��>�	��d��Ɏ����(����)ʠ��,���K�;F�F�=U����|}G���[L������zJ�%4�����}F�y�9,ohR��ط��f�iL(I)�z�Z�`���Q,�1�R�%L�D��j�Kk�yu��Y�Y�csu��f��k+edsj0p�39X����*�x�0�\�ע^�}x����19����D�F���̞Bf�k3J@�Iʻ6���z�rp�Dl^�f3�@Wt�ޭ��F�(t�!($��>��e��MPV0|է�Ηp�8�w��V�a�Q`�Z�P^:��T��o)��O8f`�Ѭ�䲵{F%� &[*M%�ʔD��dU��x��)U��Ϯ���3=U�f\�T�v�!3J��e���s&����Q8�K�*K4z W�'�xZg]��Y����{{x��;88�_G�WD���Lc�>&�
�,����/}�&�{f�JNڸt<\K_� 2����3:�)�I:T3��s�wF,9PJ=^� �I���r�2��+(�ԧeOzJ�ҜU��]�b&��e`�+w��:��3Do��XZsb�;_�_:3U&�'�
'���A�<g}�mc�A�JjX�,��8˜?n�9:[�Fi��崅z3���̤�`0��TAɋ�-�+�l���͑x���<��G<هg���2�̿�Ћ�]N�%d�k����;��Y�<%J�ܔjZ<��)A��%��j����_�����@��|$�����������o�����)�Ԉ�9�gT|����f�� �ޱD��� ��7�u�!i��e�ʛ�Fʳ�>���zd,��֭[x��`�\�6�G�@r����P�65�(jP���Ys��N�h����:^x���q�����Ν;8=i˹s3#b��3�ld�#+	�5���u��K��9>rǅ&�f
�{R\26�r��}j����.��#���]�5��ZE��h�J��,��T%7��!�!|/�k���0	�~��'�':��)A����_xy�ь�9a�Dd�"K�ء.�*�|�=B�(p�v'�!�I�i���qQ�5>��@��L� �M���;�E�e��f��e}GԦ�=�4gz�k�糼+��w���"�3�'s���
�%��]XV�4���2�D.gP�*,�ӥ�Kg�j�2��lq� ��N�������,����6n^N&B�~7��ߌ&3�Zm��j�pz<�ݻO����Y��H0_��,��h~�٨��"��W6��?x����KY	���6QuM�G��>� �vYFv�E�%��NXa��A�A�/�A�e,(|Pj�^��biq��-�D�]��Ü<����t�8" ҀY�.���}>/�F��|��s����dRB�K���{��/;�&�B�Ytꔶ��)Iuk�����e�C�at��Kd�����ၥ���Tl�k����� " +�p��i��(k��{x��F�>*e:�1�+5�E۳+��h$>cz�	���p��$FA��\��@gШ��lo^���{����8��ޏ�پ���������ͻx�`��a�Ĳ4C�¨��F��?�2^~q��t���P/U�nw���vvw��Uz`^ڬs@<F���^�SO]C�\[T��o����}(��llhd���u�	3'�7�����9�Yr����@s�:;�I��9z��{��Z/���^��&�?:�ݻ�Տe�G���ֳ(_����5Ǎ79�ϣX�����'�8= �'@�dI��U9�Gؼ�ĕ��Կ�M��0�b�����R$��J��h�:��x�h/�<����27��<��L;��e(��5F)O	����(�qh{�2�g+�]#`gCJfwM�]=�ؐ��rP�;n�+���e�t�d)�̨��u(^�����ud�k��h���-)�' (/�eM�_3<�lϕVS�67�ު�lC_��6��>�H�R��A��ɽ�{Lr2�V^̡��534=��%J�����*����s������z6��ʮ�f���4�B���
��K��@>>�H���5��QO�_:�|��liqm�q�����Y�K�������<+���+��E�R�l4Цx.&Vbϋ*�9����`:��I����%��+h46P��i�n8�j/j�P��fH4G�9^+�?c������� ��+`<ȩ�r(�9��}%�x��.ՐX���}��Lw�����Vה}$�P���tz�ޝe�R�g͜��C�IV0���-��D���%������$�R�����g1$�Q��ް'�X��m�`���l�u�hVEfė��x�A��S�O��c�KZl�Ř�~�m�|�8�r�2r�e��sϿ��k���?��m��8����ū?z��y��	�۝�51pDo�E.?�t��Z��?}��Oc�z��Ѯf�j�:����������.��{�iq���ի(�8k���XB�e���89>�/���-�1frظr�o���Ǐ���#eׯo�(Q,�?c����ZD�z��{ʐ��.�Yk�Ν�8k�*�V�x��簽}U���X���;s�\�M4�eo��IC6�k׮���>��O������^{�<|�G�?d�D*�S����V�)z�M_:p4��9���}�=~��x&:��W�������&��q�� ��}U�xnV�M��m��\`#
� 9�ŧ�f��v(#S��zxևS92�2�9�DG���șݨ�V������M����a-:��}{3��¶ ��s�Ҡ5�ɞ�p02U$��/����1c0#�e�� *,��=F��#:y��^&N����GS��
X˳E���eI6��m$�ˑ;���-1L��73rt&"
�q��_��x�˖�R2ή�_V:���r@�:B��]^�$���D��0]`4!���#�#i�x�g]DQb�(=�\��|e�Q�EK�j�!�,��/<�o��i�(FϾ��zC�_�-�Yd�-�3��t��5B�1��\�V���f�Q�_B�ZGT�	]M��t�eb,RR�TyD��T�k��r�cF$��>7����i��)�
�_ΡrfWU�@N""��v��"����*wt���.��A����c�Ȇ�=�0%"�,gۏ/:������QN3�0$%��̎��sf�8cE���(��-��U�JE��7-ǭ�Nq|x�v� Q<E��Ө��C8ڤN�o���_����)u:�P:�E�ĳs1�Q%m���Z�q��2D~��_��}���_��G���޾s��G��L�h��P*Q������'_}��ۘt��c���޿}�w���l����*�z�TJe	sq�]�s��I�~�<x�H�C��p����W��
b��/~�Ew�ꖌ3L�\o<���.Wǧ'x��7ԛ}�������צl6���K�#&����{{���=Po�Fq&���Ej�1��d{11�R9������/p��U�<9�~�S���=,P���}��oVpu{S8�ɣ>K�]�<z���=D�66����� b2��9Dv���(��<#�P��t�&b ��{�5��e�9d�nP,C1�oe�*UF���A0��7Gʾ�=M�L�J:/�w�<�dbۦ�Bp���m؝	4��e���F�qC��p
`�&3������{H����/��'��,��<T�qΛc��zԲK݇@�`M�d����J��m�$�cZe ��4/�0X�7�E4��G]E�+ lx�NE���E�MP�>����G���u���.G�Z�rV���}y���n�U��3�����������"��q-Q�՛��*������-��KI�9�*1>����?�VW��L��dmM�-� WI=�� �7�����7ZA\���c�X��m�Z�i�j�m]e"ą2&�Fc����H�{�|���f����[о~?=�U)���͚s%�b���De%餲���~�L�w{�.6�5�Q����p�+��]
%2�� ��`b�|�����)�:�u���u���т��Z*T��372�e�5�u6!Wvg���!�2����u�4V� �d�cQG���>)>ɪV�Dik�F��+R�Zk4����3������p��}��������go�>Ļ;}��s�R � ^����O�����E�+��<��ɓ'x����d��2�f���5*f�(�9>>���*�,FG'��u�ޭ۸}����I��?�c9ٿy���C��W^yE��Q���<+g��K�Ң���9į�+���7�|]�Z�F���˸z}���:.����}CZ�Y���{}$��&W372K�,3�z���O��׾�;��{��~���I�H�z	�B�Qʇ���ԍ+"�2n��'x���p�X��O�̨u�N�ݣ}���D��z��[JS�>�/�a�K!PL�s^�b�"g�Ҳ��2w��?MC!A���ލ���(�X4va֗NP1+ka��c��@���l׌��i![t�$��1t�U�h���_��c���P\��F�!J����GC��d�r��Qǜj 
���dɹL�w�̞x�%�l'gá�=�����!^���esx=�ʄ��4�d�-P�1)3f4��@�B�pQ� �#E?�a���p�KG��'S�"�4���ҢH޷K�.s���T`�ʘSg?��G�)l�����������"�"�z�Zo��/?���y��^àҨT�=g�G��q����5�Ŧ�Ȇ$�7d��Z$�����UԪ�!*�Z5BA�ˆ<M���_3��*��̚�����+
����Iu��ܶ���%�*ڰ`Ъj̈́�?��Y�N[�����rݔ���03st�,�B�F�H�`� eEJ{H����,�z�سm��qy^�c�,l�H��a�l��5BD�
���&�G�;���w���(�^V�

nX3\�"F��@����=V'J%��Y����W�������}���ٛ�q�p����l$��i)?�F���O� _y��KD(+3쏺�H<�����J��V��QYҞq�Q��S��w��;�h��X����g?����_��^G��o�ڍ�x�hG�������.���/�c�����W���o���ܾw[�Q!����x��gqrr,g{��9[�OG4`@vn�NZ9��L�92f��r�����O��?���	�ſ�k����;`��E���|�޸�f���u<}c�(�ɨ3���prL*n�2
$수9�73ǰϬ�����fC�:�R:"��t<��\�Z��#%���:�t���	����-hi\w�B���(\<"݋��J���$		LE.�.g�N9?c8	�v|�CT˕��d`%/�-6
?��q�t�2��W(ǥs�l?]'K`*��5��U� ,o��8g쥼ev�m(պAU����|��Y�P�1����IK� ��X�M�@������+�|�=�T7���xLw6r��OC�[�{h>�\�,y���rm˺��;����e~N}J��3x3l{�=�g K�yN��d�1���&����pi���^��Z����ٔrF6C������TF�{!g-.�����
Z��kX_	���2�d��k��R����Y��G�\�y�´dQ����V�b	L2lCҖ1P���W����=��5GmN7���$KG��l��zm��Mmi�`Ӄ:�Jt_,hЋZ����ن��}c�t���yx�����Þ�#@�b�eƯA�B+���g)|����r9[�a2p"9_Zˋ)�����5�=�,g������{� �����}��o3=�
��E\L-CY�([����qYI%�8�+UV*^RIU�$Ne���I�r)�ٲESA��f�`���g���w�o�����n&�`�
���U�A�t���������<�sҹ�H��X���~ﵗ?�SF�}b��W���o����@���ݷ�.���������J�e_���ګN[	�ci��zC,
���t�Q�e�X�R��׬Ď�P���IN�a��{c���޵�/�U0B9���9���[
�T.��G�s�>�n�N���g��o��o��~�fgg�_������ا�{o�cw�ݱS�l��!���c��7o�������I0�����Ӣ��)y��I����_�d*g��7�����%ku��Ul��K��mj�l+�Sv�Ȓ2	��:�ww�l�L[6SL��4�鷺e����]�6wlñ��7*8�dPe*kA��S:A	�Gc�Q���`�^����y��9�S�� #7V�1#ָ��X�pq�@K��%�0f�Z܂r]��{�+"ye�6d^��'��Z�Zb�'�/�V�3��aL���ܽ&����m2a..gB��`�|dU�T�2Up���=_*r�O�o$�D(���:4W9������xS��p��i�pBNك�I
4��Qq��E�C�G��\���~��`�C���iDb?���>����1��Nt���A��xl�|Q�6�7Hz���࿑'1��EFl~�l���6�����?e�O,���}���	�}�瓴���'vt�ת\ޔ�x`fϊ�M�7IX��b���h��B��#p�c?��A���(��������;Be����q��1v.�C�3�&��|Z�r�"��F�����b'[��W��j6uO�j}]�8�h���8�VELB*�O�����5���=ĕLog�h�wX^A��=)�����;
��ڎm�<�Q��*�TN�� �:r���-�Oz��BA����nAv���M����d2�3g�~������_�`���k��7߾�_�w��xܵV�oZF��T�'F��_x�^8w�ғ�3�4�^��� ڶ�Hة욑��9��m�gMd��ݡ������.�pic<�\�`����+��ĉ�v��	�s��{p�N�>m/<�������>uV���_��UJe{������w���t��_z�;s�z#���v�[Όs�-Bf�@���'ψ(Ł�I(����w���j�N�����������hR�Q2g�Q��U�+�
�l�^�RW�@Tջ��\Z�X�A7�7�>$�r���kq�    IDAT�l:|��ǵ�.Ds�AĄ!�U����u�͡�~0���h� ��Q��D8,Ja��a/��`��L�(⡭�9q?j*1��bZ�_����A��j���s�~I"�l�6lAK*��tLo�� ���]���q��J ��)"O������6�X�A�w��i�#����6�D;�׎}�X�������2�F�����;N0�2wB�C����.ҵ��m�U쉇�O���zP�����T����Q����e���u��FJ9jLD˚�5�{��A��g���O�b����sG�㯽`�چu{u�= &R�O��MH$��|6'#�Q��
R���k�SSv��6;D���a��m�RC����e��'��)c%�	I�!פ��;2ŵ+�@�]�]�]���?)+�K�}#7�̔�`�wyaQI)��GܯT����M�
s�C!~�H2��g&�d2LC�$m��� �JN!�|ʙ��RV�V�(e�n�ꭦ��?��چ|�I�%�g)g�F4N�V�)�Ř��ޤ���1i�|�2ɒ�se�����{��/|X���U��\���������
��4~��Ⱦ7��-;��������©��VHO[�2ŠJ�K φ`�^C=Hئ�T��ʚs���eZ޵w�}�޽x�u�af��¢���Gu���~]��ڴ�� 6@ɿ�2���W^�{kwU�@z��U[ZX��'O��|����L�L���?+F3_�nݺ%���ZC�toa`��S�U&^-b:�Z.��?���d?�S���/��?���o[2S�I�dM,�����|֖���ȡE�*��`C�Qk��]��b�t9����?@'�RֲɁu�;d���UR�R.�]��� �/�vسy��4���]�?5FC���0�:�wI~Ae����g|cƯ�U���p8R�8L��/ė�{c;,�$�Ø�����w��f��K0i�uգ���A���M��:�̧�y%��R9L
�Ѓ�6T�(Z��EH�:�Ej|��k�!��TӅTV}��:�׉�|�j��*��(�g�}�21���\�#�����^|�2x�}��FD��x��Q����҈$�d!#����+1^�]��ٜ�e��
�Q����;;]��9cn��L�~�K?��ۭm���~S�Lth��=$)e���>�0��[vq
7��5�c��?m���	�Tr��!���l#����= �:Ɍt�q�`H@�`_�?X9���>{�ׁr{A,&7I�.�B&U�0��9*i�eT��5�ܰ\(�;��=�k{Lu��Tqo��:�������g�����m\�{~.Ȧ���;g�ÿ�3w0�[�TT1�9�ڽ5�p�C��qN��9!�屘�gyb��633��}g���Q ��23L��>}��gN�������[�߹��_��a��ִ����Q�z����ZJ����Kl�]˧��9�Ж�b�Ϟ,9��-l��6��#Ű��ٗ���\�f��\����+U;|��fM޼y�6w6�̙3:	�de����g�	:^����flan^�K̴
�4.<mǏ\{��}��-��݄����� �Pu-�2y6F*a곟�����d���}����߰La�R٪5��G&} ��c�Kv��6�����#?z\��|��{!�QJ/��׷�uU	��g���.k��z�g�&��K�3s��yTS�3�8?���I�[�|��1��Ze���a�R����G�.�'yMj��v�� =OVLɀ�x0ƀϟ<3�=V���Cf�G�Y���H<bU���VE�7o:m����������I�=�ZpR��,U�!cU@���Q�H{e����r<�� ����v��AE8������OL]��C�1N�r�]����������H��U�M�}�q$p�X�)O�AO��G` �&؊I��X��X���-��7��Ԡ߶����8�d�o\��`�𕟵�_Q�c΍�1�+/خl'"�龫�8{>Ĝ�`�p�i�̌;y�fgf,���������x���`�P�#���:�8��@]��ε)i
�]�r�b��'T��>�ش�bA�5<�YC�p�����R�a��;$�J�۸"�]|8�1�<�DGÒ�Jx���דN76	�Y|F�V+�拗.٣�G��n^��!�(E	�	����e�.e��y�HyX),����o���+��h��|�o����o�w�?��[���˷7��N�v�)k�K�u��)�g��pפ$�X���ĝ���ʤOSo�(�aD�������i�����׃��o�#��EevL[[�x�lr*��t��j��&k� /�u�G�^x�Ο?�E��[���;�`?��&c�1(S<2z �&�<����c���}�����Y:?#�?J[��	�_�N_�����<!��m�lskW�U\�苑)�;�֪=��-��l�b�B^��*˰IaT���j�`eA�wݩ�T���<�88 ����l$�p(��%B�ܛ��$�����X��I+�b�D�(�sƾ��Zá�6��W�*&��� 5�p�%��@��+�x�E(�u"�[��y�7��v��9u��I�����ߓ/�C�C���5����'^O�<b�+��ˋ�}�>&*
p�u�]��9h��Y�Ѭ���AO:[��?��K���`��R{�K h	R�bŊf���+���?�1��G��1�;I- ��@d!� c�AOi�f*��8mwn\�^�f/=������Y=$UC�߶tfk[%d�+��G0�qs?pz�|�ɉ7y*m��o�n{l���C�<��B�I^	˧�=!K�Ӛ��ɓWv��-?5���.��X�D6�|��,{@�wi��J���x��9� [�l9w��k�����	"����*�=��=�p?�OHb��`���H�u�-��i��U
T������c8k��\�L=|�n�������0���c X)y�-��
}�c>#ݯ�%�JM��ꊝ<U������|��W!�P��~=�`���n���o�޿�e���V$��^���Fu;�b����=w氲�䐩>�J���'�8\�j�l�^!�jҳ\���lu���˪lY\�:��>L�~�c���+�g`=U�L$�P�abᐴg���믿*(�$`����,"2�t�.zAf�r��p�d͘q{�����v��i[���6jmK�V�0i�((��S-�ԉCvheF�	���v:��hǺ��l�
��؜b���jm���n�l�R���%�����{$���\���;�u����2Vo6DF��QWkޣ��Q�m��'%�P6l��!|ps$,��X!� �:y�����I�R���^3@��s4ҍSB�����X�/��ZA�ʡ'V�1Hg��]�$Y�y�{m�lB/-���0@[���{x�S掕�-�{�<@w��%Vl׉l1���� ~�H,�	�'?=bn�}B^���}�^���˩�WE��8`��V�+�0L=�43�1
09��k(���X���:�'����5{p���ZF	I�,�vΘ�	2�dE�r`й��U+y{��f�VM�����h��̧�.��][GDO>��丞[�d�$�-�CZ7���}o}�666?�dG���CV�m4�B&�'w��ېhr�0k#�㉶��B(B[$Vi������`囱��{8)�-_,X&�Q�FҚ��9O��yMf]�T��oi����8ΌliaFxġ/1эg]$��^����Ao�\���C�H�?T��Z~J��`bY�]���¡-���m����ݽ+i��҂%�}磊����1�q]�c�v��pW@)R���O/�{h�ЗΞ={�C���şH����_�o���`{�1�� i��I77������C	�3_��=}bɒ�'Jbr�9�T
ZItqP�@S M��l��ҥK�(�"��jX�5T�޸uG�,X�ׁ�΂�Й4�� �����Ci.���cP@�{��Yk4�ʎ�_~�*4V&ȑ��v` N�/3p�'�Um�-,��Ҋ5�#{���P��Zk��RF����,������nwF��g��"���U�>X��}k�nJ��<?gGW�X�\RFO��g��\��ox���<��� �S�����a�x0�]�f�S$7�g�7a<`�^��i�u�g'f㘿Lش�c�%h3�l�51Ľ�����޻������d�R��N�?��}v���D�L08X�F�hd�D�����z��o><ȖV0@�!`��M�<�"��+,��c�0�������ݶ�*�ؓ��?��x�.|}��뒡�����d���sFIm��L�[�[LaT�g��[ujZ�&�z�$\�Z͆MU�V̦��ز�w�A?{ꤱ?_|�EkvZVkl��J����������*Ri�����d�/�Yyj�r��5�{�pS����?rԎ�Qk�Z�(ؒ�RY�4F":�σ��<ERԁ^�Z	*c�&�W��P�b�ޓ��82�I��\�Q��nO6��o��nmmk?�\D���ft~��h��znT�Zo���`�����O|]�P�g��#��Ϣ�ù��뽕�3V��}`}�h�µ�G�)C�|^�?��Ġ�v�Ţ�&��.�\ϼ�����"g���[��˿x�#�g?�@�{<�`�'�]������`{�!#�2�Ǵ�6W2;�<��|�5{��!�7��#��)�R��[�e݃W<��U�j��v���T	[[5k�[v��=�}k��=z:��������W"2F`k��B��i�GJ&�,ꕏ�$w)�kknI��C�T�gtP3	hw��E�bG?��U� ��_\���kuG���["S�Bu�{��ǝ�&��ꂭ��Z!;��d��	��ng`�|E�ݝݖmmo�u湇c��|h���dLF�K9|Ȫe��Fq��t�������U���zh;�X'VT��a��j��ڐ�p���M�3;��1P�j����H�=�ZA%�o01����� ������\{>k� "��bY{$��$�q,B�^	f��=Ә0Ġ�F�������t�v#�$1��$�أ��6�� _�*�|����Ī �H���/&� �D �F�� | 6�5���P(��}��5�J���=�g�uD��w���+&>�F��K{���xkӮ_�n��F�Ӑ	v���[� B�>>	p�Ӗx)�����Ma�){ȗ_|Ѿ�s?gK+˶��@���Oo~��q��\�PG��: �`y&������̊Y�5k�%*�Jv��I;��ls��4�s O�^��پ��-Η��g��D�H�����h	j��۰�)O�H´?¨@�X1ܤ?���8^��6[�sOv��VK�H���g���U�C���+��g�ؘ ��,���@��T��*�%���NG&2��Ǡ��5�Jʆ.7"(߽�>~dk���fϕ���u�nZ�T�b���O�)�$	,���$����W������[?�@�ă핵m��e�T�:��n0��Lad�F�g����1���6�:�4W �a3�)�8�\E'�j�v���r�r(ld�[5Ut���2�Z����0�3`�L��땖&�/Y��݇�������Z>i�6�ٳ�5��#��ې��vaa��SӪ���I ��m�a���dK�ׁ�����[uz^~�T��Q�2�i�����I%�?�h�V笘ǝ�������`�{����:��Ŭ��k�n)�r�!J�8�:w�-��:�>µ(��J^�b�Q�%h�3�"Ǡ���2���5�:�vxq/��=*�?��9|"��(8A��űj��F֨���G|DbT!&���a���Ǥ�/�f�B�˚��~pί_o�����`Z?k$������2�."�����Ҍ�2�?����ȃ'~|q}��c���(�R2���:���C��rܫ`c+�I���7�q�!`sߣ�T��8�%&���M��!.�i�=�ݿoW�^U�(g��y� �L֊�ґ�g���L�	��~�!�O:��i���W_�O}��6�0/�؝�{�?��=m�b���g����\A�%������p��v�i��Kv��I;��j%zʖR�H�����`m���J�5��Q����EdwSuh�	ߣCc��@l��
�B{Fc�ܪK&���i7o|�j~f�j�<uޞ{��.�#߻��؆ *4��I܃��xvƶP0�eN���=�����(���蠚 :��������P��6lo�X�qB䴂�qξ���"�ægM����4;;��zd�/�?��o�(��o~����[�gW���Vm`�d�:���P�dӎ�������"��7ǚLA�f~~N�%I'�)���677���M[�[i[�]�ĝ���|/M�`g���*M_��؇p-�[A�{���CU=�l����	XL�aa>���6���ꪐ/i!=~�H�i��N!6U������/j�m��W�mt�E�
NV �umv�lǎ΋ U)cٵ>0��iKf�S��i7o��C8���rA:����O1�I�Lر�#�8���Q�9��^.'���j�|������}1���e�٠��ß�I�}��(�����2��b�� ����� �B&pރ{��éPt�(r'���Ý�=K��P�r��Jƥ=��������4����	b����j�����U�b���!�F�j�g,��'�̀��}`Ӄl`��מ�0�>��c ց�u;��~��dB�UX��GE!u�&��0~^I�(�w`89��cA�{w�>���U=���w�*�)����ߙl�R��&cŪ�gOE�v�V���F�����=9u��̗�d��9��ݶw���=�|lI\��0��u�G���vK�xqyI��ν��ܲ�����ö��d�BY.eи@ށ����mA�!�泬;O��&����z���w�&{��I�HmZfT��_�U�c=�f����C�ur]|��Zӕ2֯G�O}�363;�g�~w�O����Vȩ�<�0G9���W~=��p�
�R�Nd4��Z��5[u{���� w�ɸG�A2a�bY���$e�q�-.IA��T:r��bH6�E�,��(��cG���s�>�����o���z��߼��k7���N�4�A��a͎�������3'�-1X�޷��׭�m(�..��<��UO&,���v6��-�ښ5w��MŒf��~���C�cOY����dÁ"$�{z��i�=q}�YA�>�(��I�ހ�_z�e;r���,Zz�o~���훶��X�(g4���Oٹ�>b�A�n�^A
o�d�"��ф)C��*ڑCsvxe�J%|ha{�d��AL"��z�+[�-%r���n�ʶf�T�*��aI�Kv.��@�!��n��ڲ)8%��`�aż�t�*�Iz���C{9�o����W�*He�Q��@Tt1p=����cSFBGtX� �`�n���V�~��Vs�%�K�
��!���UH<�NU�I�6S� ��@�Ht�{��b�P+�x#{�nSN�+h����"��IK�V�,�AS)��d�Pc�͆��I�b�ʚ��Z�hýQR����aEUN�!IU��@�BB	T<W�b%ʽ�{�]w�Jx<������(��~\���Rղ�iKg}��={��iaQ� ;��/`� -S�jfd6c�y�^z���޽tѶk[2��t�%[�*[1_P���[U�eF]NTm�����5�>��V��Ҳ��̪53=5�y��l�L=<8�5]���wD��ВA�lH�;��Ar� �8<�����s�&֧����N�a[�]���fn߻{�vj[�V'�~��?m���'�<0�ѹ�����C����XD�#^G������+�TR�<��8R	�G�}��ln���[T>(���T�b���Ҋ�K%F�����^����wt��_:}��?y����7�{k/�6�Y�#{ ��`ˎ/��W��Oڋ�ؤߵv�k�o����{�h-.ء#��D�?�<����m[�{���]I�Q�[�2m�"N!EY_�"��YN���?��8���_
�&�2;ql�`�%\�����0� )8\uSB    IDAT����ګ�c'O���`d��~�������[�l��UM�2�z��g>k�>���?ڴ?|�-[[߶v?e�T��c<bGr���D�:rh�P� #��O�ZϘ��Y"k����Ff?�lgc�M��R�������Z@���hu|,�ϪV8��)V�� �Q ����&�� �8���8����X`Ǫ/y���4�����}��l�s҃���)��CD�������]�OL8r�"����Ņe�n�*�80��a���������L<�8c����WE��&0�#���.�AAQt���l!���`���zS�1{�y80��v�%��ߣ���YB�3��=f  �!Γ&��c?>[�X���w�u���M
a�,� ���$�~�o�o:L��ͺ��k�:c��9�"�@�l�������%Ƃx{�E�^���i�{v�����S�`�5���H�g��e^á�m5�z��"j��6��G���Rz����L�J�g�D�Z���i ��A�9�G��0���Y&���χZPO��Y�V�m��3�HIh�Ɋ_-a"��͝���߾�f�/_���{����.�s�?����_��v��R����p�8Z�� {�fXGZK`��"_��k/!K��7��w}m������-��	%+�v�s[=nF ��6]�Z)�S,��t����8 ����o]9��=z��'h�X���ۗ��7߹�רl��I�
��ć#�[�Vg{��?���z�%��4Ѭ>���8�t,�0	�WQ��ҧ¬��xd�5s��65p,6e@h��Aİ\T��@Y��6���>I����1\�V�{_k4��	��fC"y*[��矺`���1;{�imt q*����߲K����p��3b~�_��U�u{�~�Ϯ�z`�A������0G}T�l�d���SǗ,���qF���5}KeK6;�l;��	��vw롭ݼd�1R��2)���ʨ��Sٲa8D4-�\
B���$V1�M����i�L7�+[`d�7T$�x��7$_�GCRd��<����{�����4~F#��%LU��6��[=z��=!�k>4�G��C�ɼ����&M��{V���&���:�ث�}8Z'�(��W����E��f�U&ú�􍹥"ר�t�o��I5�[��שC�A,���ѳ��+�|����w$�ʖ׊R�X��~]L~�O$#�V9<6A���#)����{��t_�-a�ٓ	���[6?k�͎�=����w6�Z�٫/�`gN�;7o�;o�����y�ż��	+M���_�t!g�������P�����L��V3g	/��5{-�&�V�45�6m��!��^�+�V�E�s�z�j�u�$C|n��oT}{���=�~
���D�5��
7�)hDb�g�/�������4����ݽ��nܸ��.�	��B"�K���쓟����hw�l������mtO��<�mz��y�h��7�-7(A��L��֦�I|�y'���G�g�f�\iܞ%CBֳr>g3ق�,���҂~�`��ȧ3*�V�����+G����B�I�'l��Ǘ�ַ߹��W���n=e;��u�~���,�G�R��O|�=v�
)Xa�@�l&�N��J�ff�Ef��X��x���8}��e�S�i-�8p��+ڮz1��i����(s�	*���6A*%�Usc����\��g���&|9Y<�wԆ��mu���>{�.\x�ʥ�=~��lr��к=�}%T>�s��+��^���rE���7��]�r�v[#A��I�2iF���Z����Ge��N㊄��o���ݽ�غ��;q�2��M�X1��ڣ��v�ݷE�"�n�����5�/����A�Z��T�����(�gkF*��sP%��
�Ĕ�C/Nԉ�D�mt=R��bc���
�3�e择>��Ͻ�j�{@�%i#�ab����Z�w$�Y1�(<z���^��옍K���i�l�R�D$X�}���Tv�Ģ E�-����LIEGH&�*�#�@����ܧ�Dp���{�Y���F�=&���q��~�W�ܚ?�0p�tI8�h�D8��]*�ו�i���U�eLP�A�R|O��s�͉뙚�վb��o��u;v��mA��ϰ�����s�.L������2�R�Z�^���Y����=��k7���w��1��h�,�Rflϼ�^=j�}z]�޸V�`�I�[�'*>1�y���RC��t]�!dB|�a�'���D�ʹ��Ug�*r�c  �MHl�'��U�3�^��B�4WY��=��m��O#"AJjB�%H�9�i�Ñ�[m���M�v�=Z`�Ʈݹs˚����g�?e��˿,�����E����NV����D��38܀��������l�ްF�m[;:+�`$&ZŊ�8'x=��D�t�JՊ��=I��s;�0kǎ��wƒ��s%[Y\�;O?u�ןt����D�?���տ������յ{4��V�i3x��Dv�j6;5��^<m�N,��BE��n�=�kk����gQL�C#`��,���$�e�m��!�`��@ءgCF�fCP9`8J�L�PtU�r&	'>=�DR�=�w��l�C}����|ѹ~��737g�Ν��Y-�Ǐ��>�=��yk6�v��5�u�ɳO?c/�����]���}�w�f��ܲZch�f�Sk�բ92c��,[*ճ4�і�F�gw�lص��ҡV���3p���:m�w�Z-�fX�i�*����U1w�w�Te5tBA\SR&d�x��4怇)I����`bg�ҟ!��T��� �M>~h-���y$6���S](�vf\��k�	s_z�$B¤���'����Rff�R�]B���j����o8��q�JW�r�d!t0�@���B�c�D��â�<�=�Ȍa����¡en04��T e�a
j����4��CZ���&�#%�j�	�z�'I�꥙����맇M�_��5����SXY�re��A�p���C��FyL��=>�ɄM��4�/��҃w�zf��p��We�B���iK����}�#0�[M��yl����S����8y�Rɉ=�O�����X3�v�#���Ҳ��-k��_8�a^�����T̻ot�'?e
�r��&Vk5d)� �����$��j<�Lىx����>�e�dd7�<���3�� �zW*^C�oI�DTr	�3���Be鉕��h��F$�lc{�.�Ů\��$�9���;;T�O �){饗�s��\`�;�=�z�d�!�d���4�LNB/˹y���f������?z���о��q��� 5j�S:�r�z]�-��u%�TP/�E"e���./�ҡ%S��\�r����c'?�px������|���~�{��������.�Ë� ױ|�o'���TibS9[��Ȅ��U��[��w���!`�-7�h2���t�V��nl=V%�æ'
�bH�H7���긥��Zg��Pj�*�A>��]Ȕ�ٙ�ݸ����>�{�\Ϊ�'6d8�����wt D�;Hi�d_���ӟ����߻������ZTǏ���'O�%������iwlYw��1Kg
����"�ڑcsv���%R}�Āq��h����{v���V�,X:W�T>m-��[O���]��d����Vg��ʂUI��4bxl���ٽ�vC�\�Q6�L_�P�c" 6�m�ru���}��i�F��ܹ]�����PI����r��J��Z�fkG�:8�\��|'�A�{怞�Vl��#�8� ��^�`_�~�Y�P"D��*�0sU��s���
�C%�"���Qgi �9	��Ӟ�t#��ܺ�4��qd��`�H���EW���
s�4�[޲�
�EK�c'��h�:ҥ�k!�U��Zvku�F�D�7_���&eəZ.i�C��c�ӂ� <�7&8�T��jD�>A"�y!g�@������ݡ5��1��ִ��o+X�j�5J��-�.(q٢���EZײ�wo	R���^��nkw��=UoH�j��@�	�\AA�>!𦯳��O.'���Ug+���5�ʛ�v$n���ƮuC1}Q>��Y'�Y�2L�G�@��Z�R�]��>)�]�
����T*' ��g�m�p���¬�!�!"��J�HbIxR׮ߴw/_�Q�33�h5��5�Y@׬W��x�j=1�[G<��%��n#q�݉j�v�"�a��G���`
k�w��0$�Y�9���0�>�R+���d�$8~�H�]���Y�*H�`����Μ;�����'Z���7/����{��6k=+���8%�`��	��;V�þÿt�qY0��K7e�7��ݱ����S��8p�F�Ł�̏T=�0��[�+��y�hs �0��Ò��IKP�=9qr�l�ZU���ۭo�&J�
V��ּW�H*,�(��*�(�Q��c���}�����i�y���eT`�T�¾w��,�_�E��t�l�~���Q��jq�ؼ�9}Ēi*�l[]�����w��Y�F�/��1�q��%'�mL�j5o�/���MW�J*8ȹg�ۅqvL��C���#�ݑi#�g&Yy���$ӳ��(�U���X�aT�8������y_A���T "�1F+��Bx�t�jZD�r`W����T�d\�*���rĮE�&Y����@F��O���f =� ��aL_	`U�``��G9
�y��G�"YqS�^�G�1p���)_�
?��_>}��5-�D��`˛�ru_���@��'��礲������׎�(���ܔ�A�	"�Vel��V*p�+�M���*eV$kTT{|f=��[
�=r����}$��@�|Ҕ�,��f���l���ʣ��ڮ��]�		�3_��]^�׵v�#�ڤ�D��S�ʅ]+�M����S@���X��qR)Z(A`�Q ���A���U���vxeَ=������h��6��Xg������w����vi�O�±J�M(��vwj>X%eJ.!YNU|��̔�s��c�Es��o_�Y�C����O�*��h�&��.���6w-�Y�X�7�
%�f�//�hߔ�=;��\�=�=���?�1�1�bY�!r:K뜤�}�ܮ�f&h��T�&:�-�skəM;�����܊_=b�٪�o�pl�����~��'����������ƥ����]�+�a����T�q��?0��UW������c*#J��%.@��l�4�~��sH7��ç/�C�PK3�Q&�L�\��J��� �Z�%8Y}�m��!��`�2�$mk5��~,�Ⱥc��\�`y�%eT�NѻYZ�5����d򑻴`���Y�) ��l#R�
L�g��P���V�y->D���ۥ�7���]�f��,i	|��1�4L����i�6�6����t��g+J �Kp�tlT�~(�GMߦ�f�y �$!4xU�j7�Y#��X()Xy���n��y�|���yC���(�6{��w�q��+k<Q ���~�k]С�}����!����,���f�S>ie4K�*� KFr�@� ��YZ����ͦ�VkWlT�Ȋ��̃����%s�զ~��ZQ�,D�81)��X߽~�D�f�\V�K�]y��{}$@�i�u�lԛ���-���\�*@��H(�>v��#/!��!��~ٍVܢ20��+d��=�dq����g�S�V�i~`�l������E����^#��{�іmlcb����8�w�..���C+
�jZu��:ڟ���t��#]������3��*4��-9i��9"����o��򶲰(8Y���6{㾞]��R5�����C{���ֈ�T�3���15R>�ԏ�s���b��|~Ng�����)gS���4,�����|J��V6з�P��4�;iv��1!@��m����Q|T�u6�'��f@�:�@i`	���i����NrB���=7�Y���/]ur�ۚ�'�F�c�Vۓ[, �X��L�b��[.��Um6��ós�~��>"�H���E���sO$�����?�{��/3���ꪲ ��m�Å��.��	�=A�����˃BH�c�@�^�a(�<M�#O=Ad'U�b�b���(i ���d}_L�n`�F�&��x���龰b�3F�9����A���'H�7TY�3��lβ9X����Kf ���Q	{fg�ņv���3n�z`ׯ�Y��.F�}�AJB�\����O~�;�~h���Y�}%'�V��M��:\���W��!Ά����5el8���Hw�L��[��x��(�!�l9bZGK��'YN�R�
L[�#��r�hY 0�����K7���m��b>c�4&�N����?�`�����Yt��q�RzMI��h���jA,r�����3�5�*V��^�c���D��s2a���'{H~`�;A�	<%U�.�+���;���J
p�����I�L�6��5@!bE�\=^�Ψ�rI���D��]��u.��S�KRR�h3��m:�+� ��Xۻ�u%��B�JժJ����c�جi����~��J���qf�m��!�V
�iխ�j��b���/J�:���l)ؓ�Ir�ɮJk�f�k�����-_gM�u7">��e+fsBG--���`�Iڵ�C����*u��=�5�{ɛZ,컄�������PPӗ��҉��ly6�G%���ĳ�=�4͇Y�2U�� Y�~nq� ���@������#���֍[>ްє�Td��lH�|R=l]_���Z��H�HعN��T�"�m6^�D�{�n��l���%�lg"��s�����V�Tu�Ȼ��fmif��?��_�)�m0���"���>�`����{��{�_�*�#'OIGD�ա��X�F�~OU��������S�*;�e���	Ik7��@!�p8��$Ӣ�e�`8Y�z���WÒ��+c�Rs@+��$-���V�
9x���߷�� ������="|,x(��;��Y\e�2��Td���{�=�<S,��[*͡����E[LYB��3r%���쳵�k�oY�� 攪[�3�;կ����{8�ٸ߱\��9�)�f����u%)4�i*H4}���$�BA�Ӭ7�L� Fb���>A�Hd�
�{U` Bp]l�� ET!l�4�7y�	�f�����&�*7���\�n~n��ż������X#��`L%b#����Peq�Il`��FT_^E�+w��$,�O��RЫ�m*3��Jۡxt2O�`5�<�=eM��<�"��lZ#$�]��Ir=8�!��Y����5LĭC�q	��?��̳W�ZZh��!�0m��<���Q��,�s���Q��cu����Ӝ��
��$.�"I�	mk[�8'.\����w���6�$����s9	_ �s�BLܛ{nvʎ=l���6�-ޱ���i���U�S��m�F�n���T����}vtǲy1�����7��e��z�]A�AsE��0+5�
�\F�RZ5�^O08lv���L�Bdu��#\��ӆ�2�F��uT�!	�\#�;��$�d�G�'_�@���oH��z�"�u8g����ͤ��^���Ç�j�|�a��Ku 9�ԆqK�h�������'�@�� �{�uP�BtJ��裘U��4N�oO��@��;�6_�v׶�NSz��;{���;~��W~�ӧ�D4����Ώ>�`�O������W�r�����Z�RQuǆ�d�3�M��J�!ːͳ@�mXWP(�ǖN���C�C�DB~?LXy����ʉ	�XYeЅ�LTfb*�sv�	ik71��lG�d�a�o)���R�H�t	JT]4�y��Q��=��(���9����C�TW8_��^�h��ﱰ ��װC��,�,y$`���ft�M��sX
X�q�>"�o�d1�������sSu���!�ß��U)���wj�8������,!�<�e]GԣrO%��&���Q���S�|��jA���`�;������6T3�!z���� ��i+�T���>Hy@DK�n��`���8����ױ6Ӡ�F6��#���3���u��*wuW    IDATu0\��=$s߸^n�Y���b��둴�b'��Lp;䎆	3LYO��>�iBK���{�^9���YL� ��F�	���g���5�+z�����2n�f|�AJ�����n?H��깅�t���c�<)�C5'�KAZD2�07m����\�z����s��qm�F��A̓)0�L��C�{���;����R�`�;�~h91�]c�$t�>�{��5�r�GtM������T��.�Z���$���Ft�tGr��'籭�T/gT<�^�O{E�s�:Iāq��5���LF&Z�B�d#�Š�����GղT���i;�HOX��B� ����=����K8r"N2�z��e�Xh=s>�C��7	,�8^g�ю%���P��N���'���c�|�?����U�H���o}�y��K�V�k�-�Y�:-W65Y1�b`U�Y�r��@���L��l4�
v�]������ �%&w�Ђ|[5[X�*��F<���u)e��a/��ovA��ɔ�6���aM�Tѐ�4�5۩)��q�	��~e��?F�9��pc�I��=�#Y���>�>���ύƱ�k���X�4%itma��_�1Ax聖��� ;��]gjSM�Y`�BD�9��	�V0�zd�7�M��C �F<3'�j�� ]RM�I "���;�g�?߈8�d'�ZZ�@z�`bA� J@��u���,�H����E��3ބ\���{�di7a���51��$�naN�=����La�j�����1����=~�Q0�94T�f�L0��ꀹ�a�$@M�a��%�D��7G��F�k�i�7���_���k ?D��?)���! qm|I.��`y��������P�!f�M[p��{�t���PG�`s�H�HtGc��%�-��J'$\h���f�6?�&�5�[\�RB��rI��5�H�%TQ �0V�U���=����4�
�9T_���5�-�L���ag�2�=иB����"8
�{7�u^Fd�d!��sQ�҂a�� r'����*Ap���c܂$*��U9��IO֥g�xj[�	&9�ߐ�	FǛϋ�E
I0m4���A!C�`m�`����*�s�������s'-����T�b�Z�㜒�@���$I��[B7ZͶ5�:4�N͇��"Ž�۹����H�S�%;~���=v؞;{�_�ُ?�Å�緞H������__�t�߾��e냢Ya��1� ��u��+n9�F�f+S���5�[��<�����Y��k�|^�X�L�����Q?a�ʈ�J��^Q�Aud�r����*[ld�㨦�ᦝܤ9�T��}�, �hXqp�	��b,��s�U���&5U��L�%�A`�1���]��'��z�P�Y��^���ii?E�̀= lyA�X 	b,X�t����	�͟h�	sW�`����TMI痶!�k�D�%'+y��+�`�nȧ���k\�z�(;w�6����C�󾢻���d�ϣ��)ߴ����͝5�$:ޢд�$9�> $lV�O�G*��\�1�ɡ9���g���ML<y��4ס�{�)V�)�q }b���5���n8�lWJ�`����^j��qq�����	��$4�������Y�� yE�J^#zUs0�9x&]M�+�Ú����{Ŝ0�d��%��~�7����	F�B���V���l��׌z�H���40rb��'�]X���h���Rɫ|���כ-�bYA�c���5�a�߫8�\��s�N4x��@�H�\��,rd)�6����N���s��4��>������H�8�!�����j2��273eG����YU�Zk����sP_��Yg�g'B��(��^��.��I6��z�ꭦ��|��8��I����܃�3�8o #*���zJ�`p��L����yqn���^�CC���hsC���t��iwmg��$	��Bkh��a��pbX"��\i�f�gm~z�NY�������������U�L���o����?���[][kd�c9�����4�P	S42��;��;v��oY6	�a�	����-�ϩ����}e�T�ȉ -�ϊX!�}6K*�@G�&[*Ho�c��v�:��;��ZQ�H���+`�;�H:�0�B=F�GE�BYA��C���pW0����Y��ł�L�myaގ?j�!q�"آ�#JN�\^��$.g�3�633��G�@���/���烉�!s�#D/���	1�6����`qz�sve�*����/	��_X�qs )	I;�4O�!b�7
n�������\IC��~(B�ٗ8���'��p1b˫�ޏ5��7)�d�h�5ل>�_���c����akKstճD��K`b�?��,P���������`�Q�
zX�-<%�D�Ʌ
yQx��88�~��o�n��&������5(磑�f�������>a�x�6ce���D$X_�����U��(�W�� 2����g�����W�zuy�S�T�$`��IrG�N�]��1uSc���mzf�Mdre��=2k�u���{��'XtB{$/w'��I��<U�	�J$�BR�� ��꒿��d�zCd0�I!�j��ѫ.��3�M�ͧ`O+Tg咘�Y뵝!X�A����S;u�Z^�����$ξ����/��"�8�@{0�d"J�-O���܇�v��#kt�J�I��5M22vɒxI�#؝r���'6U��9+�P����<s�H	�B���~wY���#�ᚢw<IS�# �b�{�x�<H�-_����9��������������W������	���ko��w���[͡m�s���	"z`z���M���v�-���ڃ��5�0͹	�t��*x{k�j����$nI�����v��Qg6��Є}��X��~)���nW�ݰ��]����'WD8�<?��ٹg�uz�L�Sz �rذ���t���(/i+K�zxI0u����faaN�_mgWRo����Gv������%�T��p�0���!m�F?�?�*/��C��)�������9�$�@!�8S5hʤ�+	�.돃"d�,��3'�ᰠC΂ft�$Ȯ�95�)7�/��'���s� (! ��`�&���\�|��znX�1S5h��w�J���E�v��B$=���u�xdS
Xrn
p��!�����J8$��$�$Q�@AR��=��L��>\H6�W�4�����~g\�dg2�P�K��ĥG��?'R�V
`�>������B0�*cX���e*�4Տ���C��^Q����+H,��$��<Q➺�����ԚaЂ ���C&��&�Xȫ�1���`�8��	,��r1J����0T�gf�kW���,���{�No�Cd�2�|w�6��֥_���T�.--������]�oHǒ����$�<��}lu��D�n��9+�:���߷�ݚ*�g�yƎ���e����#�Dx4܏��C�s�{G���$+d ��$S¶qcgG�}Y��rY�--*��������y�𦵾���9P���sb-bY���#�(d�j!�@�@Ue���#�dZ|9�q1�ڊ��N3+T1���ű�3�¹����/��cN���^���?����N}�ۃ�5�)�������`�͖
�7���9�do�O&��^k({B7�6W�rwg[�\��Tjb�}ڞ��ia!��=�Mn=��1<�����߲��Ic�h�����
 �`|��Rk`ԅ�W�F���W	�
Dr�S�8}Q>���v��s��	����O�6d�߱;��ڥ�?�������#�b���5,�I�@�T0�NE��H��RE�!&�7�E�;�U�lg�v��E����نb R�O��	 �sE�O�pIXؘ�zE@%�ɸ�G?���أU������c��� j���Lh�轂<��O��`�S��<��VO1�v��lspNak��=�lԳF�}�-�n��&��ԛt�#IA�C(�u��;V�~���z^����|�c��ڧ�B;`��=��9�Q�3P	$>fN�"��/�{zi���E�&X��_1ؒ��|N�T�Ť��f)�&���D���>��F�!I����-�-��(1B� ��}��
w�I�|A���D0v-U�R��@G� �,c	%���٬�`�' n�X���:���>QU���h�V,2F�-76��vMϓ��|�-�,Z6��������j�J��A��K�^(HZC"[¢C��D�3��?�>Ӑg���=u�醃�v�/�]ĒjE8B�O.��!Zr-ZkHGc�Fv�Κ���[�ش�4�އ���6[��\6̌f$����b^s����r���	�l<�Y���#G��Ғ|����l�і�Θ���åI�?��H�(x��Q��Ѧ+٢��VlfvQFCǖ�셧V~�W��ڏ�pa����'l�������m~��]`U�_�4@A��M"4ă���5�����vݶv�6��3�L�C�G��,�����8jǏ�r�(oR$������QY'v�W���m���� mQ/�Em~��F���	9i��y��c�J2AX�����˦���v���̣u-�]!ps��	��B_�پ�_�a��(����T~��1I0(�3�Q��Vc��XL²�g�@�̯%!�C6f�	������}�������Ȇ�f�r��T`|Q�C����sPq���0�/@a|��*B�l�W.�Q�zZ�6B�z����4�[T�AU$jn�����R,���H	�$Le^W{?��6f	Tr�	������0;H1\��2�5�����x�u�-՗ ������!��A�80��FT �YNg�IzK�j�V�$�rb�oGk�4A���݃���E�i4�dA(�4����w�6=LؐX�?���Jє�[#x�������U��>�NEݯt��0� ,�8|^�P*!��6����\�������v��$�ʬ���@+q���C˲�$���@���ݺu�z��$����/.��P�7���k"���ST�A��U���&%52� )Zc�T���C�<q☽���ҧ�̕KE���p�"ic&u���q-Rz8��P��{x4�f�c7nݱKW�ڃǛBX�$��7���\^A�����l�A&���%��U�l���g��`�Ν��7�cl0L��@"C��_�>�i���0�Kg@�y/�ꕧ�����KU{���?�7~���p����O$���w�}��i��֌��p�Pb���k��h��� �N�R��i�ީ�Í�5:i��eɢ~װ�N����*3'm�h�(@<�TK2ψ�V�Z���l�Z�?�f��j� ��#+5N��]�*���� ��bE��j��Lz�{H%$��\Z�٥�[Y��驲�Q���H�������"R<XߴZ��,�K�,�v9��e��shiHM Z	����)K�_*ft�g2y+�+�<��d*"��
a�)�Fdq��h��,v�v�h�M� �TK��2{����#	P¡�$�Sp&>.L$��!8;MOϑ������^�Ϭ�����3���3l�~I<�ܻV7ë��KX�������.ɜ����?��:�Q���I�#%
��E�E���������U�;2�-�W1WT��^1��t!���@�a��X�t%�W�$��Χ��]���6=����	��+�h��}AU�i�3O��EUHz�NTŽG"!A�B&��ґ ���{�8~� Ċ^k�w.��v�偈v�VEMB���2l$����ԟ|���~���D��y�1�����'OU����I9�`mm�+	�dcyy�
����/�U$�ɘ���L����$:�S���d�T���A�p>#9F#��6,��QD!d#;3�dPR;[���~MD�ǍE���ow��Ʀ�[h���,Tc�
w�i����ԵN��l�y-٤Hz�L�IO�����Nً/=k�ϟ�������v�a��l謯�6��s�h��%�����)�NSn��Ȗ�\=��`u�d/�_��_��Ǿ�Å��~��v2�$��;ߪ���j�۶!�@r�Rt�,h��Np���5�۪2�Mi𒉜L�7k��9���t�k���r�D��\�l(!c`Uz�/�b��P`������Fd�RiiQ���ᒘ8��CF�A��7^Mި�iɡ=h��5�6�pڝ]�*��z�gΜ��}F�w��m���mk7{
�$��跢��uI�O��=�R�nBF���d��8%O��kS����rْ%�D!�x0Ҍ��g�]�g��1�c�#?�"�(��<�[���!)8��S�Y�����+A��0��	�h�%6��$y�s_���u�cJ3~>�I�8��~�Nj[�z��UX�4�7Jǜ����W�g��ajc�A�>�-� �
4����bM��^��=�T���O�G��4�:ẕZz��Q���A�U�F��`�m&f�T�m�5�g�f�Ø5$�XX�B���!"|�,ቋI�@yy�+�f�(I�1����ӢZ�g$o�$��@��`3I( PAU�S�&fl>ڰ.�+X}����׀��L􌜐z��;�{̜����T	#!'�����عs�l~aVH�|ͳ	��!*^~�m<ڔ��L>�k�t��>�p �*��#���?Z&"~��!)	3���;��<���AD��\����N�d�ў��9�XX�2���M_bKNV����9�Ԑ�v��@�	�ם1�_m��e��+��
rhV���+�Cr������W>��]�����&FCk5zBeh�3I!w�.�ڝ;w����g}�9�m���-�:'�L�J�Pٖ
vd�l/�_��_��k?����U�D����w����z�f�gM�P��u�I��/e����ö�ݹn�����Ma�^�fk`�[={�5�T����AOF}�a�ry4���h���>W�v���flL��5��>���u��a���<�d�ꅪ��!�t�q���||T��a�c��*F�4;7m=�I��pͤ��_�W_}U��+׬Yo�?;�"dCQ�ɩ��{}�\s��%����u!���#�67[�~�a�\B�6-2�|��H����3A�bB���H�}��4�T��~,TiHC%*�6$z�a~��F�C��`��/�~2�D�*�RZɉW����%x��@ �PDr��0�6���R���=���ocYz�X4�JFcin@@" m��*��It��d�R�'h3%��W�'pF?�%�Y��Z�G �����,��-~_�?��� �:������IВ�2��fRR5I����A�T�d��<%<��v���hb��Me��LjT!9U�C�'68ȃ�vŲN����t�L[?��Fr����CBBKIˈA���NOZ�8gWD��feM�m�Ǭ�����+��[N��,��gqa�Ξ=���T��k�WEVحk��֭;v��a;y�Ξ���KW���X>L��5|�E"I���I��p#��4.�p�*�r"��4��T�Ru�
e7��Q,i�_��f]p>�\��ȡ|�;�=S	$�����є�&/0��P����[<�5��}��r�#_��HN@�^x�y���`"3h�i&q�Ӱ\��iIԀ�9���`�u)7�/pݸ��V(�ٹe�	�.��ŧ�W���/�pa����'l�����^���S�����bW�,�_F�Qv;�~�}p�=�hf^*��U�X�m��H�Nc(��v;��m�kY6=�~wۚ�-�5����Y�2c�����X�����ϰ�(��݉u{D_���]J36����L[6�諂~b�R����T0�( ��%cN'�k�|�����}+S�j�_���y&�UU�fz9g �L�E���$R�,?�g{�����]�-{u�������^y�k�E*�IQB�D&rL��ι���� �>=	 @�8�9䠧��v�����_�ˬ�7<;5^���%�|�jaorF;���    IDAT22&	!<Q��Q���\��!�ML�,�epB)�xݚ���y'D��TBR�NP��\�ZIb�7���B$I�.O���d��VD
�X�o���&%��rUy���.��7S:hΛ�M�j�Ȫ�e����k�;V��+���n�]4E��
�����[۝v�RSjD��NASuH���N�.Eb Eh�)��H�N��E�y=�Y�>�͗��;Ĥ�aE6]�9W��lVV�}����1±��Sk����'����TmX�C�g�F��ű�a�*#
�ڴ�sZ�ڰ�A��@8h _,�m��x���T't��Q�x��'�>(�iKs��8�U�2i�]�v�؅jU�q�w5Í"	B�w�c������艀�,X���o�
Ԛ;�J�\�t������Ǐ����޾n]��𰼶dg�\o�R�w��*�C��		��(����J�"%�4Oa7M"�[�ƔegKlF��
�!�3&f�u;��xvu�HLb��hNS�G��-�tB�2ZC?�J��F�?%�vS6�U�ē����ح�Q+���q��L���jl�\���t�W��!���:�x)p6�o���id�1�,"�l�Gƅ7��Rp���_H��=�K�A*I
�k�(n_��O����gߟ��ޞ���غ���_�V�:SI&Ku���̛���,��<v��Ί�Vc��$Q(�Ȗ[���O ",�l6�P��F7�)��ʥ4:NAG �D�����2��� 7�z��c}�|�(l̓j͒NQN��r��چx��F<M�9kUx]-	/&M���R��SnX4C�e)�%/�Ύ����#v:�w��$�� B��P�rW¿����Y�z��2����iIry!'~jy3��0Lt�(.!�Vk,F#xe� �+�*�@���C���g���`��������2��<�3mv��YP9��E��F�S,?��߁��*؞�	���-;,e���/vdU����_v6z�������S(���U|�9s���N׼b���9��m����-@�&%�"§��"��Y�ӑ�=�	�����]��v�>mH�]t��'�ms���*�s^gKs��2�3	�P	Aj��fz�b/���?r
�ֳ�������h�Xe
��C��4ֶ}T׉����v�P�:޶D_t�5۾�|~�&FYp��H�x�ܺu+FF͡�g�z�@PB,]y,W�,^�~��5]����%�g4�>ܨ×�r��|\��Hf�3��I�b*���s��$�,�3�xӀf����}��ټV�)�C(��E~t&E{�8���C
�����"t�*!ʮ6�Ų%�խ҆dmi/�0�%b�&��	j��9���J�yޯ��z���\Cu�W�B�
D�h���� q�$�7_4��p&�*�E�j��9sj��+�Kju�:f7�[�1�Δ�nu-��6��/f1%׆0:���n��q���,D�	������fa�˟�����;[�]���r�O#�ۇ*m����u��@��"@6dn
f����r�����S= �pd���)��s#�"3��X,��X����!X͒�H3�%��p��+��	\&Ox��Z�YX=H${���Q��rӊ���s��3� !���&RI?f��.����`�9>9����'��h���w��PMZ���}6#0	%H�=3�r�$���0=e���IevV+��OK�cg�v@w��+�Q�PpN��B$������8�:Ch�J����Q~�I��zl� ���^=r�u$)�6d�a����E��М���"G�$7�È�͛�cb��Z�h��i��"І��'h�b���[{3��� YG��t���Β��wu��t����&��.TO����I�<��h�E�!�0��:ŉ��-�%�ŨKm��:�O:�޳�׽�:s��k ILZc�{�����
9�8F�j̡:L�����aG@5;��۝��Fz�p�"����/��w�~�9$�C�z9��.�-�G�(��Mi�	7R�ՆƥxK�$��a�Q�vlێ���������R�	���<,��n�c)e�I�'��O!#�����󈑾K���W,��xJ���ߏ�Aɢ^�tRIΑ���Z�ov�[�n�hk�e�d�ȅ�5Ǒ�0�[�b9�����^c��F��;��qF^z0�,���Ur A�bG�4���xVb�%�}�Q�I���ʫ��X*@�U��*��L����SȦ�&����rNK(�ݹ �</#����ij���W�E������(ZnQ�$
��_�ٸA*D�*��� K�`7�C�U*��W�.��C	u������:�y�����i�7�c�����u�ls�:�� Z�"L�+9�2<?����d��2ٴt{}�惟��3CK[hX������aT�������
c�[�TRK(�ĜE��09�P/dQ)L�\�B�Tn9�H{z�J��gkrӊ�������T��	���e���v�t':�]��$4B�`���΀��,�^�"�F�:ْ�+�!����f!�	$�.z%�3�d��,#�VN��d/��ɮ���Bv`d O�>]�l,ZЇ�������N�$�E���R�J$p�2���V涄�tț��^�ga;&�yX�！��V��(��t�YZ#����|G#ޔ�-��M��ϛ��Fº�%si��"�:5�Z,x
~���R;��d�ZR�R��f)�T{~*Y���4%��c](R����������TM
��HMT�ª�NʔC�F���pDi�t�2S0���*=(	]mF�*���Ն����7�-1?�6QK���>�/;%��b*3�\���א�'�����N�gY%��X��ߔ�dG����?������![x��W86�9E�5+py�	�d	=|gO�QkO�/��N�d?
�:�
�̙i��f�m�:�4�b�B�9�@����/�-["����m۶ahhH�}3��t��RI�ۦ��p��oQ��%]�X`	����y �]�I��7sbU��f.�h؈ǃ�����튃\�d�
��W ;h[�n���̌�1��,����gE��2!���i�#I�4+ȗ��f�csS��3CCH�Q$�:���2+ɖ��R.	<�k���b�A��H&�5*�=���&v$�}%��D��c^��pf$'�uFG��J��=����ρ�6��G8O�=Q�]��ҏ~잧������M���6N�:�����������Ye%����'7iH���5�l˕2�IqG�5w����TɅrM��i����@��G1?ۤ��dv�����͖��Zj��(WXli��٪}=s��P*6Q�0��d9����"��\�Hz�n�<,_>a�߉�S� nl�|���������$��y�n��9�*��i�]ؖ��dPF�qt���Oz;�8����As}���n�i��F4څhl��\���@����������4��b�T�jJv�@��FW� �"�e�T�"5$���J|�3bf�4��a��Np��车|��������Q֒
�Q��ܸT�!�E�(��*v
��L'�@�[�h�5�!Y9�;�Xۖ�RP�;lkH�qش�&�g��4ܰ�:.E�����NҏD�9d%98ݦaf�C7;�e�؂��49�2�K'a�B 0$�f���)����+sb�wAd�����d0�ʠ���șC+ȜUT�s�����q&�͓EQLQ,5��fUL�^��Ȧ�χ�f*}>���H����O^I�!�йy�ͽ3�e���cH��|�".�:%��%O��p��w&�&3��,�e�t�(���gW\���C�ң#����P�6��,Z��/�d�W^yE��\^����u��c�x�嗹�I�i�L��>�v�JCm �����.�F�O*��x�n�3z:�kM��~��y!�MNҰC��,2?�l�;�]�7�+������=L���V�\��l��dH~"�A�bU�rA-8�#��^�f	� �6'�V~VbCK{J�#V�nW@�R)��L�8q�·`�����ҙI�9�}��}��Q�GR�xxP�2Q9�㚒\�C49C��f�İvQ�K���t��rl]6�/-m�^�l4VT�ե�z��6[A9���ZF��F���Dz\`�����O���AOT�+�BFP���@�<z]je��*YCn*�o0�J]��WG��C��EKS�<IB�5:�x儧H.��ݔx��X��wܶ�3:�у��Tz
����å˓x�ͽ8{fH�Gh�VF��w�0��ʊ±���2@�lź*����S��Bw�{����@�N���\N��@j8���9]X�|���3���D�b>/�?�+u�$:H��H1a�FHP�M9/V�7��/z>a��Wi����:Sz�Y57on��ѥh��Ɛ��k��Ѻ�N�F$���E	���UX��I:�>�:^�2�",%sf53lä��r��.�=�{��T��]~$,���wI�Dc���g��U,�:�(�͙�:��W�@���4;�em���}:ߗ���|�6[u�cӓ�y��dg#EՑEq�gX �d!�K�EKĒH/�I�3m'%9D�Jeg� ґ��6�fк�{JC�Iƾ"��*8�����yHy��%�y��kH��K�[¿B��҃�=OV�gJ�$�I�  ����Ξ��j	y�P�܅K�r�ĩ��,q��F/#A9��ZRsfv���m:"A%�y
�gϞ��˗c���^�u9ܴ��NŰl�b�v�H�ꫯ�����Y�>�ɊX��p���>£܇��G�t��w��Ƭ�ZfU���������$qM�ݸHP'�Z���0�����V����M1E�n![����4N�A>OT)$kN��l���B��a?�P�LI�UD:���O�X�qT�m�������P�Ѵ��U����#"����į<HRI#Q B.J3,(��3�^D"1D~��a����̳���&H��}0�O����b�8�Z.m����F���c�SΜ���5.NbׁS���EA�_p��"`��DT���7(�p<	�f�H��Ġ����@�X�ɋ���dmN�ӢE#|LS�F��X�v֯Y(��� �(�����Yȫ�l���g�8�d�Q@��KH�)n1��sd"�0�E��|$��N3J����Lx�p+��wnw�;
��*2\�;�8�²��t�L4�YL�;9N 	\��x�@ p��\�z�g=^�y_��֠�V3j6�^�4=?ږe�L�mkn��b�����tM7mâ���lY4wӶ\F˶m]�M7��鵚���ntӶm�jZF�l�����8��^�9�N�?g���i��kv���А��^[b��t��u]7Z-��4�0KȌV���n��0,�����n��[��ٶ�[6E6�vٶ��4M�5��̏5ڋ:8����V�0��U��J��l����KT�e�����-n�-!�H���lw�r0p�y_�"G��ֱ�J^3�����S9$(���!z�`za]+�Xu�����t����>&匿GNSl<T	�UYh�i�/�E,����p`�gb��$Ni�[N@y��k8Y�'����M�!=6"rv��P-âe+p��Il۱�B�bU6�wwۨ�Y�^�!�����-���c+C�����ѣb��/ɹ�m)3�fH�ߑ���2%W|�WC<J�J�|^�?_u�K����#an_��֮@w�jM��j�$c"n�"g�^9�(3����I]�|Ot�.F�y	��AY�'��$DC˰P�4p�Ro�����;�uE8j�B���b�JRl{Z�nW�.T(Q���4�#L�YH�mc!o���z�9�%��1ǖ�A'ዟ���M��x�zT>�d��k�����d#�űb^�7?�ܽO��zs3���F��78<<���ÿ8:2���/k<Ο�=3``(��{���s���T���l�B�`�	�@rd���!�*�]b,B8����ca�6�L�Ã�ON��!�FCC��4����V�fq:~��YK[�_�k�7�|��o~c3�='����M�X��]a���}�(�7M!Zp�BV&	<������	f�z��a�#]c2H ��
;[�le�yi
�հr�,�׋\vS�a��$���J�\H������}�ҥo^���A},�Sx�:q�t�4=�F��L�XT�b�h���6C�,�����V�e����h�j���].��l6��mۆ�e隦Y��j�<1���-��ې����<��i���T_-]7�e�-b��[���u�z�˟���-��]-Z-90���VK�m��l5�iz5`Z�Q����tA���2شݦ����i�v7ZZ+��:Ep^�2��H���;w-O�e��u����-�i���Ms5MS�2pϴ��W�4M��W���,�ú4��|�a���a�ݞ-�SRLf�K��tL-J,�*�v��\�/]B��.�<!���ڀ+o��S��7�"=U�$	�,���DMؼU��	x2�ptĢuB�S)&�4��寰��{P�j�T�!��:�ȇ�����.Z�|�7y&$|2�Qx���kd���޻o���n$c~X���%,R�b�BSy:��E.�P
B����˳��8�����D8,S��b��#�f��&JU�c�>;���2,�Jkh4��\�8g�H�*�y��UZ]a��G3�
���b�Vi �д.m>EA�>�-95��{�s�z.)�#	G�c�@�F$g�Ļ�b���X9��O=��_���{ݜ����Ǐ;�'�l��Ŷ+5��a���"Rl
N�e^����2�qH2���̈4x�|"3&�5Ǚ��*�W�5Q)W��1�)���e�~ЏDW'�.��eKf���I�r�){;v(�7hx���ؿ�m1���̔t��&3���+�fn,���[�XB͒[�	��S��$�j%��iT*�4L^�*���S�*
ڪW�ɸ`n?ғ#���������9��WΚ�}�������Xbl�O�8�D"F�P��.]*$���d��ш�u=�-�˱J��u�\#�B.W���f�i����zm�[2�$�e������@��4e#d�J��_(���lv���D<�̈́�F%X��\<pr��x�2���v����?���g/��E�]k���T��ћY�@�X�퐥�K*6�IQ�T��'�@YJ{F�B���&/�G�=�g��[8��_��H�d�*�Ͳ ��������ᎵX8o� t(Q	a��&39d�u!�ۣg<=����� k���4e4��:]���Zy�B� ����8p��5zV���@�\���H�Z��"�4Ju���A#*W��<�$�q�m�Zd^+�dI��Ywۦ����5�Ȇ,z�/%H�0�"	J'՘�!(|l8�D(@���ܾ�Z0s�?q�C�;��پ{��۳�䩳��X��:�ܶ�H+�/a4ü9� �z;���F�!y�J_���-%����ʣ��EY�0y3p����Q<x�)�wx�Luc�m˱r�lx=&<o6M "#bP�E�H�������#a�u��#�5�BR4���z)�.7�����<'���Ɣ��$!nz��߹Jل�r�D6_B:���4/L��̝�/^��d�;=�߼��;�|�.���2�W�ǏM'b�r+U(���Թs��%:��G�����o���shڴ<����ZM�g�^�#A��!	S:2-���Yrw�t򢍩�)(9C/hZ��	�#sfՎtJ�W��Q���$$A��8�3a�t��i<����a��>���xt�]������z.Wl��Z����5�7m�V�Qt�|c����2&�۴�-_�QNTK�5�rey�R]W��"�_�������Tk�04Vƾ�g�I7�ĥ����2�#W�Ex�������w��W�Ԏ�g���������,_�+2�q�ԘB�g7���Yv�O@T�/r4cP�7�hLbE�0��Ê�3�=��;ￚk�f=�*�\�C���86:��ͺkV�Xî�G�G�z�RI�mڰ��2v�#ur�#��Խ�g'�CJ��ܐ��:Ul�$5��;Q�R�    IDAT2<����Bn��}!�`��a��~��<�%ֆ�mG��,i��o��Ǐ��@o_
wޱ
�v!���6����3� ��H7(
o���ޕ�t�7�ئ��"�)�����i5�`�"��9�������ksf���%K�\�Y���^��{������Ǟ���;�&�{�~;z-�>�a4l�m̴�ۊ�L�2�h��s��d�fSF�Tv,-�Z�4�o���bbC�&ۤ;ZP
<M��dF�� ���lF�ْ1	x���M\�p�߸\z���
^����MS�,�%;�K{{{+ײ����|6���l�^[�dWi������<��?��ᢐ��rG-8��pA�W�˜O01K�h��ғ�����E�z{%�^�L�"BG�.��?,P7�]:�1[X%#)�1���Nx�P�x"��j���%��H0`n_/�ϛ����w�������[��rAN?������]'.\B<���5�����B����5�3E"���V�"̓]����Kje�K�\%6����h�wB!׀�@s�n�mX��K�m�G�!�a�����pN:]�k�o��S���zRx����M����� B�=oBFeї�L_����@�6$ϘuŴ��g�Jż̛��8/t�0(U��x�Y�����-]���+}�/���^���/^�m����p8����K�|>+�Ha���h\����B�=A�*5���^欱��|1�JEg�C䋉c����B~�1�t�P$" h@��u���铓���!T<^03�x($�Q�>x�߿x��w��V���u���ȹ�~qhl�7�;h��0&ŶPTNy�Si隈���E�[ɵ6�� �L8�{�)�"C��ϙ�P��X��ŒΖ
���W��Q�\�"6V���T���|I��,�m-�?��?7~ތ�d��D�`Fω�ߴ�.�u?�-YlGFF��?ܽ��O�D�3��V/��Ӟz�	P�J1��Ѕ��D�)Z��!8'���dC?b1���nU!Ǚt^�m6C�S7|�8�ް��t��n!ȹ��w7�1A���^{c+N��$�3e<p'f�H �7��2��Ŗ]9�u�8���� e��]6Vu�n1��g����Rqe�Y�t��RE�G�,�?������{�W��L��pv��ާ'''���<4��xiPؾ���>NHŀ�N]�EZ<d+njr�fI��Po5��!DFp�%J��B![P�⨥�U�D,)��D��''M"S������lSS˂D��G"�8��}�G{l�߿�K�mǶ�9?|�O9�=7���}'-,�y�H�Б
����F��]�|��xA��V�UjV�X��IԞڇ�5N��t��'�;wbG�.�V�LGw�>��lN�K�iH|^>.��
i���TW�@�Zӂ۶��DF�}����sݮ��o�b+����~o�ί��0��TkV/���F��lYd9�$|,
�+k�\[	�➊!c�婌Ŗ]����i"Ue" �j۪ػ�02�*�U��7>��:�ؒH�$J�^^hlÃɉ����95 ���	�w�z,Y0.�D����������<!�IjJ�U�VY	�Ŭ2�P��dr�BM^Y�n�ip�x��O޾x񼷮�B�~��
�
+p��q��Щ	���ti �c�"�sS�b�P�*i�L��}E���t���D�]�K@��ӭ+�&>6�ɉyG��渹\Nrlɶ?b�d�ЙH"��Vm ��R]��N��~��%�::�)��������?��=�ܹ��^�W�x�K�F~i|���m���V4���.4U!rr6ʝ��NK�9�K���Hz|̹%�I��Q���&9a+�pD�\�E���S}�l���p���S,
y�$>��%%fDb��t�~2�� i!�����4M��} �n�b;|)w�w�������Б����K��0|�(Cv�����b
�IE���'�bQ*�[[��DGF0&.��F]�[�z־k�Le�(V���Bx�Cbޜ�*�n]�>��.~@&��RlϞ�_ ��$�k����m#N)�P{�[K)��J���3�T$��hP+�v�L�r��R�"��zC��mC�O$	�l�,=��Ǟ����:�~	�+p�+�c۫�ʚ��d�Y���˴�B�.�V9P�\;�H��N�Q�n^����O< �1T���rA�$v���$_�ja�v��8��b���y;&�Ɍ&ш����D��aFw�4�>���wܱ�{W������>����#�/gCo���ѷ�	�_�X(�r�G����9%��|�.ѦLBb��	axF��	mD3cYHZ3z��C�'������	�g�g�ݎO�4�י{��li���ϫ�� �(,z�V��n�3gN�=.���[��NL���~w��GOF��	�^�7O[E�D
�__��A��%�Vή�f�KN��T�sAv����bK�;���
�nۋ�t]�u"�q<�if�&��F�>�,-����c|��o��g��I��v��+�J������W^���xjS|
.Xݨ�R	o.�DC �
C�Yh���EԪMq�ἪX�fPa�������;�W��N��h��[S����rS�Tjbg*���U&;O:'�����@ɼ��gL���)�S��jn��|�T)p�Q�*�d)�p��( ���/�	��a�W�<Լ�&����W������-���~��k��Xޯ}���?|�ѭ��ay�ӎ��@y���̸���}�Hu$EJE��ɩ�h�ň�A��OR��>k�߲��AmW�r�ĸ��P�����>�U��B���}�ӕ�)\�D";I���=ntœ0kuX�f��O}"z3��j�-[lm�����o�}�����f�j��1�N�ζw�C�b�)�u�;��2����ӛ�tf㕹^�Z���B�P��-�11ZA������6`��>)�~�`	Q�L�m	����q��(6oރ�Y�UB�Ѓ��M�C{8,�a�.Wke�GXly���Z):�=���U9M��R���XB�r�l�J]�;؍3��T*c��y�^|�S+���~��
܊+04tq��M�G��,p�XS��Z�x��dQ$��e��B4��mj2-�d"����ф8J�����eť�$E �'8�-�1�J��n��e�� ���u�dq��Y���D�P44$cq�k��g�]�lٲ7�s�ގ����}�s�����5���!w�l尟/L��[�{=�n��#�	�m��R�C\���b>�&&��,�,����bPb�.�j.���Ï�����Kt�{���t�b��PH�m�T,�ΰ�f��矋ߌu���q+[㥗�yl��cK��.�X�D��̈6�tM''����N:C'�5UX�99�$*�pI���!0�}J4��l۷�Cz�a\�*�~&��L���6����	���Il޼c�94�e��^|�������uǧ8��`+�I�pir�-���R������W���g�+��ސ6!�b��/���6UA�P�sv<��{����W�V]�m[�v���3�8�-��V�d���x3O�E�HŠ��#Huv�O��ˌ��nm�>￀/(�~�ٜ��0��	z��ł�,���Q�'q��D�'���#���}�1Cq2�&�^�C���zj��U��n�������}�y�A�.��\*J�fSf�S�,�VU<�a�n#p���7��F�Z�@��}n�	��
C f��9����e����&�'�W�U.�`�bW�r��:��~��-�X�h>f�'bQ�-�'��Ii�ef�}����X����l��|�o���d+�/mt	���G.w�;E�'�#���*��
Ơ`��uxAH1��5Y�:���9�|'3y��f3�MFć6ރ%�g��|�k��R��2l�.g�u�~Nȉ��;��>tRQ)����Xl	�脹��F"������@<^m�'_0z�s^j��Ų\�<���R^@�U1�0g���=���U�j/���M�����������>�{�v����J�ru&L�!=�+�H�э�-��#�(��)�\��a�1��[M3V��5hK��e��SR�Y$:~sXM��m3��{,��K��B�:�	̙=!�O��\}ᅏ.\����#�>�ږ�_s�~)�4��Ix��AT�Si�����\	�U��ք�Ƀ;VA	u�x� Ie�4�iӽ�W�E�&�,�c��8p1	c�"��h�%�M��S�����C�ڰ?�h8$��Ŗ�p���<����rͼߏ�e�-���կ�<���d��^�.�&!Ɯ�V%m-}4U"o.�����IGب���iY"�23�5Tf�,UD���鏅Rń�J�]�`B:�
�M�*�fˍ��v�:���c ��/�G6m@"FRTMY��-���ar�*�bo��=~��kKڳ^Ȓ��P3![�E넾���;o��7�~��M��E5���+�ϽǏm��CG���y�	4jn�5��[�����ʈk�e	����Y�G�{b���Œ[z{�c��\{||<Y�����ٍ���O�'Vf�?�m�R�&	O*X�hY�Q�N�m�(�"�P�4�~��1�'33��#){�G�����?��f�c�|���;��y�A�.D�Qt�]�yY���b�L��S��#?Sθ�����ܣ�ш[�{ ^�Se#�|l���������`��ǵZ�f�f�Z���\H����0��l W(H��s�e�
��sy��2�lԧ��������ݿ�V.��?}���>qz~0���+���VI/�8xg�R�^����v{vx��=0�3���5]��ͦ�V5o+���V+��:��b[��ԔZ�$�6=���=��X(�0"�����j��"�Ug�Bn3y�ncd��=���q)�3fD��Cw�#��LK8�x�H��$|n��f�D���[���>�nV A*��|>���1!lp�D*>!-����+�?��?��O|��tN���x?V�����ȑ���la���n�*M)�,���[�[��<���]�p�˳f������{]/��Ҫ�O}��s���3����$�;n��4/J}�#-8��,$�q��:��	yמy���-�a��F���c��[w���{�T� �#恟�(&3�(��҂O�H��*���B^��ю�"�0�Ʉ�sĵ�R�U$�1!)�\����#�Ͻ#��d_�*�lv�չ�܋cc���zJ�
��H�� X)�!�G_��׏�x\����tg{#.
>�����Ǐ?5'
b��5W�-���b��*�Ű�������ڙL&/j�F1���P($s�̦b���byٽD0x�T%�$�Hc��c(t�l=q?��,�����B64��h=f��Z�c��#��b��܅���:%;u�}a$��t�̹P�!#!%|�GSL�Dg:�����SF�X Y����LȌ�J�q͟�蛏?��*v�F]��3��^�#o���o�<�����k6ju�hl���D��
1
�8�Q��e+��ڳ��׺�_�O���7d�̅I!��k�ot��.�,4,R���$��e��02��T"I�n�駟��x��k}M���G����wv����t�+��'�k�9E6�e��[��C[�G��)�!��#�,�f���IS�4DCat�:s���D8��K�,�����[948�����G�G�Qm��d�&&#Z� �@�hT2�k�r����|/��~��-���r����r��������[+�˔�p����*���.]��X����.����yS�����'h���f�d34<�=���R�o�Wă��Y�y���w��b���N�U����v�9���,���� 6>|z�hTT�I"Ì�>$�1a��*6dCh��B���uB!�a*,K�P��� ��<����L��:�MMA}����y_����<}��0����UW`��W���c����R�2M�I��Z�ôta��"�0�,^��>��/�����?��_8r�į�3Yaʊ ����GQPg�r	��b�n��cQ�.�X�;Յ�=5�~��7���`��n�{��,�SY�HF�͢��Jy!<IC�)ubS!�t��XQ���Vlg#AA��u$�3g��Y�f�ܺիw\�Z�:u�����;y���$ш��*gۺK\�Ȑ���b��$�J�8���ϥ��w܌�ݲ�vd�бm����]�a��c��0x!�x�nx�.��R�E-���u1��/��J�˕��	��R���}�[Rl	EiA����)9��J��XB��6�ǪI��wb���M)��>z/��X��5�tw���CI$E�"���9���Dx����	E𾠐�ƇQ.�b;62$?�����k`�%���?�µ����W�V[�];��{�O�ٯ�l�"sr�z���Ծ+�+����ӫ׬�x��g��믿|s�ַΜ=��h!ζ[���ǚ�(�P������b;96�d<��3gѢ���s�͜?���X���w~~�[�~u�����L!�P�D~���[#�H �U�K��uk|��C��16��$�.Y�����+V���C��}G�����̖���-SE
�F�%�AOyf�K�<�l׵�����l�e���{Ν�x�C�ښU+��Jw[�U�����|O$������}fl|��n�����ĩ�g�{�A�J.�k�����5�?�����z�(��6�����ؾ�-��r‒Lz����ˉ��B�`��4����+���ڶ=#�ڔѴ����"���@��EzbD�~�����se,]��ˏ<�����zL���
�*+�־W~sp��o��J�*�9�2�5%��'.F�m�/]�?��_^�{����Ë_�[��X��G!QL
k��,dJ}¡�J�1t�Ǚł(;[�6:bqv���|��+���]���޹��:y���ܲ�&�g�BGL�iU��0�C�^V*	]80��+W���
� ��Hѣ�ݦ���*˗.{r���߽����s��[wl�:82c�e�^��|^7�� R�!H1O��ˎ?������z?~�.���];�]�t���p���j������\2��[�����������f�����ⱱQ�8y;w�uef����m�VbFoѐGR̋e�$ۑa΄��F&A*;�;�Dҋ�=�H}���)���l%RkKTܔ@6��9��Db����.E�(�xǐ������Sl�,(�-aْ��C�����?6���
���<����֪
��I��U=ސt��` ����w�u��'���m޼9��+�\�py N���2RS*lZ�z�(=J�bQEp$��,�+�2*���:�	��ܸ���ׯ߰�z_������[�ǁ��_�޶��H[���Gg�@Ӭ�4g,=�R�"����S�ļl]��� �A�_t�$y6ku�BA,_��?=��S�|�^ůny��:���Fu��R��"���HI�%jP�eǞ���=W�o�cn�b;ܿs��K�._�y�n��0::c�9�LM�����p��<EK�Rw:��
g�FCC�x��)l߶Ŝ�L��Č����I������Rf�Y+o8ہ˓ضm��\Z�=a<��#3ҡ����4 e�N�EWA��|���Vy��تt��22�q��b|bDd@f]͜$�l٪�޴��Y���^��8��_:�%�;U�9n!�WIYl��n�Vԓ�<��?�3�o���������{G<���X�m�_�򋅞m[n�ζT,�Z*
Y�Ŗ���}���>��7o���Aϳ{�/8u�S�����t3f�D*ΈQ����ؖ�U؆W�1���+���V�h)���`X6R�ܳ���-��>��}c�w���Sj�Ieh���.)�,j����'^|a��^���F��ܱ���A�h�|�	t��"�iu�:���C���b*_,��=�U���A�9s[��E.��D�G�{��A���*s�v��ْ�X�/�a�=(���4̛ߍg>�aă~a�@@qx<����Fl'a���~T���`*�_Td��    IDAT�Z�eӸ|�&&G%2�R�\)�K�.��Gy�'�gM�vzn�8���ap��o��@�l�D��7IbT���Y�^����#7�=���~�ؑ�o/�HK�Ѹ21b�ʑNЯR��=��j����7Hܪ�Й�Rl���G�ܰ���~��=x�t�����K�%���0>5�R�&��a)��8�2ٶd�S#�?L1���M��}��>����s�߈��?_��7Μ;�
I�l�Ồ���d?-��^�ԧ���X𡡡�[��:584��Q|�'��J�hbr���D��<��k���+r��[�`�S��1���������]ȤM�eJpE�x��MX�pZ�:<�]�Z��VC�C��ضu/J�2��b�<����%t����)WAnɒmۓ��5l��6�0Zz��j�h:�6�h/Y\�xc�^��J��E,_��O~�#?{#��9�W����}�K�C�~�r�b��L��R�)v�#,:HYX�p����'��7����~����GV�x�𣳫K�.�X٩r�IT�r<�ݖ�Ff���~��R.��c�/[����z}?�yv����C'N=�e��N4���'0rˮK��d.-ŖV�F�%���͚�K���#��^?b� �O㑍-Y�p�U+B~��|}���صk���b�c5-q�JDb�Ffg[*��_���3�q�\�4�d��]'�GƐ�㑍��MÐ����k�G���k�����O���?���ȥrã������X��*��6<p7͟�Հ� <nZ�5�d�E��q��8�nٍJ�
L�q�2��O�+{�L&��u�2��_r�]���~��w���%�
N6͚��i.�,kU��xĶ�t1�ϋB.���"������	i
%,]��?>���~�z�d�g�W�VX��������S��.�X�cj�!�V��$͜���/���'_��&���/|�螽{W���DБ��c��`Ifn��̿��%����["��Jv�>��G�ϙ󃵨7��عk�+GϜy|��C��@�x#7�2<��s�(�	���-C��İ�ٔP~�=1��f>�3���3�X�z�S=���o�kݶ�Ͽ����q8�b�2I��Eg�b˙m�X�x�����7b��//ں{�)��T�n؀޾��.i,^,�?�L���{ȗ���B������d��W���^�귤�fKM�����u+�d^?<�-�'���Ƽ�T���Z8w~۶�A�\�f�q�}k�O=�x0(�Q,�s��������\.�AM�~h�m��f����wX��tCO�}��91�P�*����˗���l������1��8��7�hp�̿"�˗Fn4ɰaڂ6��vvv������{n�{��/~��[�+�� q3�����)ώ�]!�l��g8[�d�X��=��S,�����]:p�^��lwn~���s�v�;��-e���V�ox1���'���2Ŀ���B�ES�AEö�A�+t̝3k�ҥK_\�b���}/����+;v��B(_g�,�a����Tȧ��Ӧ׻��yv�۶o;108���.�}���߃@�����������H$:_}/�/��<;11�z�Y�0��B4���z���-$g������l�
"�$˒��l-4��.���Ѭ1�����_|a_/N���_�ř.]ߛHt����f۶����o��͟��ŋ��/&���2�`ي՟����v-�=����W�؁o�֥����ޝ~��<��^ѫ���I�\��&������+�_��f����^}���O�=�dsB�d!et�,�c�U[�)1tD�8:����T+��3����$rSY�c��+V\7S�j>�-[^�y�셻w��6ҹ�z��JxQ.d�+����u��͢�%�V���.�^I)�8��D�D�` ��N���~�0�-�z��|�#٫yM��1���o�v���GC���0���2D��G��r���/<��4�)��[��|��Ъ�{���+��Ć;�#���%U�Y�crb�`4��L,�x-�����&_��
��Ѳ�"�Q��k+�Pm�g��^�s�t����g�m���m�д���z��(��}����`%>��S����`�9`��D:}��4�s��Z^�m��f��#c##:6:*d-���f�b[(c��՟۰��-�=����W�������ȹ?-�K�T8��HG�-���0<���c�mk~�ɏ<���}�/��گ�����ӄ�����hm�A��Բn圸Ѩ��a8T�6ͯJ�21w�L��P���Gn_�b�[��ڮ��7o~e��K���<p�&f̜��T ����'�|�(b���2�e�T#�^v�]�1��g����X"]4�/�]��+W�z��c���ߺ}����pۇ ��t{şyFW�8Y���I�R����n�����vt�����^BwO
�߁X4�2!)�E�Vo�q$��`�s�joʞ��'럚LO���TN��[���L���19��7��&�Q��^ܶv9��I���ѽb�&����YB�a���a�8~�"M/rX�~���#��������������?4>>���+�_���r5������Y�L�FGG?6����DF�e�S�4��ª�k��������}���M�����o������a64�ccY�-.�Mz�6ivQB"�D$�s��{�X�n�5;͵��رc]_�[{F�&fCQ��Up+u�Ȋ��܋&�S��R���|n��ԥ�Ι94��������M��vۛ7�sص��WN\x|��#8����>��
�Y���R^�l�ZC.�uۖ���L."S9��D�\B*GOW
�xt���'f_�{�������T��
��s���Зꖀ�l&W~����������n��޲�v``xÎ��v�F��}�:��>xt�P^:�4����\^��t�];4�S�o_�m�bfA6_�D�X��JŊ���.�lݬ��#��t���=�r̫�"�Ս�n_�y�pi�,�իe5�V�z�NO��/����Z�a�<��F̙5�-�m����v��������~�۝���������a�57���j�G''&~��J��l[��b�A��pc���?�d��?����sM��q.����c��^�!��`tt�� b�Ζ	=D}�y�]0��?�싿�^ދm���~�o�t���?����&Q��Q,W@ so����˽����D�Oeq�ZRl�Y)��Ѓ�h�ڵ����u�?�}��_;qi�ѭ��ƅ�*z�fa^oV� �2�/da�&l�%Ŗ�#紤mҙ��	�egGB���|�b	�pH���S���oÂ��������ٻ�ѱ��{S�KF4�4����{�l#�͖����b{���{��#��ܻo���(f�����"����,��^��>蚎�����8ʕZ���n��=���n�k��Ъ���Z�V+���j�K�ULiѨ��U]WNLf�xc����6!\��!љº;Wa�����k�|[c��fJx��9?v�B�R�D��#������Jv�r�V�<x�g��B����02�X��Tw��=��m��P(Ge�RI�zca��z�R��t�R��lV��FS�))ٶ-ej�b�j��Y�`�5̓o�g5��+p�W�������إ�3�:8?�(H� �Q���:Lآo��/ؘ�x�o<���x���[����;�����QW���ᒮ�.R�|�RY�2w�ߺ�5��y�^�#Q�b��l���I�y���nZg�y�+o�ش��I���9���JV�n61���is_sC��������
H�����U�T'��l�0gf?����˳O��u�OMN��ڹ�+�N�������&>�O��̲��wfO��e1����=]�0���y<����{��Nb��YX�v5.�D0�F��S J�"����H�`�@�9I��� �6ZR'P���!�XL
i�,�bILfJx�;;1>I���xw޵Kv���MC�Yl��o䁋�:9�f�)<Y��{��}���"�L^�e�b�#C1^�Ԫ1E���ex
>`o����`YfW�l�i��yj�TA��b����hHG��C��������r՚O̟��o��O?��
|�W������ѱ�?g�M�rLLaZ���5#���j�(�bƴ��f*�����~aݲ{/��7x����/���塡w��O�VC2�)�Q�d'�j	 ��0�q�����4~��V\��&ZM��w2�e���c�޻lٲ�N��a������q����N``����1�;�e\��da��BKږ���I�;̶-e0c��m�|NH�^�!��K�-��M��h$�\����`�ș����{?GĀc�2a6[�ǎ�c�����B6Wߴ��x<���u���g.lڱ}���t�kV.��c������;]]Nc�ܛN�+OD�0���A��uKE�*݆��A�ސPv)ht�F����{[�cp8�ZSG��[���E�pUxu�c��<�R2TE�f����9'��`��8�A����ғ�f'��L&�UƦL��N�,�<ER7[��d���$՛Rh	���9#B�	��� �{�W��x�M ���1�׹������?���r%L�P7q���(]��z	>�[
 ��Z�^�G�͙�ծ�ԞD��HzN:�ht��^�F�f����V���J�O��k��%dܴl�O�x��a|lB�E2����p&+���+�~�G�\&��3���V[�M�i�m;^�Ι�#w8�KcuF�CotST���-��`�4.Y�f�y��^]io9C��,�܇Kż\�K�,�����5so2�,|��{hh(yq��#�G�>s���G�ryA�*��D��6	����i��Q��b._���R��}���{��[�؞>};���)T��Յ��������1_��W[�|�Z6�]z'�Eׂ�d��7 ��,aֱx�غ� m�&BO�'�L�������PŊ�xG7�w=�.��U��:�K�-'�r��r���<:�f݄�U��EI<��Q*�01>�Z�,�Z6�v���7�?/^��'7'�*��mπ�Պ�NXh���xUl�U$�GZ�ė,_������/�=]e�?4�7y�~忎O�U�r�t	�̆!Ŗ{��fp~[����w� ��z�`0�	�Be������4�!˴�9o�l��L�%Ș����Wk5��8�䁞�,�����:��⣮��D�Xtg��J�⾳�፫-Zt�f,ߖm�~�����݇N��}��pf�z>�Q�%4A�%UM�d���&E���&�Vlk1��P2=��^�l�c�?��HmŢ[�8G4�B�J5Ѩ7掏�dpxtU�X��'�"��lZ
��ڻ�����>����Ǟ�۱�؉�qqB�n^���E�*���P����GE�V�JP�V�TQ�� ^mR0	�4�	�!΃�1��g������[k�;7�a<�վ�5��{�=����[�o}=��d%0mm^�w�`�Tk���~ۭ�l�`����g���w�|v���Ԍ}{w�2]�U�*qI���\,G�"�G����^N8�B��ST�(
�*G���5�>��r\�FG��>C'N5h�m�2<Aw�u]w�n�F)i�K�=xz�	i~�M���=y��0�P%4���C7_MSm!�%4=}�ʢGC�5��0<L�Cüp�	C��C�FÀx�k� l��i
x�#���g9�숮��߸����������8���?wf������L�sK	��%5�9%	J<!�}�.Y���T��@+	Ҹ�gh��T��P�q�96��Ҍ8�K�%W���:�q{�@E����� d��hƘ��x���pI|m�F1b����\}�e��*}�y��gOM~���Og2ڵ�bڷ{3�E�*��
�Q�(lq���o8����t3|���2��qn���arbG�8��Z���-k{nn��ACWhdt����n��8/HW#�қ�� L1�6��ew�~��k�M{��=�����/,���6�:9F�22��
�Dy����\��R_In(' ү"9(�|��j(Fz	3aѢVi����L���4x{�FW]{�x�>ں��`���#d�B�tv�E?~��>5G�V�	�Rھ�F�#U�ƒv�z�� ���رh�GX�fxh-���� Aɂ����^�.�B*L�Q1~���4�jvi�]y��y�5X��Ǐ��ߜ]���v����V��� ���N��@�!ơϣ�J8�M��M�ƱË���FT����7�:�Z���#���2wZҪ�H�^��~��b�À�_d����������������+�����>tbvᮇ�������/��6k/�h�FrV$����n��@�B�z�.�n�שˌ�Y9D�l�0d�#B� �{8b#�uY��pZ`�0���l^�-:�7��-�u�� r֦��{�׽��-�v���� ��sss��?����={S��4�$Mn�P��!�3"��M�V�%><�f���(�5��<=c|�S+ ����b<��cʩF����3m�9ۡnY��ݻ���Ў�q
�V�"���BөSg��ggi~v�L���H@�.����L�A��g�SN?W��kr��1#����`!"(L@e���0"&~���@aS7�i~n�tX���yׇo� ��߂���Z�'���gN��)X�YJ�3��=��nU� �x�G,�������c ���$〣�-;��ý��'�=^�N� ���o�uУ�~/�� �5IHI./5{o|���߿����x���|��������Ћ�{���t�ދ�h#�U��
�QG��p0d6�L0�R\��̔s����@�@��
�D0~�EʒJSp�"cCAje�e����7�rx ��3<�jk1ö�s����#���[n�urjjjս�km�lO���3ǿ~���p������W)�`�����-��͂�>���4�r����G�e�P�`k��$ZD�>�B��P�V�hv�MgZ��GFij�m�:FcuQ ��)uL!jR�U�7�^^��!E;��h����`�1��5�`���
� }e\�Ml�e+Ԇ��#��p �� �M�Ann��.6�_��ۮ�����B����H8��/}i�1�� �Ǽ��@�
i�
����c��qM8䬊$<	 	������J�oE�,4���N=����O;0E�&{Q��}���EtI
���)�haa�8|�}7\s��'^�>��C��_<�Б���LF�쾄�?����9�hG,Ʉ9:5
�R�[ɣ�V"N�;�e[، �,?�{Kx>�����!�XC3�2��A�\CB��`3ͭG�,$vVP�P%�2�V*Upmʻ�w�O#��ʙ���6��|n~�`�"}���)�DV� /I�p��F�n� ZD����h�B�ܰ�L;|�PI��s7��5J(��E��ҹnNii�h�@
pbvf���S��qޔ�f��QIM�h(.i��x0����|F� .X�������.�� v!��N6?K��o����ל.o��43�@��_����z�G��#�/���x�_|��5n�r��
���%X�=qƵ̀1��P���N�1Hc��(�G�5ҊA�(���BH��<�V��s����H&
�g��E���UW���Iiz����[�~���_�v��|��GO�����#Gi���}�죛��K:kPL��̨����� z嚭M�fh_���
�S+�4��\c�GH�r�`�nq9������`���9���A)��Z��n~~Ѽ��;'w�ܹ�Q��Ξ>��fs�3�n�Wt��(v
�~�2R`�� w��	+�AԒ���`-ᕕ�9h9jD
����o�!AmI���Y���U���甤�YS,h�5܃�c�m��*L� �i�UECUM�=kHw0+)W;����Aċ\jA s�,k,�����
'�$ ��2������[''��"�ʍ�P�}x�R,,����=A�لhLһH��8�E٣ ���Ƕ\9"�Hi  �IDATsNkYH� �b2MP��A*�Eul]����^N2g�lM��QȈU(�j���L/<�"���x�o�ֻ_��~>�;r���O͟�����ť����K��EUզ���G���  ��e]{�!d�X��'ס�����sbA�<�B&}:��, �l����+n���ëę��8S*�P�(�B���b~���l�i�U�c�_|n���,y��bW%%9�# N���V�9p8��&l[���-�lצ2�Ԡ�*$r�&DA��S�T�=��.4HK5��Â�4#mb��T�� _�{#��툾r=�H��ʴKqH���.@T�{F��CP�B�ͦRd�J�Vf��P.=�.7�zkȨAmEj�5��-[?�o���ʏ���[`C[��������/Z�GZ��B��2%a���f0N��>�=�jHR|�Ij���`�)g�?�3�����e���������.�� ���!�(�R�47�@�>�"Ml���ݰ�����}`qzqi��G����wҍWJNa����B8f
�� �B�"$���S�W��KP���M�BC}�EFJz:b'2f%�}"I�K�"5�@�l�@W9�87�����C������)]o��?�W���}z�ūgN����,jpE�P|�&V,�0� �C�ʵ|���L�����67F�F `� �KM�P��
 V���P'�Rty��e�B��xhJ1�V��K�XH�jD!@�g%�ڎ�L�Lכ���Ny��-�x�跕:O@IW���-��x�D$#���o�kx�?�ܵ힭×̮����-��,p��}��<���T	����[� �1RPJ�d�CZ�Q#FH���FFwwK�`2`�H�P�Kp�"(��������=�/p�y�s�s�|���5��UP�PKm�0)��. �l�f�
��n,�f 0��afǳ��Vo,TA����[�����9�|���V����9��9��?U���xL`��7{�@��+��l�*Eq��z�zu��Vr5��Hi��O��?�>W��(u��=�Lw�b���O'���^��K�|��HK�Y,����Nl�a2̟�_�t%t�~��U���p�ʦ)2��� :��)��B���_G�=�`�J�2�q$.��O�o��E�O�\�x���ѻF���x@ґ!�	��`�p�#^΄~�HB$TT����
�R�5�rDy�e�N��qL��(U ��ܧ�
uɣ7��\
uqh��D����3JUt�����O�[�p�H1���4ፗw6��1�߆,�B`�L�o!�gJ��n_����}.������hS�3��Y;wA�i��JW���>A�$~���:�-<�~Pƪh�0⾢Ədsq�0k�Qھu�P�Fx�1��vԌH���$�+xw�=��)>U�,�Q-d`��ZMW�X�!�}�`I$뽑C��n5Ek��D�!��FF�&#�sW����J(��,�����t&۹�։���'4�Ɲd�^��}������`���i�{��Y+a����H ���L�[ca[�H����������b���X��<�n�'y��V��R��T .����1��@�N�u���>i�;�z����X{���L'��Yb��=0���.�#�V���|v:��X#���p ,f��@����`k-�S���q2^�8��r/��~�Ct�S�᱾A������L�SRS��REv�\���ٜ�E�yY��ؤ��������=��n�q�y�.(T![�G���m���0���椢^����ORm٫�3����fg[�Vb�����C�	c�T2b>.A|��E���Ӟ,�۷�m������v�
�1؎�9����]ka;z�G�#Q+:ʲ�Ee�F��!�o}�??[yǆ����]�&�u4��Q�n-��o� ���Ӟ��A7A��T�D�2ڋ8��c��~v���|�l����JS���aɷæ�rѣ�s:�^�T���S�/�~rD�����W{*ve3.���b	#n�?��޼A�Ї���=�⢣���3�,&�l��`�^mb,��d{A��-����W�|P/��;Z5���E���|.�
x���������$�&gw`�}ڿ��~&7��c�H��OK��rS��,�L��rI�����7�5�vFY����rcc�]�K0�Q��:�<����ڡ�:���x@�����`�W�K��.'��"]��qΗ�;{��BV����Z(~���<�7�r�oۥ��AA�)^�wD���+��\��(�$ǩ�ye~p�n���ě���|0d�t�U���-��%l��u��hȈ^�.N+�S'��
�-�j��W;����w��{��ϦO-��~/��}Bҿ ɰ���2����j�ǒ��%��t���w]��A�ɯ��.�� ,$�aH�A��g�&��L2���L� �	�v�{/g��u~�D�!�kZt��BͰ�����T���������B.�,0={������O���3��s�v��.�ƨKl	e��B9�&_)!�oA	 �O5"�^��OD ���&H����?R��q�iz۩�u��zh��,����{8Z��Ia�lN�������;�8G��\��O���>���8���X�F:�2��y!D^5��]�� ��r�sR%�uK_.<�֬|�(T�_���e��(v�1B�
�w��A��ڷ'�,�_��}\��b��(r7�m�KP�?���g��瀤VÌë�q${���ׅ��{	�II�^V�r/	x���@{�K ���'���~�V4I[~���1QT��wd����C�c�r�����-rD�9&�'��@~׌���(�L�(Aj`I�ǖR@���o(�=���3�?��2����BP'S���q�J6��}b�u<�C�"@𡐳<KK�M�Q%���~��h�6',�-��d8�3�lTBcDSw-��o4��C���3q@�C�	��/��-}&��I8K}�N��ԿP#����݊��N�����[��j(��[��3��xiU+Cx$��05�p�t�v�=.Tg/{�~����g�7�xЍ�4I6��S4�z�#�{��.���eliJN�빙m�)��u��#5{w�9�������3�kcs���{��� 7J"�l�غ��������� VM.Dt��)+��5�T�9�]��+)�v�1��;�v��F}D �SmA%׵�f*v28��2k���X����"W�h��ݭ���
g�@���ܟBH<�t@_�b59n3�jHB'�i�.p��1l���9�w��o�$�{�?� �P�*��g�]-��?��.P�s�e��eC}���Z�#���ݺ�����'��^qbgm���}t��Ѥ��9��3�.�"u�$�Տ?������vP�y��>۱jq1���*�|��|2����f��e1��N�E�a���}~���۠���(.�)�6�M[�e�%�tN��gu[��GҌ�t(�#T1�mҖ��"�����y��^B{�Q�7/������*����y�����5n"3!���B�h��n
.�#Y���=m�'
 f)-F#���8���&<�d'�aP>�������@@��=�����������MP�ۇ��N��>�swΥWJ����m]3��x�Íp�~�v*Y��߷=Ô)I c�)I�=�>RwZcs��D }$}X�!{O�zo	�j�#�v[�M��2URJ��-Z��6������+�iQ������6"&w��bHt�6�+J��%d;.�	QԒ�`0�~#�1��i��<V�V%(KP�gA�����Y����N�&Q\��o�{��c�B�1]) m#�Iy�oǢ�	��d�X?��Ȯ��/b2��`�d�IFq���k���A<Z�t��F�X���������a?|{HCr��g��*t\�lw���Z{@:����H�6��ubm�3+��F����z��a(��0��9�m��ظ�4i������<Jai�����E�GÞ�s�So�8���:%��Ώ��2N��#�7lRy����.&1�<ZD���'�zR9	&�M�s��{�i�F|�U���j��
W���%�Bx1g��ce�I�{�m��*Z�Dh8�5��{J�0B��W�y�����@F�.H@s�1�l���IG�/!�%�a���������O5X���^֝Y@�F�Ʒ���n�	��f�]H���4�L	.�b����^GA^������2]���|�b��;�I���QD�[�����7��/ഒ��� �γ��A����X\JJ�-��%��=�+f�G�L�uqM4G�<Z�w;���.��� t,���]7�]q��kN�T�J�kD5��F/CM�C>��fL���4r[9#C�ilt]�؎^���1�{�ˣ�O�W	�m� d���g�>=�`�YT6����V�
�L��2�M�#"�u�[B*!k�\ % 6��o(l�x�ޗ�'_�d����vM�[~6�1����WJ�%8��*v�A���弹F�72�;��x��lQfs09�; e+-/V���DL7��r���H��}�����9���3�	|6����#��8s���g���?w'#���s��O�V�ɐ���ٽVZo��]�n��R��E6����>B:�E�Y�w?�,RZ�Us�����Uc����D�j� Y���bˢ9gЄ���,�D.<y�EC��7g�WY4��}3�fEL��Ӌl��G�%�#�+�:.W�裂�K4?!GgGy��s�O�S����ԟ�f�Bu)�1
X�Ss��i��3b�Z���:��B1�P���N)*������՜�y�}#�K��f��\��)�A�p�r4��:=�R\��/y�˙������n��ľ�24�x��}3&�����usn�{�u��ع;�eĪ6����+I��~@V����_�+C�K�SH�Z���
߭���vs��-?N�kr�v*�_�RqX�g$��F�d��!��w_<�7r�bfc���>i^����l�>0i#�b�s�C��'匫�����\Hs%))	�bd�:��2#�z���j@�w/��������M"��:�`rȾ_�#`Ue���`O�����kˣ���6ۜ�u�Շ��ŀ��[Ǔo?������Svl�rc����9(Y��'���7'/&��Հ� ��9�\#��셼h5w��4+�52N�u����1?�������v/N@T��]Gi�BR�Ք�����͒�+C2��X�=DmLݐ�$@V_M2�i�5�y=	�Q�E�@k�$���~묹��K�E$�a^�V�1T�	��,Bδ�M1˴a(��,���s�\k\�3ҧ��
��ed}0����R������������xm��0"s��֣='��A����9ܯ��:��'�(�$n_�`ya���̷O��]�~Ӈ���֎L�?_�_�|Es�9(z?�-8��ݐt���J.>
ܲ�oHT+��Yw9ˑ:��<�|����<*e��Qk�G8��8Ғي	�ӷ��cBG��<E������5������r���hH�D0�y���^��n��NM�hwM��M���r�Ƽ}�٨Q[��U�,��L'_r-c%8���ݤH���-�8E�>(zz�U�_n���H��t���X��B����K��D��G�X
#�!��x�66������BMӝ�{��~�]ѝ��[����_΢?�D�y�fӢ�_QH�����sǣ�����C���E�� ��_Mh�z�F��#��/���R���C}��v#�g�Oh��A�U��PK   :�-X�L�,� o� /   images/6b34e9bb-e0d8-4181-9662-be6b7300858d.pngl�s�%0�-zڶ�i۶��i{ڧm����m��}ڶ��}�֭���I�Vv*�T���ΎTV�F�Ǉ  H�2�  $  &�$�w��?�����f��  �J��{\t[�ٮ��<	�/�2�C��"G������C�@�Jb�*�ȱM'Mӽ�_&1�)�;dc��.0S�l�Q%ÆDE%�b�$g��?��=���W�����|潕x�)}���|})�;�ݺܺ���U�c�^����W��Xg��P�_h��1��8��q���/���F������Ai��������?VXdZ�����������u6���7���"��d��p�@�l-� ������9�r%,oM�?.L�)3�ͤh�L����!�H��iۜB�%|��D1�LH&I��e͑�qe��:�%�H{�%�W�Wz��ꙺ���**C�ɫ�~�T=wI-k��/7���Ì���e)?#)<_n+v�\n�j;�x������&����Z��~��mઑ)d��U��۝�И�ѳ�<-�x���]�hS]�-��J��zx>������T�H���K?�v��k=�{Up��p����S�����M�Ae�I5�ID���5
���4u�,h�G�uR)�?HQ˔O��<�n���4H.��l�����IbfZ �(4�R�*C]
��&2��*u��
x"3��M�o��}릊"_Xl����a�2����A������/]�/��M*Q����?���(I�WCD��� ���Ec�o��kr>�i�U��4��~Y��yެ�U�FCRE�S婱kI�_z:��k�mA]C=�\!�8o��mU��[�B�r9�Y�BQ:���	ċCT0�YJ�8�]�%f��f'��T+�j.B��A��h�q��-�ApL��Q�%c��d۬��@�7X�̈��D��e]\tp5���VխwV��+TdO���m��T�����0�N�=�4���4؄���bS�}R�ca����^��_[�:�V�_�:,�l������^��e��s��ڊ�#\Z�����{�Z�{��<�[����Ϯ�>�H��1�޸�Pf�d���S�R�-�ȱ�իhT'��� ���e�B�C���L�"��Ѧ
���2	��� �$	�XU��@guIץ$E�✒��*r�?��ֻ^�v�n�ȱ@B<�1�J=�� ���gn��)�Hq+��[RE"����q;A���w����O�YeT��n�5i�#�d�����{]���!>�� �v-�i�JP���F�BRH^��NTRDJ!��R[��<﮺�5�&����d1l��x"eq�2�iYK\}Rj���5*Eno��"����>�k$����2U�X�)�PY����m����#�OB��^���jUU��3������=�L��($�*+�����,�R���6a�7�9�b��/ӮG��"B�����ū\�v�z�-�Ӝ�q�4n�$���kMQ-�9��sz���V3�-%�ZjYE��1�A�kc�æ�:��Ovy��dko��N�#bP����1�>���+��	��?|�x���N���NeP�����u���4��c ��ף6�F����ݴ��+z =�%x���Y���L�а�+���^�\���G�0vЯE�1��`c����HP���2|�}NC����~g����� ���b��4�K������׵Z���[n��R���L��ETӗ��ЙN%���"8���u��t(�o�����7���J�}�����׊���p�8�]	M$�D�t҈&6ڰή`�#ިL#.����%�4���:�q����}�'E��d��qʜ��69�K�\�!�, :�6>O�?�|@��JGZCw�C�Ġvte��A5�C���v�����ۃ�W������������?#qW�{�]���>�[[�<բX���x7�ퟀ������t��؏�x�w�\�o��{O�S޾��w�(uϧ>Bv���6��`c�;8E)�N��Qɱ�X��}���OX377���,�Kn��zDZ-��P{&�aQ=�&6Zc/�c��q���9�Y��f�����_
��h�"������ۮ9�Pz���?L������V{WG�\�Kȗc�Ê�gc�aIdlS,H2��~�nw���v�a
$]�IJ���*yg�0F�j��p���=��lu5 ��������JA6;�-���$�ʵ�p,�,�b��&=���Z.�K�Z��*Ö�1��X+�Km�vRl砯`��Q5Îf�`�qY�5)�io9r�Mତ�>_�Z���N�D}�aC[�$���UÐ�M�͡��F�8G��[&sV��)lr� mJe�&-l��9I��b�ֺNV��]!�i�S�sml���%͚UY�չc/�L�b�lAos�9q�^s-E��MS9-�
X���i�0�U�	@<���6�d���L�s��F�{sŶ�i�tT�5��<>�"��V˲�Ȉ*M������Ql�^6&���0p�G,;m.��>EA����:�F��
����T'��������n��i�_�}nl�Ñ<�\�?�f��<��/54R�~�^ϴ<�P٘�Ud+���ũ�Y���q�۬Uw:^/�
�W���[^_�	_�=E����޽��|��L{�Ѝ�@U�R�J�BgQ�,1����f!�&��D�Y�h�F�MNc������;��������|F�&.#p�� �(*@X���0�a}��/y<i*�7�{>�z<�2gϜ9����&[�
./�B~��v[��T���`O�aac��H����R���$oHY~�(���#�뱈��i{�70`qrK�!��$��./bR�E��|����ndp$ؿˀi�����P�O{6@0+��(��iW�����x���D�w� 6�� �)��U�dl��e�c������_�F_��Ӆ|�gB�R�wx�@7�����Aϡ3����C��ځ"x��nE/�TҦ=%>Lf�X>��r�磍%9��F2F_�Cp��U4�zp�j~&�P	
peI-�^����ԑ�
B�����v����4�*��!��'�^*P�y{� @�8xxΤ?��ܷgMY8���v�G��?�����nyw���E2E/��p6ؖ��k�����D2�L��-��l�T\��6��3͙��g=��`Z�5cw��
[�<��pb��GB��?M�KaM�ڵ�@oeں�6s��\��EE^��V�:@�1��\T��òg'��v1�gt�d�m#eDx�>`h��k�;*l&����7�jL�LD#b��k��������ga�s�봘l�3��%z�U�`S��WSJu�_�&�F��F�q���{�'1��9k�/�����/K��}�y��?4E~��~J��ߵ\e.�E%:����r�W���։?���ڹ�2���v��N�-���g���?�V�gQ�.~QB��;9��ݎ���oUZ��
��8�� �<�g���!b�;����Qfq}�;�_n��w-�[	�9�r�&"�009ӂ�����~�	w
͐ma  @�vI�� ���+���1x��퍘M�������l��#"5��6�0����wj�H���ؾ��,Z?��}cF �P��qZ��Њ�]7����2����#�4-�?�!�WF"E|�S�f/���u�>$o���ieaZж� -[�ʸ�����D��l�@���F& �����Q��p��}P>�[���$�x�C.X��2;��96�N�
QQ�a��>�cpg��X:�a���W�d�XN�К]/#��/��:�>D��v�?y9�ZɋMsX��I"F�o��x@�e��\k'1uK�2��}		<������Y�x����:2� �p�JeG���s�<(=��a�!���a��΀�ߞ1��rGh#p������A��Ë\���\�d'&�b�OX���拳�ǓZG����J#�«r���©)W��X�?�<kQ��a+�V�U�m.u�"[a���p����UF,��/�;H��h�0��d��k�kAe�T+\˯�p�[�����,��<B�u<�՗Z�'�>������o���Մ��A��E��-�KG/�WA���$�K��~X��x)X����ʦơ`ϑϝ}x�Yc{��КZ Y�h�n�sE�҇s<�
�KU �
�D5����]#e�}�9#>5՜z<Wy��k5s�����ޯ]��u�Թ`�$��G%K�\QpO��!u�ִ��g��SA^�M�W��s�]���/[����~�wGs��^�=(�w(�+����R�)qP,�h���Z�͟�"�����
�٤�F�`��l�:�"8���lF��0	FP��7+�Y��>�[$̉��C���pJ���.`gF�R����n���s���l�|��]�u$��wt�6�ɘ+�NW�{ �|��߯�(?B��o��4L�<��;���͝��`�	 ��B��o`�-�V
�X�M!�oR,���$��D뤣,�5�_T�0����d���sy}�l�u.�>�'�Yd=��X��'��w�qШ�G�E?��L��
�}��4�Y�?�ά\�h	K��-���z�v�>pA+b�*H���n.�
l�F'�X�&.\�*��Yoo~�V���F�=?<�w3ǁ"0H��~�XR^t:��;��҅�$yc���Fn#�Q\,�~36c��k�n���\�H	� �ѡ3�1O:��W���ī�2�t䓒���V���K�b�� �ݮ [�t��������=N���4ʦ��'p�pw��&�+�}S� o���k����ɕ���܂��"e��!녻�і����P	�c�y�̐������,�:7��:{�O�ֽ�Ɯ5������L�~8JY�^�[��G��{ w\��7�ֵ�%�	 �_�w7�%.�y�ͽ�c�����W��f��n��V1(�o�|2$ʅ��M1�<���V�Q�v�.���>Ә�m;31��s<c��X�n���N{wE� �<3��TJw؎o*I��r�7sQ8
�]ߞ��B�/7���Nk�|�&����E�zߟ��r�.��E��Īb���a,_%g�Mh�ġ��JE��n�iϯ�Ks'�|Bx4$�������ml����J��$�ρk�l����ZT6�������k�Kg[�DBI��<=m�3SI���7�g��H����~h2��u�!7\��Ԃ�0qjY��X�̽��ɔ����EO�)�� �m�m�"��'�����,�;��)�Bބ���F =I��
}�,/?^TGh1*����"(Y~���˽�O���}�Z�xo��2A���=aO�=5����5l�m�}ƎZe-#kmS�3���'�ꀝ��d�� �5��,&��^j��5�@:5���f[�'
#	׶��0����T�!O�YUwe��y>��j�흩G ��4s�vY�F>p����������S�9���е#�An�bL h�9"�GR�`o�%%&ꇕ( �$i*Z�M�.H;H��B��7B��`��ӣ�U<%�"�WS0�A�d>k����X�Fs��D����z$!��LJG��@IL�9X*lU=xJa&0t�� 5+�tT�~_s�^�$�>��NUZ�q����Ӱ8��=�&�P������l�Y�/�H�Iy�:�i�� D���߁ف�Q�EVx&&*� �X�^�-�$sH'$i8˜99{�7�ɨ�����R�*�\C�(l��H*.�+�����e��1�	A�h/�S$΂,{��ޘ��|w@�э�̍���.D+�f�i,���+e��Α�X��ܸ��0嘶���to��v�v�`��AN"bVx�4}`��Or.���C��' �lú�5���QOGb)j2�
yN�ܨ����8�jB��j���̡�K�����s����C��e�^����1��L+���ؗ�澕a�w���gao�>L�kΩ�6^1:�
��cVRMA�5Q���x���5-z��𨿨,�j��՜x�)�G1I@��2>_�n=~ߖ��苷���/#�?�(#�&�r��|6��w]�4�w�܃~��О�.�KܮK�~�/g��hd�v	�*4��I���+T/Ȣg}�u��+U؜���a�=t�$�۲��MX�N��]M� ��A�H&F�0B��u�5K���6꽲96����xF��h&��>E�&�����f��N��c�l��t��a��r��������T�>RRҌvaHȣ�,��=�Ta�@���{2�#n���z�;�p�Q����'�Je6�XV��yC4���`�����~�|��3?�@i��k����I��WR;��`f>���f>��_Q_f�����_R���LNI�������ɕp��{���<�w����Ow���I��s��S���<�]��9�X�sh[�r�H8�6�[:�	G�U+C�mB/X����7j�puu,&�M��ʐ��x3%]���Ћ�^�f�r�� oS�T�D�|,(ٰ1�!r86Ҭ�1	'�4�N�g��r���҈Zj�!�^,,���[""�Pˇ� `�u,��61�����[и�5�����~Y*���Ime�'�B�߶\D��c�S��4xڜab��>b8G��l��j��&������e�#���6�tT�� y�aI(r�4�ۍ�g65�)dbS�;�>8qe�^������m�����~ 8^"^���>+�H7��/)0�Uy�˨��#\���:�D�щ�i�'F�C�ǿO� ��I6�!S9�O��T	zh�Ҝ+�m',;�q�,cCw��I�CC����@��7�L�tn�-��1����i���N;����D����]9��g� s{|3j��s����7��`瀱|C@���} ᮳�KW\\ܪ)�3`�nK2l�8M�\|b>�	%�R�&b�^��*����=���M��Ot�ʼ�n�(��Ƞc�.:�c2"v�L��#�Q;�!��`{a6FU���&;�tĪ�=�\�R����Q�﹕�7j�W��}C����� r�
L�F�(��v������z�7�.{�d["�%���I���6��y���m1�f�T��+�š�n�G��t���Nk��A��ټ� �r��MP���o�V����86X�Y��K�J����.�\
63��� �z�v��f<�Ƅ��ۏ$�|ΖK��US�F;����g(�#�^mz�J_i�E*����y��j�=�ژ&k^0#���X�u\��Lc��#�Z��o7�7wf����:�-8��B�B~X%~"��A��yΊ�/�"��8��{�ۋ��xO W�!	�ԑ�rϤ�s�SFu6R���b`x)W���ilT���V�c�c������A��޾��}�ߟBx'S
�Y�����Ǌy�ӿCx��*g�g���e���瞤��O���1&4p�m�r�}υ=ϯ�;��[W�O,U�K=>�_����l��V\�
�C.xG��5�H���s��㫻�n��%�0�H���ϋ�QD>�'���OB���`���}�b�޺�K��6U��<�I耒c��G\�o�\O�5��a�F��. w�#mL�����ݭ���(R�����V:Ȁ�.��ՠ���:c�d��8��ujȿQP8��t�6)�2+��S!,t}��c�Y��l��8�O�</84��X��m�z�z��W�?�9ݤPX�>�!/G"�$���}�ģ���^�y�1 B�B���Hn�NI5@5���aT�"p�)=�ǿ�G�������WK�f�l
S����|��y�T�����.�8+ C���M��c��#䰉��V�e��M�{���[�D�bC� ��+
KZg���H�S���%�3�b� ��XƐ{���߆��i��[�;��eÏ�@�=����/1��ՏQ2�N��Z����]���U2�;�D{M;=��	*KY-\.;�Gx��l��X������D�P�R���� ĨB��I��eø��y��f�j��p�	TNf�8:�O.�TP!ъ%�����z�2'��:������ľ�G���9�����B-�����>�a�Β�Q�N{o�_�mY�c9+�ư�PA��	$Q�-�tɀx =�Cb������Z�����g�����CǊ���L�9�#�O���^�O��|Ɍ�t�j{���m����8�]^���g���&z�u��!��HSƯ���G'��pv-�bqi�4�2�硫#PCP��)��ʘ#�Pf=k�����z�?	2Z��O�Z�d:�a��6ȱBf�NΓ'��P���)����@�5�O�p����|Ya�O�?�C*�xuLp��]{2^���UvN�}�[��A�pF�2r�E��y�4�0Ȭ�^<�%�BB��&��2=�і�앖Ҧ��%:��Y�aS\oo��Z�c���g��!\X[  ���3,:�{eK=�^�d�}j���Y��^�f!��?cL���*m}�B��O��l�`.v����O�1�
�"�H���j6������6���ԺԮ%2�-h�dI�A���%VM���`��a�����t4�VҎ��{ߐ3��oK�C��w�/�OC��n�?�&�w<N� ���lv|�E�v��^�BĻ��/��5x�DCl�!���$A��g+9�Ԡ�g�S���Wb��L���Y�v�5�7���<t���8w�¬
C�4��tG�GM
 ���bzP�JR_�Y���]�ˤ?$�o�2����%O�l���q��L{#]4���������ޕ�GI�����|�XpMg�z�^��k�u��r-k�/�'�q,�57��1�f���'�K"�V]0�ߙ=�n�KYRfG��Į���x͌��5M�K �e�C�K�g�Z���k�F1���+�{�׫?2a�W�\8ͨ�Y!�b��TcF)JadS��Cc��a��'��7r<n`�#=J��$؏�أ��K	��/8�b6 ~�?�|��n�ĵt����tY��������A��/��{���m�<j�5�I�tEpZ [��)T�o�����-1#]:U����_����Dm�C���7��t��i.?󼤙�)Q���+�~w�t�z�I?����U�.i��\:�o���v1?��d�[�m�� �5G�@�g�������ɭ+^�I��H�w?���;�y�$t	�ONR��X���j���=��)*��}�1���������5��C�����y�Q�!"�I�� VaL��C��OT���7�=&��~��yf�,�E˾>p��^�zyE�`�O�?C��'c"��P�q��A���,LCǇIq���ҳ��ic��#ݔt��t�_��93y�d�<g�[/�e��K8�ݳR��;V{��{v�Z���k���^(B�r���7���?S�_j�_��%d�#��q����#�<��|Sa�	�P�?��[B�5�a�E��~�ĽE鈚�6�;�I��b�̽��-��7?n�7!��<��`vI��۵E��]:FM1e��x&�>ϟ����������J�ϐ���2�aخ~~ɒv�P'���`zA^18�q���J�B�;Y0���1���6�Ȱ��{9-�%�k$;�sr*#��5�>KF��L�5?�|h�����	��ǃ��[�H��V��a%��h�-2Ō��߂����������C�+���i�8N0���e܀k|}C�Db�d<3�g�p<�Q+ I�� `�0bۧ}����A<�@��{t�8ࡔm>o��[@�5�9���_��^���}�=�Ad,\��	��l��d�����I�{���	�b����0|���e�|��.�}��*#7df�[*F���^�,7vӵ�������LV映A�,j~7IT��tX�$(B~TZ����Ƌ��9uǞ*ke���If�>��@�ҴUu��G&�PYR�Qw��]<j����	�����m���LC���7x�fk�u����8\������B�ݮ��kV��9L%�C6�<�=�;[��(_0�6��'|�E�"[q������C���ޯGLqM�*��B�/ �������gR��AJ��v!]�ɼ�	a��kn�Y@��SZ�JϑZ���� * "�Ӊ`00�j��'M��� '�~� ���?�6����6���6��t�sv�9'��	;+1��no�=��(�CUE�Gt	Irc�{~�ޝ$?�[X�zd�p��M�7e���u@�Ol�|�S�� ����U�����{8������gv�"y-���e�idT���h����`�M��{��[��F��W}9�,��@H��t����j׃��L!�Ǹ�F�%���pQ�L�/�n}H��<w�q-G�����[�4�7V>/:���z^�"`�k��z2�;�#�&Cn���q�%�����I��6�	�Y��;�c�!Z;������[$	�(��B�}��i��?Hm�x d�{�e����F�x��:膦D��;� z&I����Ƀk����~0�k�R��(�PV}���������i���d�@�������M(�M����4��_9���!4�Ş�t�#���dpȿ�����Z}�7�;:������FB,⟡
�~3�N�,a~gm*ZQ��_�����G/�$ѥ��:�v��F� X�0���a	-���H�T��<Pl}�F��b�1�M�h���z����|�Yek�M�Y�rm[�xNЃ~��uɲ��[I�� 6ۘ��1��T��kb���x����wtX2Z�y�}��bh���P�z�A���N���ӹnfrg��� ��g�Eʙo�Z�P3Tk:œ��[Rz2W��g5X���H�f,�'��f�(�d;*��5W��MG�{������箣+����ǇJl��͠?���wJ����u���?�7G������7>�Hq�Iv܉�Į�]� n=eb]�K������}Ut�w����<����|���;[���D��k/��V@�^����{:>���������y��
$����E������ �l�#�8C,
���t�p�����K�rQpS��<��! �Xi"��|n�<Ę�;d����s)���A�����)h6,Y�����$-
�%.<�*�4��)ę�t�$�Pw�ڌm�ｂQ��/Ɖ����tUbf��w��]�&�fܮ̦F��v���Wx^_�ǯ����^]�"��EcUA��#Q�8!ajj�-}���kޝ+�T��f禼��8���۟�.�����)�{ ��Ȟ�!��r��˰��������,�Ǔ�73)T?�:��E޸�):8��A]�SLy_�)��_;��y('E��wg�:�Jb�N=�A�*@�Ρsԕ�w��*	�d���Eύn�h�n��L�̏���^GC!�.���w�JY���\��h��K���Z#2�'�py��E���5���}1��g���cJ\d�?�0�1Z=`�g$V��|�~Pq�}x`��^�%���֢��=��S�P�v;O_���u��S�ʫY�Kw�
/��������w|����d4��W(�شV���5�ʭ�/ߔ��AǷr~���O*� �P�v~��7�Kz���D!t��H��z�z��8v~�tĕ=�¾;;�r%"�����ɟ�(�F�[�O����ԲB8]q��T���c�=3�!�Pb~�b�_�څuؓ<8(�d��&��o{ѿ�]�D`u��]��c�$U�9	B������?/W���P�U��OB9=NV@}���)�
=�|����]�<�q5��%�Ƕa�J,o�a��$��h�,���|�[�|o|��)��2�]�Z'���E��g��b��$�J��{�}�:�[�BWq!�55�H6����D��:P���3��)��6
� x���H�`B��<]0��/�կ����[Xfۭ.��;��ҝ�$��k}�r�n;�����~jXA�;��v�1V�"U���j������*��V�� ���A�8�9�	h%|@ã�O �5��Ob�4yMa鎦�=�3,EF�t3����w��e��iҨ�	k�!  �)�㡬,�+� ��r��� j��T(|lvN��=��E��l��5s���1��)�awE4���Fw��2YϫZ1gt���M���\/�
�9&��z%�W�gV�P�F���Y�>X�߀����
�����AZ�?i��z'�����en��Hf&�
�\f�M���i�U�$��*�/���|TF,�"$T�V�"�ڱOX�j"7_y�{,t(���z�J����?g����\�Au{!s	������+) #=Y�X%��=�佦�O��ջ�>#�GLGk:n_�:��z,�%񦲩7f=9$��HAOL���&��m4��-?�%�Gd�5x�oy�� X#�Z�>�n�y�C�h��*�<����8�0s��Ui2�j��z�c��R�?��a�z#���g�[g�l�+ �mLl�`h^lQ)�V,�x��eWp/F%����WxAD7��Y��ud�N�{�-����D�a�.�+;�ُ���u젃��>�ټ.󗉙�wo�E3����Î�9Kr~��q>�ݍ	x[7~��j}g}��BY���]��OW�։G��W�W+$����J58�4fK��N����ب�ɛ�J������Y�j��	����9g�u�Z�$�j���J��TT
2��5�3�-�ʤY�\�Z�n��n*�MF�Vx��Ul�qQ͌��uבc�K����qy�K�Vl7u~q���%I��E�%}��W>�hn�u4 7�j6I4�F����C���]���O�o��޳�:h^�oyK�oɎ�z���E_��$�/+�'���b�]�}�x���; L���.�]U^<��ǆO�{`Nb7��oc~O����;K<
�I�f<*M��u�;Ke7F�r���G:l�M[�$^��'�$>���`ɁTj�U�Yit?�lռ���|0�
�>8�-e
�	�xbA�� �S���W#i�;�"�� �,��� ����n�jH(0��^��y�=n��`Z�9n�`r8>�����[�c�W��L�nO�Gd�pH06`<4-Ȕ���8�/{*��ǀ%c}K9ܯ����j%���Ji�:�/X��G�4m���ABR)�_�U7Rþǜ}f�k)vz��p���3}�x�7�Zq�ew�U�c82�7�fy��$�;�M-.g�������jT5�ޖ\���|�,�2[��V�����dՎ�B�h(�ֻ$#�F����5���Љ�Ԕ��e��5_'�e�4�r�sĀt@�Mӏ��Rz+�Ty���^l�j=)��V�P3�%C�&؄��������d;��Z����yɼ|�6Yyz~i�����R}�U*�[}�xs1���C��e����`"�>v\��%}|%�2�@�6y��#A�Gѭ�2��2���4j���:�I�'�'�����J:�� �a�A�r�4m~�՞8��������9N|h�� ��1��Y�����g7a�sC�߿����c�Ѻ�X'|��R`#��{绖38����c���}��b��9�z�����,�2�!�?����R� �*�201�0�d� V��@��>oje�(��s�\�"��Px`�J�4C
\<koR����i$	����']a� � ��č���"|0���7v9��Xɮ�j���A���ɜX#͖�{4Jvz�5��y}��XM��fT�q�L!��z(�b�.k�����=.��V7�Țey�wr(N��ƒ/~�#3#{H�x��F�Z��ޖ�S�K�$T��Ş��t#n:��A@/$r���)�F�9�v���������2�,�j�f{Id������Km"K�r�:m�Wѓ�"_�!���W��ӊ�����=0\��@��*�r脗"�����4;I�L�P��\|��fь�6N���7j��%�ɨĕ6��N7�Z��rYWE㘹d�dTwgښݸ$.W�'L����o�A��2��0�_L���E�֠c��Z�B�B�W�@��y��F	4��>���|{�ҝ*����X2�P�����,oY��PSI&M'��_�Y�Ww
�r�VGhk�U5��B�ߖ���)4�ja�݅S(olKc V@1J�<���ZRS?��+	s����Gޚ`���u�Z�Npbx`�Zs�ȨezcEc�c�0�|�����kJ�q>�X�=b~b�Y4�:Q੊>�q��~a\k��Qc���u?'ga�|�c��5i��qLj�����V��U��`nJ�Ҳ)r��X�@\���f�L-�l���+,0�Nr��|o���������|�ǎcY�*i�	f{(�
g�KQ��O@�IsxQ��nYw&���]�mჅp�d"�Sl�C�W�Ǻ�0�8Q�-��g�^�GZ7�!�M�UXi}��`Vq�6�!(?;�eʣXyc�	t�/�X!�r0�u���g>����o�� }ɓ��ްSG���:����	� h�eH�k�c�6��2lkRɡb(k�5�,�ᬾ��,l�Ϝ������D��^�&��l՝x�y��>9D��J|ӘT���r �Ƃ��̽�[�}:Ӝ��7���F�� D�A-[[��K
ʈ ���}q����%�9c�ׅ��2� ~p?ʺ6�G�) ���o�V0Ӭz��P;�q�/���O'�C}p�09��8)��R�܎��n�]0�=��|įF�}-�C�"����4���.�Q~�{Z�D�m�i��>2�v���CS����i�g%�*��(<�M�&��@}�@�B)H9��l
�9���S�l��\1��F�Q0*	y9Xlr�χ������Qbx�y w��Ve�l��
'&�E�������Y�fYF"aR�?:��� �4	\��'>]���y���!����oTՒ�':���y�|���ݡ�"]�C��T����U>� �]��Y��^O�2`W���s�k~��Ӫ��w�7��0�v'*&L�m�<,�tb�<�O*�h�$�i�X�{�#'�d��/��ig�<j��Z_1x��Ǻ�����
<t�Y�RK	�
�B����F4%���z3��a��	o�y�r��6d�O®1s$Oy�R$�_���7*�����$�<�%O5<���+�ϛ���J�_�V'��5��#ϴ�qcޫ��d}�2�X��XT�f=R,���A��0��6����<iƱ_�+�T��(����{��"��	��䤂�ʨt���2��#�{pz�����A2Z��Z��`�G�
*��2�2���%�s�a@d����p���Li�!��A�71��U8ր������
�����i�p(��?k�e��D�@wSRRѸ擫e�qH^H�Y�m���o�c��[��y�����Zw*^]���ت �Q�ЪJ�3�SX�q~*����O���E���[oz�X�����h��'�$Ȑ��e�[f��PSr�����2����"S��Cf���]���ە����b]�PO�!Sm���ڑS}��L�=D��qAs��5��5��ɔ�9��3����,=n�ٟh�����k�@`l�gR���wh���?�Ǖ������l�>��ާ�<Ⴏ�.T�����I!���3:s$욆�iA���TD��ʾ�{�Ӆj�9������"q�M��ͽ�B�۔p�,��8�sw*MO~��a!9ES����p�t:P6��� >@Lm�pAY�=&�Zft���# �k�(J�E`n��x%g�K����Bbd�Y�FjLԘBj���T�U���0�Ǎ�$vSX#ƃ�ݔ���ҜȘF����M�;�z3?�>��G����'����Ҍ���b����`��?f		��ܟS[�;d��U��^��4�VՖ�D��$57#�-;vy�x�k���;����+٘��O��훧��h�8>9xp-r eLvm&�f��=����0�!���狞K���TO�<�WY��mQ�6-�9��Y6����X�^�������U%'�9�{!� ��%�`z��Rf�r�
�|��� &���n���\ �]�D�%��Z� ,P���(�*!q�
��(�r�x��:�'�^��܉Z�4!:����[#DD��e�6�}��O�
�Yf�����f�lUl��:j�f��jTrt�Ҩa��$�Y����,u�JF���_T���<����7�n^�3���B��@����3B��.�;r�V�B��c�Z��'R�%�'瓬�]����!n���g�	R o������lP�E��e�rF�
m �f�)��X���YX�%Փ���%txp@�1IF.�0��0�LQ�=(p�,���p����O��C횔�~��a��A�c��u�R0���-�f:^�X������LJ� c�>^�+Z�b�s*z	�EB�;��֭�N��dlx:�� ��ƖlB�m�y�����:�s<����3/c��w�d���2���oX/d\��>�/�c��~�DQ�Qǘ�����=9[�v�b��Y�8�y�:״!�B�8R"s���1���xko�� ܷ�졨w���d-|�_W��r��}qA�C�<���}���v<�P3�W)C����y��k�^��$ԅI ]�4���6�i�Ϲ^�ĺp2$6Iz�0��1�6�8�26P��H��/ �(����(����3Ħ���HӔD�n��AA�~ϝ��Rw]8O���^:��Iyө�u��\�Ѱ�Ӣ���!����콡���Θ-��NbM弡�����3OPC-�kz��-���O��{wsoq�(w�b�E�k�m�D6�3�!V��#O�t�8�lc��DD�Бr1䉶�q�A�P�Tڵe��^���_~�;?�����x����z�	��/?��������#�{0�8M�,�lب��Nǡh���Y ӂ�E���ل�\������7���ȉ��1��gEHӂ�J�z9=���B�����Α�V���sJ�$�¤]���X���9/TX�1��
y���D1R�ETk�>�т��4	�b�uz=q̙{!�(^�<F���V�����j�7|G��u��껰�{7;W����~A�@޼��4xm�nehB�+8�U��C���V�`i���o��yس���&]�����i
+��N��
qv$9>�	��b�Y��cZ�!K�bJmY�1g#���bB�w_����來S۔)�Â�\�J׮^��W}��I��r���o�bt�� �.�B[w_bm�k���\<I$r`} �] ) ky�2�$"=��\t2u�Kr{�b B l ��k�DD��Kp�z~̇M X�%U�#�D��|��-	��p� ��X�B���)�q(r��Sl�A�!�;�\�J���.�-^��YTP��˃�`H�8椀^!@]Ѝ~�U��26d4i�^@����˸�.��8�	y��EپZ��K?wǺ�ܓ�@@
�3җr�F gh;�R�dV�Gq�]��!�u|�0/Ej��0}t����Լ�(�����;�~��䞥_@6���b���i���1tC%�\���C��X��_d)�����Ue� m�P9������%Q�X�qbX�|"<b��4q0>�W&��g�k�΁[ק�%�c�GQ�Po4�b8b�N3m ��Y>�/J6�s!����Dn�g�K��"&����9�׶r��A/�(�t��C���V-o��`8B�w쏘�0�ixwB��-���g��d��}��`�	�q<� �Ή��ᾏ�Ր9�|�X��~jѰ�B�V!.{�����1�I!���Z��1���5d� θa���9�ܣ�Ϥ��q�3������'��H� O K�T��h��d�>;?|:t����F!��׆��nz��_A�~۷�w������|�*��4%S5��0��IK ��G�s��|!P�8�.��CT�9U�	�2�i�/]<CgϞ�5������SO��{4��TS� ���:��ݑ��BZ���1Xk@�00?�} ��4�Q���3����0�3�ktv{����q�4�s�%���9Z�q�]����e�;��8f N{{{t��u~��ic}�F�u��$���R�"�ƨ���tN_x�+�ȓ���/?M7v�6���Q���؛C����@��)��k=�Dا���(�x�-���5���4ۿ���������}�G?����~_rB�7>�����>�u�`��E
F0�^�R��Ȋ��ؒ��O������ɕs:�%�=��M���t� �v&d���iʋ>Q��M�1q��S7���������JS�Q9� =xR�bb�6����`��8,~��Vm��[���A*�f��"\�U���7���l��+&	h}HQ�'���F�u-7��hi�2�D�TX�|��T��e`2��Ӱ^�D�8���A{���	4ZRQd4��c2!���nx���ɲ�� ��~)T#�?�g�1����{���Ƶ��{�:YΌ�?OZV<�T�'��T���c�������s��g���[�Ԍ6�<K��=�A�/���h@�h@O|�Iz���|�H�� ��(�CZ�Y����.H���s+���%p��	������ґ2Po`�v\z�dd���
��bߝZ�����p��B0F0����)��Z�ER����mC�b���Ĝ�;YZ�;��EB�$!H�xK�{�1���S�lyo��B��N�]�]�=[�N�/��v�r�� 0�CPê��|�-�	B�J��ȧ$v�-Xw��t=1|� �ʀ�:��~�G ���v%Z/FTOy�#]����1��O�d˒k�����$�br0k���Gbb�Cpr>�G�Kλ�O�ɨۉ��cl��͒g��}��ҶB��״]�B���>�O6i��3K���l.@�d#������.��C �)����n\y��	���7b_M^\��ڐ���i�1�!a�&��Lx��f%��:�Lh:��Y �_K��~�T��Y�A��s�=�Ȁ�/!>
/6t�������Dx!k��Yxލ�i^!yDNk#::�gC
s �}��W�&&/ �a>�D�	P�*�����4���� x2H�����<��&�n��D���q\��e�s6�=�뺱	=�!�8X�CF)I�,k�����?q�R'�P�8�2W�X�� ���_^}�?)�"���1��oK8Ѵ�OPB�a��4eq��c���5M���aoH�.�[<K�{�k��s[��D������?�ǟ}�667�-���iNv�lr�x$J�jN\U��fo@�V������}��O����҅�b�[D���g���)z��}ڙ֔�=�)���U�9$�>�/H��!�����/h��Ҵ>�Vv~Dq[��SCz�+�w��Az�+�;�l�3-�ᆐ5�	����iw��n�i�`�IM@�ٻWW���G�nޠ[;{,??s�:w�Z���E`�7iP�TD��c���.>?DѻG5=��ez��k��S���2�KJ��T!&�G�K��c=��� Y�L�F�x�<`�PY��
��vB������t��������G�r�/���o��#o��_��?{�~c���x��cR���^�
�kG�-��re�$���)�㜴�i)���<H�ַ�9�:@��9sn��P�%)M�g�x�>�[��ݱ&�SKY���"���q6!L��:~q!�B6^, ���@�?�H���6XU!MLR& \iªy���`b�\�8����k6��E}��;�ã]^�Ξ9��݃��eEA�ۧi^���@7n��x��8M��O֣�����o� h[�= zl^�ꭒX-���$d�g�����V Vd�(K&X ��zt��5�y�:�ءvQzw����D� ��S�z����d�,^���nHT;e�,T�56���i��s�������Ӿ0�&f�G�����V���=	z��C>��%�fbs�ݿ0���v,����y%�P��),�b�|1O�.�Y��e��V��u��,2>��Y����S�.���ĐG^��m��,�!K�Xq���Q����K� �ˠU�J���/�z�s	���c�ޅ ������Ɏ#cT���?��dł�c�)@��y��%0Q4�́��6�����w�{=��6��^9�[C��6��9	��9��\�s�c��J�Y��*k��޵�{}����%'I��gm���S�a	���['����`�$AH��� (������B
� k㾉F��X�y�ܐa#p��	�������x疯BI��5���y�vk�E�N�>́�oث��f� /쇸o�s������ߣ[7whr�1B
 G�u�m�Bb$��4�Gi���2��I���s�"�tb��钨{O������hkk��#RR�p> �G@���km퓍��a��]JJ찞�y��p�s&0��{8��ձ��K�����G��x-���W��X /X�!s%ǅD��hg����
`w�A/�``2�rގ���������Pl��^���>v���1.�ťd(�+@�@ X����h"A
H�v�Ջ�C�1u��!}�;���tn�8F��=�,��?�i����[��V�ѿ�#t�sH��$FQ`N����*J��"����=��c�g�gt��e�#K���|�w��wn1��b�DtX��<J?��E�<u�����Krr:�iYq%n��:����U̗�!c4o��܌6��x����7Лx%���Ktv�g�:<Z���!���'�'��_y��\�Ee�Т	� nHR�v�⢵T�Yc�b��%cSQ�*z�;�F���ҝw^����
?��3C=�8�٣�ӓWn2�r0��yCM�Qel0#���J�OP�+��'ƇWq ��=s�NomSY���gh�}�-�����_~�������4�_��%���o�]?��?�3G�{஻��͂k x�T5U���,x�,,�����v�%�QJ�`�־~���oz#}������4�xNY"�d!@ʶÊ�w?�}�c���)^��Fl�iLI���eI~��/>l�q�"*�Mܖ�� ��w�1��Ŕ����vT���CS�T�3j�9-JE��"EiQ?˩���&��.?�4]��<M�3f}���>E�.\���5"h^[:8���tΕ-5�MQF�l̓	�6*X��b�e�Zq{�,� *p):��=! `Ɇ_����3���s��7Xp�{��v�
5�Sjf�wq�}��,C�&��DtA�2S
�A@?�^�1/�� ዘ�Մ�.�2G��@���w���u��sj`������ <yò-�ʎ�̋.=�M㹄B~F--��! 'A�H�����! P>� �9��� Bֽ��,-�'�ju=B>�L�%w��r���t�������aC��R�O ���!�N�J.�G�1?��/&�A��٩��ϗ��;�u���sK�mG;��ba��_~W��� U0$6H�'D͒؅�� �,#8Q)Y��������4�l�.��N�� +�c1
 �s���Jb�}���{�uw�.=)ᠥGF,���LAÒM,�a(P&������ϫ�[� y���C��g*>V<8ȟ/�k�XQe.t���&	��(	R B ـx� =A�w�.��I��E���!��l��� �m�`dr�τ���h6�����⥔���-Nz���A�.��� �&��0R�:t�'��ɓ�"-��Bk���[3��_̽wp��}.���q:@ {�$J�dI�-7Wٱ�8�'Nb�nO6�7s���&���l�Ȗ��b�rdY��e�.Rb'A��~pz/;��/ �z����� �9����W��3%�+Hnn1�z!��,�J"�Չx"���>}	G�a(��fQ0�@XA�5�S�jq��҃ό��>vdjJx(}M���ܜ
~�]pݲ��`��F-o m/�i\�f��:h^�nx*�1�e�C�7x���z][�0ӠQc�]7�����R�v�'a��z-��1�T�A$4���'i�	Ѳ��6ձ8�t���q*ڎ�ug�Cys����l�L~v\-�ߺ��ʢ
���!7��g����+b��9>!B�Uq��;8��>�;T��66�4����
u�{���w���C�����F�J,(�G�4c6��w�5k�?�h9;1�'o�u ݝ	����qގ-HE�z��
5 �����,��އq���hh����F�A��D0J/�P�V�?A���j�r�zmO�������g�F�ٲ�{��c��X���xo<���yL�;���9u/���&~��A��JھA��c���z�e��j��J��R.�Pȃի��ߕ����صmvn۬d>�c.SÑ�)�|�8^:|���#]n>Ԫ��H���\�!��F�T��5v{L�)~f��b�]�������cx��>wr�ͫ���?�����%����~��S4ٽ��.Þ� �m �EǶa�(�Ј�Ag����_��o��v�`ƺ	\�w/nz������d�j7Z���#�-��|?~�����t"ڱ�vPYr$F�e���J&�Z���wgpl;�X0�7�%��zٴ�k��3P!�nToPP>OS�lJd�*�Ky�i�3�j�vD#X5؋��AU�'Ξ���3�Uʘ��B���AG�
�NmP�)���/���>��"�3 (�IY�6Qap��iA����A�LE��ʩ�O~�����:��h���F-g	BDU�zM	I?t[�C?{gN���TC5_D�R7	�HS&�pd�`��0��-2yLTf� ����"`��B�9�q�6z֯¾��BW��STj�fL@Ņj$}:���*V~��n�K�6lۊv��/K\���`忣C��5�3q��A�99���M$\����@�܆��w���,	z�Lje��3��=��ҿ2�w$Y��J¯�^��mp��� ֋wE}�D�ARܳ]	���__y�+�s�VT�Wv����wH3!�J�\���%K�Yj��G<�圸���Dp)p'I>��w���W�	C�\�Kq����
������ݼ[�3�_9�~���Dj�/�7V����0kz�ߛ��T��5���XQ�zg�b��������GBPk�K�X	u	�f�J~�6-[��9,8�;����;Z��9���=}M�L�T`���VӘ�Y��@�T�db�+HB��xϪ>��[���"��-r0e��: U|�5�̷�֫"!N�&�4h�(�N�ҕD�B�
��_�������P�����^%�8;�B"١����G3�VP��Z��:�w!o��`H<�� <j|�2��)ty��*igF�?mV��!X�Ph������N��V�%La��\��"n��!|g��g&��?��v�0�`��E(�)�2��+;�,�1	 $��J���AC�V[�A�V�Pzz�B�\D�8ʵ�&��2���)@����NO>����ќ�9�W�B�xN�O&����I�;����O���r����0��������}���җ�� �}�O�{����3�����/�1�u��o�f�-4˸-YV��J�ɩAމ�3���-�5WQ(Vqzb���\�����`:SF��17Wk�C8�D��}d��j �i"�i�VȠU+#�c��Q�{ׅ�x�6��I!�"m���Gq��)=6������ؙ�N�2�2�'�?�z�\PJ'��f�Ĺ�j![.�ή �lIpnӜ�PO�Y�>�Ԛ�d�'�YF�[�Po{/؍�����۷�w���86Y����ŷ���I�gȗ�1a���6�6E9_�A�
�|��R�H�\}�mۂ�x��_��3;���Oܶ��_��2#��?��+����O�x�������7�r޽w-�?d�A���d2W����?�o��C4�1��Q����w]��/��R!��%��5IZr0���`�<��!��'ϡ��@$>���ļ �=d!C<�\f�$�	.c�Ȉ��nA�"�����6(�3��MUD�A�� qg�2���E��yx<54*%�s������n�F��<~���̴���BI�~2���Bv�"%�B��w�w���I
����"    IDATIt!O"�ę��#��cl��2mJ��r	�ad[FUK�9�47T���Ȫ	�h�E,�i1���c'�xf�lA�87n)1�'i��]�r:\,֒�/�
��L��觀�I�j��!��2-%׽�twczvJ$��AW�R�$.�ҹ<��Ym���Z֮����j�w*��j����0��k����X\1Xq��*��	�J�y8oo�sfxo�p)�/��گ�נ/�T!^��k_�<\U���b��̱D�^�����_x:�A#��5@l��.�|��_�A}DE��Ļ�w�7ᷫD��!Pm��/uf�ׂd��,���s���(��2�{}�,��x�qj��\��;��g�y���H�.����I��^�ڴ�_�ߓ������R���������		��U�Z�ad�n�~�Z���+;z�?���r�l6��N�����B~��G\ �J(?�zK]��"3�g���t�����O���'I��Ƌ|-�ZS��]<gR����X@����ٌ��B:��ܜȓ]�$�����Eg��+�1r�X���L�AX�G{�l�+�f��B�N��<f�&�P�B� ��5�C����4f�^\D1�C J�ZL :�{�9�@�ܢ�� 1!0P[�rF�K{�t����b�H�֭�b�KϿ�N�:V|��5�&�$[����!�k(`:�ũZ/� �	r�� K
Z���T�*�%����4��"�,�ݝ��	����H��HX�=����l�F_�b�S���F0G�&P����gǁI ����u	�zo�������P�;r 4��Š!�2��3�\�ʏ�k��d���S�]<���.+ׁ�"jo�<A��,�GN���(#�(᢭[���W12���8�u�w1�0��/���̧�k�J�*�&� �bx� �(fq��YD"1���Q����5�F	�)fpz�,�?���������<*M/�7nC��>�"'�e8�V0�J�:�h�Y) �:B�*J�9�$�سs>���{�ZtG��r�N�A%���O<�7^ۏ|��b��Z˃�� �y70$�/	��xP�V�-Qn�Q�7��V4��z�ZEB�H}!�,B��'�@:�Wǫ�(#�[�h�0�ߍm�7�]W^����80����๗_�Ͼ�����}���C�/��/���<2��y�y�z��� ���ء��?:�{��W���+���}����������o���Sg���n� .8ob�&bl�0��ߐv���|z��\�?�����q4�>����q��c�7O��f���*\(�p�(�*�c�ď|	�FB�h�C@��!�Y�7�gS�1���nx�2A��m���Oh����׊���Z�~o>V��y��i,��^��%�C�F��A?�*[����<�3�L��02|�ή�� �x��Qk�-�7�@(��?G,օ��at�E+�o(���H�n�W�h����B�<7nHt����d'�洕Jă�H�'�M�Q����dB��ݭgƄ`�3/��-��h�=eR�C���['�@ΰ&!X
nY!vf1V���R]b��hPثUT��o�����u���Y�,�����S.y&�j��ʠr)�uxj�q\�O���`�ݟ}}zg���
fx	�j1+���[ɺ�%�qm��|�ex-N��(3(����b-�g�m����%׽�\E��c*Ӂ%<�6S�I���۪�Z�"׵�kc+�.! ���Ҭ'��Z�T��Q���D�ni���V��4�lR��r�<+�U��ߙ���ǲ����0�<^��!���<
7s~�iu�)1`�O�� �V�F�w�k�N��D�����G0�����Z� H&�	��XԘ=;_̼p�� ^��s��C^+���m����I-Ã��ip�vM(R5sS��k�$�J*���I�f��	���K�� �s�^.�����"����(�"	�;ܼ��#���診�l�O��xƣ�'�.qf����W����Mɟ���b:���Uv�\�������:�q�z�^�U���p����oFc*�*/�7L2q(,�b7	vy���(gq��+IpI<��n�����|r��8���/ޑT��{&ć"����3|�/�f]�+U�R�ཻ3��7!=;�g�yF/
hpn��G9#�@4F�ZV"���$�����$��Pz�)8��U}��W�[�v�S�|&��ǜI]*���8t!��Q����(�s��!��GЙLi��;�	�013��^��N�����l!I��&����AK֧���
|��;;�u����A(���c�/�P*V$R���£<X(���IX]�^��1���	*d]���7�=�5�>2 �W�?3���t�pZ*El�W��q���8|�4��ޝ8t�0.��|�S�Ɩ��xk�1<��#"�_w�5�������O�M��}Wc�y;13��$��؝��S��Co������019�3��X̔���h��(��hE:�
DPg"f�°��"�&��ڕ�ߺ��&\�qF��-,�6?�o��Zf�G�P̗04�����'(�҅�d��:8,2�d�T����͢P-#W� S(`!��\6��LN�B�!S�r��l��\�"�"qd�9u��s��
�����p��ׁ�G�$��N��o��_��|�'�SB�Z��&U�
3��ٿٍ�2W�#������,��g/ٶ�/>wӥ���K���g������ppͺukї�#�E*�@2G4��UCW"���A��c.��/���'O!��B��@.W�ڑ�8��]�Ivjc-䲠c#�]8��|��S�q�C���'܏���u~��V�)�F��M��i��Zx����C�Bh�.T������R1�z��Z��z)_%����|!���
�b!��&P+g�!�0�QՁ�W^y	��4��L�%�����#�CzqYV�8���K>�����5��$:�=0����m��0�v��
&�"��͕)�CK&����P�++v��X�!P27e��
*�p�e0�M���/��7_z���ޫV�9���*�
��X���A���LB�T2T�
6��ÊR�K��
�``�(n��&D�b�MσF��G]e�\m�^��v�ו�ʯ��ː�Q@f��qwPSq[V����8/%���d������3�)֌�k�I���,���P0�7s���@����Y4��8930�O���*��� 4�%r���6 Jx<�:�+�"]�hx���DQ
�X��#�x�ҽ]�9�R�"�3�?�C�P2h�[���e�;q��Hu���]'��u��͆���ф��b��`O?�-��u���Y�y`�`a;Kl'9(SR��͍�G�5߶�X��6�v~�޼��
�M������e����C���I�ҐMH<m���9��;s�I�3
i. �j[����μ�R�1�� VKɧMd9^"��(1Au���.e���(���"9I+(`�^K�w�1��7LZō"&���A�#�;�c�9t����i�`>^���T6/�J�V���5I���z�T��j4|~]��':0;5�.1�><b��*��F�C`�_�D�TCde|��4*U�6i6F_{��"޶|m�y�~3�$�l��S�a��N�ԅB�K7�~�u/	%cXI���'W����(�Z�*1�}MNN��-H$"�م��!�T��L��Պ ,�/={M
�@��ȢS�^����P�����Т
��-��?�52dANґ�:Z��: ����p��{�g�Vv'Ѫ���;2dW����D�v��k�rUr�)
z��(�S��������VG��]�v����E11�ų���?��8:D:Ht"_��� ��㔙��j ��VDe|��}�����@*��!�~�~dE��s���p_�g�M���	��P��1cµ��d��=��Bѐ)Z"�#�0����l��Hg��� y��?u�zE��/����}�Jg�ϟ�9�{��Ţ��oæ�k��/������?�
��[���[��?}���w�N�q�m���[oUru��I�b�Y3*��'p��	A����R�3�b��C�&��������x�	�Y���m��9�PEg���m��k�e�0PΠ�Y@{!���$r��"
/��W)^X��xB2�{�L�#��v�����B蘩Ri?*���U�(��(q�PF��Ʊ�q���~8~���D"]��y��_g��5Q(����[�����`����*f�|�����+G�&P��P��W*�MO%��LY�%4�Z�[m��]H_�q�/?��������zu��C�}���>67����v� �ѶT���Z"��VB?�����|�3�Huw!�J��<3�`ڱ-�Ѭs�-+ �?TB������@�cH�Cd�S�2\t�:<M���!?H�����9s��k6��Zt'�ڐ*�4rS(��\ *y�B^$��o+Ȩkf�,�!��d�H�O�^�jE�l�d�b	_�Rֽ�C��F���`�_����DiV%�w�D��#X�q.�{9�mہBӃ�s3Ȗ*hQS�c�*�_p!TM{2�ep�GA�,�me�k��t��N����_�th6�a��~:�&����o%~ߙx�j�H������θ@�U|M{�%"��`������RBp�-7!�����������^�eq-���AȚJ������vMlB������T�J��]7��V#-��7 �=?��*��Xղ�2��T��}3�bgȨo���#�J��l��Ir0<V&]�@d,�t�c����$0�#MG���*oL,t!\��|5�pQ'>�ڬ�lF��FU-{����� VA�#�Ѝ�Au��S �b޶��;� ����J8���~�� ���Z��2��`��u7�ҬgU�9^L���P6n�����~T �P�.�^b������U��2,A�ͭ�lӡ��Ս�<p�flAK���6����I�)s�H3������r��3�3a�oeB��v@��Ѩ���2�% �1(�d`��$��n%LB;�VV|���6	����O�@�! n�td�cI�-�Q�	[S8��h}i-؎�2*�_��sNΔ/W�dy���[35��`�<�X(
Z�f	�X}=��1Д�G�9U���K����:H��G6�E�X��S�呞�E>�E�#)�p�3��U�"�P��/r���VrA\"� ^xoJ/��.�c�g��q�@���8������Ln�߇���I����Z�H��78 &|f�F]I�f	j8^�ȱ���uV)��B>/֬��/^{�eL��1�k��NX$Ԗ�f�HTѮ��،���^\q�&�l�Ƨk�i�z���@`-����9eJ^.�g�yw���YY�O�;j٨��'i]�E�����?�2����8<>�H��`TYo�K�5{1;V���F��������7��2�i�;ͺf�`~nOC�7��B�Y���Jf���"Dl�3���pU���_Yj�^l�ǟ�#�>�#i~����-7}�>�
u;�&���a۶mX�n�{�E��?�?*��Ƨ�w��c�?�o�q��������jt����:!�`!Q�!�0�Ο�?�<<����'x�WQ���O����ƫ�9��QDeq�VW�ކO�|.޹�F	�����<�
:�~���Dc����1/��j�e��m(v�!&�"i�}$�ý����ڰ�ܖt/�+�ް�;�����4�x�U�]�����MT|��J	��s�>}�2�1\��qۭ7`Ϯu�xK����^9x�h
�ҥ
�ݨ�����1Z%߁�̞:jS�nW�����n�������#��ï]���~��3��j�Q�@��T�I�X؃����^�wm�&wZ*1��8��q;\����ԼA��L%�	A"C<F/`�<��|�G����E8�J	A��l��4ʁ����w����J��uL�{������+hיT4Ѭ�[�F97�v��-h�R���"��J��[D">�c�L��[jʕ�Yͬ�5[�S� 2���g9t$ސ�Y��ڑf�{�a9'3�+�Z@�6���v�ً-;� �H��2��%��X��$ܶ�2���!H	X]t�o�1�����E�"T��N�b&��'N��+�#I�:�1���؂�Ky.�2n��&n��Z��KL%��Q�&A����:�o��T33�tc�T���7���/+��L��`=���0��j:-�������d魐���Vvڴ�Q��!/�N�B���3ash�."���	�2�5��d�,J
��ŐNB�C&4Kɞ��aaF
�D�RW�kMs#���IV2�0dp���ҬWѕ�𴦅nA4��Ye�aƉ����)׺�L.���v�,I�-w�J��׳5�!)�����-CԖaΗ�[+�o��(�g ea7K�dU=˷K��@�ڎs�v�%O0r�L�Y�6	2��m
.).���t1�<��t����t�򚨁Oe*cH
�8�R��ΑU&����2o[�3�y[�+\�uEe��f��L:8�Y!6��Ց�\3/�DMV�U�5�-Wp��F��5���i�b�=��HH^<C̼�uj�9E*;&@����,��b7j��M�������kv�:�b F1V�	��z�:�
����#K��٬�WJt!.���bf✤�׎���uk�>�\3�$���P���|=�C���B�X?�ISٰ<\���\wN���>�s��U.�07=���iq����.�����l� �P��H���,�*9Ƅ�r��1�7 ���c������t�?+ۂ���Kч�|��Y=M\y�����n�e�C��:/Y�[�k��f9�5��|H����-�����ߪ� ��� ��)I�۵I��X��WO�������W�������_���;`j�bA����}�6���b$e�\����<�*�
�'�5ǋs_?o!�=����w��ּ
*&��kr=(	["se�z�g[pōOfp���kwܩ��?�">�������R/7��8�5�n�3�?���D�q|��Ob��]x����;��1��cþ}�FwWR0p���v� F�x9i�ZφJ��ߞǽ?|S�|�n��^T5��_�h�sH۸x�z|�kq��;�Աx���Shf3TH�H�B�X0)�U�Z�JE�$�sMG�q��uͽb�B0�h�'J�,����ɇJU�H�D1��1�^,�#�x��i�J#Wc���o-�XT,P.,b׎M��-7��W�E2
<���{��819�L�^xC�u����a��>xCDoTD�Jhff�m^����=�{߾}oo�-��o��W�!��^�����f���e�4X��P+���o����>tûq�17>��o�y;w`͚5p1��ӧ΢Zm"O��d��x4�v�Y-����Ӈ����l-o���	�=�1���:2����=L5�A8�xe��J�ê�D�'hPzn3�c�ΟC�݁v�vٙI�|�%��b>�ba�RA_K� ���KRTGO�D��>��bk�/����l���i�l������ڋ�T�p{�B�<ۭ,�%1zޅص�2$�EV�Y� �/"ޑ����r]lZ}iI���	�������Ot���r.�srܜ<{s��A��JMʖ͛�9`����	BV�
)P��9oڊ�	�����Z����5���Ϣ���#�����!�gq	��C��w\�rh���XrKfpo	�a��Ӽ�$�DUR�nW`�MU��4-{%Fݶ�e�D�Z�vl]�<�B�_6�!K5{]D�8H�Q0נ`_�|��8�����^����B6�AC�s�u��8N��t'\�k K���t/�ī�U2���5�K��)7�v�\;����DR��5(r`�6�C��V+�I7�YZ·�Vf��������籙P���R;P&0\�x��4�A����N+���C[9��)w�T��z�1 5�����    IDAT�ָH����d�u'����b-Ui��ej���r��f&���|�����Ӷ���sLE��n���bCX_n���
�����̾�=�R!�|�~$Ti37�N��`-Ͻ��d��p}��t�h�5�.�8s�-u(�I��l3XRUۨ��9� *@տ�:IX�{�p�x0xf �qd��u����;�1_���s:�]���,��:	�60!i��Q�Ǜ�`��&=�?��%�[�o�1���3�2�R&j�~	r	�k��%����(Q5WĩS���f"�?�
�7n@G*�t6c�&c���֒�bR���3G��Ǒ�19~Zɀq�6��*蒫�"
�^kH��Y/#�8��+���o~�\�szha���T���<���4m`���e��@�L]{�LQM��oQ����}��mE ���-�݁B�{��¿�y7�{m?��$"������_���:%t�|��O�W]��}��غ������"z��Ou��J�	[�w]_��.Z�n����&�v���"�l�UM��U'��������G����u%3_��qۭ�U��z^䌁q>���q�]w!�H�c���܁g�}߸�N�9|����믕QeB��Atv&���i!��h��ٶ���8�{��:>��'��T��� ȳ���6�*�q������4Z���<�����,�QX��3��nkr���NXL��$�ٮW�*dr�۔4��4�;����4�PYT��ĺ�ѳqH����px*�W������<�m��$��]�ɟ97���p�V���[pյ�� ��ٓ815�v8��B�&]�)y�H�>�4Z5ʙP^,^u��/^��?��o<���� �}_��v�z�;����^��,j���
�D#�c�;��p5�ٹ'�<���86oۊ�n��*��~���uشi�	b0���H9Ħ�՞k���(�}ߋH���'���	�&~BnĐ���a�sS�;�!&įS���*����*��8��3'09~��<Ъ!��!4�]�O�XXB��E�VDoO
Ѱ`;̠�\|	�٣��?D�R���H)Q��h�ݡ����ge�a�K������1P,�
��i��.ր`���u�E�y�%Ȕ*���7���#��\mV�e�`�kӴ���R�ȯq���`=�^�b��)���їH��ͣ\,b����8urLwڔY���V�]�@1M�̸�M�X Kҵ�����
z7�ƍ�����ŜƓ�(iH��WXr*�>�r0m�M�7��`86 Y�t�A��p���,��@[�J�pӖ@�Pђ7I�d ��]�z����[	�=(������%I�G�ƃT$TV���%2��Ms�4���{z-�[��\b���V_��;e�e��J��+�%F,��yZ<+��̸2�p���I;v�P�$9�䏁�8&�6c��t
�������8G���-Mpv�l�$�w,)�Sֵ�`�9,���]���=&rp�LŪr!50O����ɱ|f�1�6�$�h;�-� 3@f�j�TPl��1�|^&@1္fC UR�"��7�ҥ��k�r�f�ױ���W�o���8^�Y���j	��R��ƵՌ9����C�y]u���[#T�`*��א�]�ŭ�L�nI����j=߇��*2�`jX���;t���3�)-u
;�/��$OL�L�����_�� �f�2'�g��c���A���b��/T2���vE)Bx8'	%b0� �&�م4�S���� �Xyg�J_YI93�\��ĸnq�"�V*:��;���:7�J=]�K�M��҇�l�Jy��EB_�������V�8~�8Ξ�T�BO�u�ף��W�b����N�M�PdSA7E�#hˠ2½������z��ob�M"����TV��F�|�VQ���ĭ�₍�d�.̹NOL�E��h\�L3��[���-���{��[�d�f::���lAG��qGV��K$B����b/�qO>�"N��F�ƛ��9��hI-��x1�c�{p�%{�q݈����Y� ���in�N�=����O�+�`G��1A��ipn�+,?��6�G��� b�{I���b������q�=��|�w>�+.�Lq�$�QtĢ�N>���p��D�>��ؼy3�x�	�˿|]	���8.�p7�Eͧ��Y�)���,��G�`����	)��O_=4���y ��?��/*�-�_�b!OGz�}{��.�h��gQMg�.�� ��C�vҾu����x�D��Eaw�|�tFIǉj`��>H^6�F��̹ �'�0��<^��J�E�p �nt��El�Z4�]H�|x��$�}�M�9>�s�"��I�}4 � ��Q;�����#زm=h����/�Ǐ�S�22�M/j� |�*������,�B��J>Oq��o��/>�����J��_.����'_}���~��-�?D�,���|N-}�
1�����	�����;p��q<���l���!e�?���;y;w���/ޫ�/�b��i�2S���X{���y�jI�{���iA��K8N _����$_V��˙,�t�:�C��F9����4
����;����y��5�bn��,��W�f�jQ�W_��4:2�v�������_��~�"�Tj^��q)�Y�W��yF�ITT���2��&��T�%�H�j��� j���ـ=�^��[v`&[D��@�ڄ/G0�6��������tu�+�V�M��3�[��J��N 7�FG'g�073k\���F�w.bf.r%���pMA�	�yo�d���0�>���l�x���4�A��Krft��B1��q|9�#��%;���`	+� k)X֢3;�g^c��|�¦jf!Ive��v� ��iC���� ~����5�H��y����n8B�����l3�,KRTG��\%R�����E�b�q�S��A^l5O|�d�׼�U�w$	�΀q 5��. fE�����@M�V�M��i�s��Dݭws��u@:���zNrrt�4q�5���بJ��J��W9�I�����;��C&q2��|�$���V?��?&�Z@K��%�}
n9�L�m�u���,��5�ƕ4M�O�p���#h���@]�&�A�!a`L���J��3�GH�_Lt%�h 5����re��r�YL�8�uг�ʄ�ٲZ�+����2$oY�W�c�^�"�d��o�7抦+�D�A�a+~����{ɀ���Z�Cbp�E����%�9gڭ��E�-�Z��T-�D-�-�%�zf� �q](U:3=-��t]�j�~���dD����>�7�ȡ�UgF?_�������Y�_h�y0���J���N�F��2�Cuu�Q���8��-���g1=7����p����ST�r}DR����+��*�R�Pa��'O`�̸$7�z���~�}J���DF	�<|��2ػ{+>���ʋ�#�B��+��_<�?�3d���]�c���X���7�3�\	g�F�#��ML����H ���OglGGJ�q�K._�B.�*�<_��EL�g�h�JTd@�D�X@ Boo?������ٹ�� Z�<֮Į��4w��[�Ց#���q	���l�ZX�bw�	�(>+)�5e�f`�AT�U��:J�%��z�vh �׎`hU��ګ�~��e|��㟿�m�Z�_��?�����1����2�ڹs'.ۻ�H�<�4z�!͍�ƓO=���###x��އ��^=t�������� fffp��1���P��]���oņkPn ���~�<�Г8>6�)}%x��J��
�}�^����"l��'���P�PFu1�]�g�aanV��J��&�����1�5Р�x:�������URvމ�`�6�L9P��Lg%ǌJ\���=���"ܳ
��UH�ـv2��3s��z�%�Y@��T?�&��J�ʅ9\s�.�Ƨ?�-�m��l��)<��a,�}H���x�:DyS&%�*�^.�k�F�
j���˶}鲿��7~�:~��|�G�S��g`���0ғ��YG1�I��k��������ә����`&�X�v�R%��{�ǩSgq��Waυ{uP��EL"C$�/�d����w?�\-����J��k�
�~�i�����;n�����
XUxZU<ĕ�P��`~�ʙ��'P�͢]��4' x�����Uf#T^i��ҷu�F���|�׭!���ڵ����/���"�F(���E�D`f�VI��_���n�i��Y��F-[�m���n���VP%~� |1�ۄ��}-��^d*u����~DS=��Ƹ�V�]����\|��x"��#��cqa�r�BQ�!蚥�������@A���
T�[  �9�E���
{"���xQMm[��?x#b]���[�k�j�j\*=���4*�8|�r�pڢ*��p��@�q��� �*U�8c=(;Y3K:���
�S�Q j!TQ"t�e�>��Y��j#LHxi�����d�FL���n�%�1�v]S�3w`����dX��;��S++�Rlj����O��E�);n�ȧ��:�q�������������1
b����Ʈ�<���wMS�3I!CF�_*�;�=�Q���$Dz/M:3V��0)�	����ov�̼���4�5�(J�aBOB�W�53F��e%E�OZ�������޴���o8��7^�:>46��R�:�ۦ2�H���=b㍳����{�"����򐴿,�ʤ^�DI+�,�[�e*0�5�X�XFn���|�0�|ZO̳�z���	��r$(�5�9��q��5�:r��b����٩k����h��.$��5�ﳤr�]2��k���pȯj(�K���L��~�s���O��ՙ����s����Z*����@oo��)�T��p~��b'�IL��S��o�5[�\k��Brε�v&��ަ.���{a����@	Yp1����Թ����{��r�q�|Z��7J삁)���#f]��Q��R����^�u�p��~��ҋ�Dp�����׋��8z���h&���"Y,��/^+��g�|��U{�C����o|���}��,w��hĈô[��X}5�K�i,V��c����!MD#���-��U�)t';�����WG���9�:3.߆��U�P��3��Ű�k��YuRXt$8M`frS���7b�M��<���sҥOuu���Cx��7p�ܔ<�z��DE)�\.�䧠�ʞ%�1Q�QY��r�:Ĭs_��k/���u����ޏ�^wS����������@�� ���S�_�/>�<��>L��UW]���������S�q��Dc�޽�d=����o �m�&���3gp��a%�?3�s����'0;7�����~�38o�6�����ϼ�W����YJ,b,����n����lH�4�3��O�!��U��\X���4ʥ�ᇶ���C��DWG(�Q�d��kv6'�Z�P�`��L�ǂ�1��1�-�:�斗>G>��X(ew���x
�~t�[�Ъ~�#1<s�z�����ɳ����	`��)�3c���>n��m(6��^}�?��fJ�T�(����\
uL�bT�O���6Q�?��t�?��y_��#��z�C����W�!��x���z������÷} �F{Ů��I.6:����q.�cH]W>hW��]���Ӹz�u8＝�X�)W�c;�CWi{���p���a�G�sTrج��EI� ����UvV��n�̨k�<��,�R�Gf�,��T��(-N�V���>�*<͊�Y���S�TT���^TC�y�Vlڸ^U$��ذq�|�i��������yD;�$q�/�u��d
�`D�kW��&�D(׆\э۪�a�<6:���]�����=�a�y�ETI�(6�H��B$�R��V�T��L��M�ٔ.��p@����TK%ɷu�b8}�0N=!'�v�h�7�l��`��a̉o�Lpf0�GkTvX54�!I�5J��Ї`��M���� �bfaVs��j�p��.*!`��%��GWS��?�
w�&�w	-S��B�x����-��b��m�s�<)��0�j������-m4��LB@�G�8��JH��R�~��eV��aBm�n<�l���s�t���eN��u��i��y�LP˟�Y���J�I2���!����z��BlTlx�.蕴�%�

�6e��:�	tww
�0unF�:O���@��V��3.�:�g�劬�>�:�ҏg"nȶ�NyI�٪���
���{`����Ӓ��0жr�L��y�?��hҗ�2�$�R֒��ȅUەR feu?��sD�9�
u��<Q��J��$�T=�z<��YUeM��`�
9�>�O�pwXc��%>�D2�	��,ɫڠQ��%\!1s�&�������NV�KV�;v~���&6�Sj:�ـRN2T2g�����ʃRu�ҵ�j��U2�������g��0%�	G�(����3j>�4o�4k43�]E���ӫ�K��P�T���Ic^[��x��<�5țb`])��	g�:��o�ǚ�k�#f:���@��s�%��;�da�]pI�SR����XH�a	�)ؙ�f~��n�4~�Ҫ�6jǳ��Y̩*�jd{��QB@YI�v��w0)
��"��r��0��	���x���T���]�a��*�;�cG��D(@�L�,v)X�$j��.ڵ��qͥ;�!@�%�����q���Ȥ.�WƔժ:[�$�I>l&�{��	��6mڄ���j,�ϡVXDw'��Wc��(��T�e2p��qIx���o �Q��)��@0��e1��_*U�Q-�0v��z�5|�C��ګ/E49J�`IA��������#�}�lٶMEV֙̜�B&��|wɹKh�G)a��m�ڊ_���I�k���}�b�P��O�}��lNyhjf���G�ڷ�����տ�k����'��?�1榦q�7�K�Et���V���A��E�V�U�\!���i^?�wzf�<�({�	$S=��>�իG���?��O=��c��j����i���9�Zq������?�ʘ;vD݁��Bu����E�i�3�H=����)rS��E(ͧQL�ѪVA�'��*{�$Kp�o!E�������&8X��`>�mb�u�E\�y���GD,���ѷm+<}8��a���\o����c�(T<�T�8|�E�������+h�x�W�!8q.�l#�\��"�_�X�8Y���5R��j(�'�n���{w�Zu���������c���W\�/���݆-�0\�٘�ŦQ-\��&�4�v��q ��N��{��Թ9\z����Ke��:��d�����7�����^��2�`k�]�P���rW$��"X�6~WY��"ul�S�� ={
��g�eQ�L����t-�iVU.��$�7�U�;:���f�n��:lߺo��*f�&��1s]��s:�z������ÿ@"�'�P$�\�dZ�0�a|�R�7V��̢`U��!vho^j�տ�?
�t���b��~�^��k6+�],���E ���aݶ��8��L�T�W�oL�
1�ԋ�j` �N��ēx�����d�O$,��0���˶��եo1�u]�[m�#AaQ����2���Xr� ����s�E8�0�s��j�졂Zu��1Ն�P�E�����S`Zւì8,���$=�*C��$z	��l�J���΍9�I�ɑ�M���v	MP{���!X
7�b6�d �l����r�r�*��ꄢ`H�`�bQB5�ë����EB�t�h#�]��4��:􅩧�[k׍����T����,j�*t~��Ãr�4R�jUt�m��ݬ��M��744���6�^x�����b�3��Y� յ�Le*b�?��{��'��|m��%OG��B^�cQB��H�;�*�    IDAT��1=;g�R@cC�N�'J�2�T�'�S�8�kv�,��c�D(@*�!����I%�D�[�!Ke��䰼�WX�+ԡ e���Tu���J����z�s��Ԥ�\�Ŵs�6
�� ¡$;����y 9Knd1ZUS&Ԥ$�uW�S��]1&��Uu���be��Q�,�=��¢QNa��j����J�}����I�ϫₓ��ڪ H�*���Kn:�"�«j>[ε�	�YP$����H(�R� S*v��0IfL/춗]戂u�5�b��w��d��K�?	��p3(pZ&�TJA1�R��.�tE�R�Pt&~^��}t�z�gV5�� Y�➃�s� �noֺh�����DJp �]1�0�Tl�Ȭoǘ��g@�P�4a���23=���oٲE��=3΂��Ĭ�pɟ�/��2��ǋ���C���H<���:;P.�8��B��\B�t��$̋\v��$vnY�?���㚽��A�D(�K����<�ؓ&R�Yo(�̂�6ދ�^���ܸ.��Q�X�z5.�{6�[����O>���	�iui��T�!���̴L�z���7�X"����r�%�htdH{gz!�`~��Y]Knq=])��u�p�9��fҒ��yw��1�g2��ʫq�%#�	%q��aLNLH@��+X��lm6���kC�L��
�܆�DJ� ��峨W�ش���ć�ћ�^R8R�5;���s7�}��X�a����L���{?y��s%��}�����o�+�I.���Ԫn�?�X���,�p~�hB�7c v3yj��,���^����i���?|���Pg �G�E�҂��@w4 #��n�W]��F��)�seDZ~��U�J��<�p$V��#&(rL;�����jTG���1���&l0���0�>ST$얜'#A�������8�KDX�x����8�jU������n��=��MJ$~��?ro�D�Mi����������?������s�A��b��|��
P>v �j��n�KA��
�g��\�������z%��۾����~�gϿ��7���y����&��d(j���D ۷��/�G�VA:���'�씋���?�3����s�X��b-���<��I�u�k�ʒ�1O0j������Ȁ�%�9�P��#J<=I�^�e�s��Ο���	,Μ���G��`�B�2�P�k��R�A[�H2���E{�Ǧ��%pj���E�H7nٌ��!�ݰ}�Cx��G��܏l�s��$��:N�9+Vn�ܜy�<��o�FpblL�O��"�6P)T	���uË�?�Vۏ�t��l�u�nۅ�JS]�v �*!U:�,,A��VR���C��#/rh��GY�dq��0s����$	�b�B|�$�9��r:`�y��+���97.r(�/[ ����O~{�� s�N��R�"���_U�
��E�l3�0������@S�kw��!4VR���%iϺ���N�$� ���U���ʜ$��h�ٜLK
��6%���ؠ���[��b6����X؏D$����(+��(U*�6�|����
�*��]���i8���>��̼<0(=����ֵ��}=qaw����аEY�FGW���KL:�Az!�r��B��R�*;w����2tnL3Bk*<X�v5v��.�ӫ��,c$J���(�
:8Ox0* �T��11�c��ɷ��[����ЮT�C��E�,������ ���qr�,�9B���M卡>7p�j] Eȑr2>��U�a�Ĭ���ݝ"�ML��R/��vp`Ͷ3�i���њT�D��뙖[�&d$&��/[QG�I�Z�'H*Eժ�U��1�oV+�HF��I�Gϖ��<�=���IP07�N��E�²D���++��Qs���th2	c�Q7]
�m|-�!<�:%��h�ZHD��U����I��ڣ챗�"?��e�U��p��~�$�k
sU����Wa�谔�H��»��e�-���C�;/옄�q��[ց���*j)hq�ۺ�=�5�G�o0�`���e�E%h�I�<��r���-�,�e�űfw��Tg���20�&���s�b�����@�(��Q9QşpD������ʰ�$X�4u�Fy��/��܁���AP�	H��>��@�#KsP�Ѻ���`��.$+��Z���R�;r� �:(rf*n���1�.sS�ٰ�ş�P1���Ů�k�'_�,��h�|~�D����w����ѧ�E��X�}B�^y�Ed�V1�>gu�B!�Z�͛7j�P���s<��A=v�Sf^�BH$S*4P�	g�d���mD��� �&},:��fm�C�:11v���\��(	�M
f�#��g+q��=�^MD���p����ȐG뻯�G?����81�R��3�f>��	t$ztمY���X?܅�~�#����Wr�N����,��|�;ߓ��W��㑟�?���t���+���oG<��;�1��$�a��ܓ��T��vr���<yRs��/���*%���x������;zә�e*��b��5��V[�
�p���a�ӏ��1D�E��'ʗ�g���r>Oǂ��b��WJC��	�3y�g��)�@��f��_u#��-x|5|�Z���,'L�ZA���S,��	��CD(�¢T�@:cq4�~���ѱf5:7nBǎݘ-6p�/�GO���/�@���Nc�����?�S9�����Cc(y¨y��7�����m"��Ga�j���@����k�������_����s���O��}�կF:���@jEx���$��kcˆ~�x�ؾe=�="�ٚիq��kQ*��o}�'q�W��/��	��#��BްI}��y`?�Q��=��������omB��7{[�%���ڵ<fϝ���q���d�Ъ�ѮЬ���6s4�l.�̸xDuv%�aݨZ����Vadd[�n����A�a��c�LϤ��K/���lQ�c@S3�:�x0����X��}��>;�*1ߗ�Z�m:;:��w��=*�������v\���}-�� ��Uԩ8I��,�:t�5U.��M%"�bRA �K�wavG�Gaj�%7���2�2 1�e���.�u0��gd�\�����9��C��F� D<����} ��=���ɹ"��?;��tFcvd:gM��w�0�|�:7\����V�}��)S�3� �Ã=X7܅T�A��HPr�M��պ6��+�r������@;���>�ZmUg֮]�M�Q-���Gܚ�u&�HD"�c�rU�Īa�#��q���LLby�.�Nn��T���<�D�Ġ҃U�������Q/Z�r�B�*�Ц�x$��e��U��t&�!���T��z|^BŖ	ܵfMJ_�u���ۉ�k�d��@I�,�[�OgEl\Hg�>G�q3D��Y^@�NV�9/�&�֮����Hă(�2�V��û��mp��4&&�U�����,M~�F�GJ���5�ke���p }���09^\L��kadt5��V�ٳ�16v
�si��\��*/'�\��+Ф�q�@�&���nqK�v��Vfi�G��J#}��ӝ@�`J�,� �����#c�x��֚d8���̀�R+[�X���d��K"N�_*b\{I�/W�(��̽g�\�y.�t��s��f0`� QIQ�L�"eYT��lKZY��ڵ�U�]׭����]_�V����"� �"�$r � �L��=�s���}ޯ�]���u�0�����{��IV.� Zt�!�/����m�0�߇d<���%qo�� Gf$s%�5�!�9��sU	��`�h��/]D5ή�K�,�w ���B�	�t��
.���p8&��
ϝ�A�&Y$)�u74;�Zڳ�z*�'���$�B�T�U������J&���w��!�Ic��s���kU�4��p\��EATl��}54Ԓ~��(D$_�5dc7KC��Dr
��^eq��Vm� �����M���m��׎��ݡ��u�Fץq��4y���p�D����-��������N�b�͇\�ҁ�MdMKQd�B:����R������y���yRBd]43��QM�2j�h�L�K�v�n�W>�Gؿk*��2R������o��7Ԍ�-[�������\D�(b�~yyY
���hmk�s�� +�I��pv�m��hnk�u��ōX��)�0s��hW��9�K�*/H(����~ШȠ�3�s)�Z�5���P_�3o�@CH�[~N��������%9Ft���@t��d��J�-z�;\H��.�#M�l� �@:FO������ć6�J�e�[^Y���+��g?GߦA|��_q����ӟ��/_FOOFGF��"G��!24�����!9�`���uhQ��x==p�;�GF_o?X",�%���W��ˇ���A��NX�������ܷ��-H��a�d`�d蓋r&�X"xt�Pd��������byjH�Q�d��03�{�܋bW]��Ӆ�n��� w�MP�l�j�D���V��d$�Ǆ�h��kZ��5`�;�����k���k'1.��sG�������f*[4!�� E�Mkh����Κ����[$Փ���х�;w}�s���ߩ������_����g��������i�f�Sď&��:�ݵ���^�w�������~���w�S����$~��"MattFG�˂U�TпX�T�Yp��,~��5�'u�� *&]�#d�G�!k���G�fE�����*<N;����E�M^Cb}Fn���|0�bAZ.f%g�v.�pJ+�:8�*�MmF���𹐈Ep`�<����*_���d�+R�8t7^�4^}�(���$��O왬�N���L����_��y�P��"��b��H��C��v��y����}��ܴ��TN��Mf]&��w�6��ʄ`�E%�r��
�ܺC��K�K�y�<̹,L���?�k\��hK�Ŝ����NC ԏz�S��u�_Ra��E�BJ9����k��<��|�c�l�#����F,	��i���#*����)�\��k�U�:��ZCP�����R����*R`QOUk��}�h
:`5U�r�t�/K��F��*"_&��
�ׅtXX�brvs+a�x;�����,�`)�:]3����H ��TL���*�(05��+WǱN���E�Y��2E'��r��n̈́��.l���ce��l�ܼ�"}�Ȇ��L&u[�̩rNb�p&2E\�1�p�3�j�T,�$����@_o|n;�.+l��5�=!��R
�SX^Y���"l��b?g�;A`����"��.�N���ׁ��f�4Y�P���s��l�t��lX�Hcni�k��'��X_QDbJ��!�#�Ci��s����q:��s*�	���;<.y�t���X,#��E$3IA1ı��Z!������./JU6�7������h4f)��N�\W�\;F��u����I�i6]E\h]�L��e�������k��p����w;�U�ky�\$�O�l�"�em-�L�M}4i�����l.���¶���6�c�L�B�$����r8�l��\��dI� �[��x�:��D�A-��L��NWR��݆m�G�ب!�_���KcB��:�K��,���01yK(՚�0]gQ��eF9/�P����f^�e���&�Z������q�8� b�����(���r%�Kf�p��3R<���s765I�µ�Be������3��z�!�8��-*��:=�_�kNtwL�Q	�k��5� _��ªU)Z� ���3|�l��0]�5�-Sj���h�˿_�&�!P�*�&�L#��9_���/cq�PkC� ��]"�|=
E� [PT<3ѩB
�T��Ɨ?�	��5���gAR�����������݉w��طg�����B�H�����	�(��x�'&o�
�uyϤ}੧�mtb�8.^������`�犡V���2���
AJJ#C�<�C.��p��D��5f�r]�@@ht�2�	R�L29�,�ɍc8�m����yvzN��x��r,h�I��q��9]�N�Ϗ;����8�V���3�r�z��=��>���5�(����~����_�����~��-�F8y�8�]�&���V�K��$-��tʱ��:����+Q����4��y�&�V����x�G��ׅ\�6v/���{�5��1%[��5;:�n<z`���#�G>��Rf�DT�v��@��]��')ƚ:ݨ�눐��JC+QL%`���$���m�@�Wj��u��HA�*$u�%⏢���d-�۫��
��-ҊH%ͺZA�fC��V�7#���7����qu1��A�R���	f�j�t�h
��4vR-IC�K`�U�7��k�w����F������Ums��_<t��ߘ]~���G�����UD�7�xػs�{����p��	���!���~��H�3x��aww�`����j�Fm`�C�-N\Z�O_���u�4��-E�t�r�Ň²�n�n�X�M�_���e�(��82�%hU�?(��Ş���9���v�Ae�_
�m[�����n��s��1:,!,"c��2xE���k�y�K+R���!������0{kJ���lA
���u�9{KK��L�ŋ?�vz�'Dw�)�A^�F�*;�B�@��6<���زc���"(W���D*�d:]�6-p{=*�����j�`azs�7�d(�0�U�5FQ*!�Q��]��'+�ޱn��I�$:�bLꫢPʠ��N���_�,|MA�l�����A6Oh�<_�D�b3.شw��5_���5(�uשh�ת���dUZ�Z P�ǜ�_m�V��Vty���$����S���i=��=#F�$r%��n����:Ƨ�qk~U`F
"}^7��[�:�T�W�D~�M���$�,X0,:" �.anv/�!�(��IQC�I��*!y�j�.���ϋ��F465���#�M���%Q�C@�䄓���N�+:A���;�)���q�/E����; HW&�hGmM�����"6x��9���,���ǡ�Wo��ʵG�(U5�+�X�B����J�A,6]�h ॰��n�ϫ?����x�h��٥5,�EK��>d�öM�(f�*!��2%��o�uu �w��q
���Te(W���5@����łJ��5L�ܢQʊ;����G8�ĩ�13�����	�E��k�ڢ�&i�ⴛ��s`�mho�I�`����c���ِ���(U��hrz�K�hl���n�f�.q�1�Y��0 ���Ui�6�LL��9�� ��{�M�L�����48-%�����nR�r%�El$2X^	cyuUh��m-�hnF{[ҩ(ʥ�V��VKR�1f1��G��%ss��2��� �6|7:�;��9pkfW��#��U�]PR�x���8�&i�|^�^�8�,ܺ���F�2d� �@���I�K�Dc9Ѿ��V�(�uhDM��'�h�f��S���]]VU(E|,����\]]�-�����$'R����[祖Se�Y�ܭ�k2�b�:�^�fq�g�A�"O~�_[Y\�b��M�6������A�
�`+��C�W��T4���f�m6�,LO� �秷�S~orr�*�I��� �3hi�M"]Ɓ�������n��,�b`n~���gq��ҩ<�����>�Q�ܱ����� A"��bA��լHB�uko���_8'HB{[���?Ǟ�� W*���'����旖eO%݋���\V&�%���[aC��㤄�E)��9���ڋtFB޸��1��e����|�8]v��,���Ӹv������� ������~��G���)P��XR�s���q|��C,Y�����O����x����ӏ�J��|�!��/��['����c�|Th�<�|����\�#���G���|�b㣄���̒�F��h4�\�x@���ۏ��V�%=z��o�T��a��Ό�RmN��S�    IDATp`t�n��a�V琎�I(%��B�l���ٗ�xq����a5�A�(�b�+D�ё�����:�<�;��b�j��I��VA�����jF*��T��[�3�X�¢I^l�Z���Z��0�1g#~u�*�?�6�e8�:�� 9͊*�ܬLV	B;뚅��ɢ52.���i-&#�w� 1@ο��'?p�7?�g�����.C�W���ݏ>�������	56����8�g����/��9���`;�x�!t6�q��e�&}����߃�,ί��������%��`����f�8�׀�c	|�'gq}.���Rjz����SX��O��%����8et"^��3o`��E���0�J6Ji/�#��ڬ���l��|*�]_*�7���~[�$���^l^�GĠ�$�f;���5+&�o���M�OL
��C�����4�XD*��Qd@�K+��r�*W�~��l 6K�k����)���rE��V���odĊt�����C�l��U�R����R6���Ħ��p���ag��"�:�b�I������@�!�Q��\��X)�&�J�!�c-�8��D�k�Y�s�Ć����ub�B�@��W���-��V�U��f�py����w�e4dR�E��)�A�(7�Z��b�QNN�X�ӷ:'Wg8�%�M���2�6C%@��Kh�Y�us:��w�����Y�s�)Q6D�߆BU���"t��2�9=�+7&N�����Zk3W��@o{36�7J��W7��3��$�!E;AҢ���6������ylD�H�J�X�"�+?��TN;
����GK�*ނ^��A9E[Y]��{(�$�cޣ��inl'"����L)(������I���<�'��ʖ��6�T�z�,���55H�N�EK�	;-��+��Ԡ8��G���'�q��%,.��������f��alD9����pІ�ǎ�� �[p�+ph%x�:<䱓���"�6������9DY�(�� ����>5�K�:,pZ5i�N�m��c�Ù��3OC�!R=T�u1[�57&RR�YZ�~0�
���߬��co��ۗo�l��y����2:�cK*���
���
vl݌�-�B�`���9�orj�c�KowXa�PC �EJ���ǟ�^Z+r�&#�p����u��ee�Ir��h&���I�;�
�.7z����
����j��1��O�4R��sBis�XX.��Ĕ8ٰ���E{s�>3�$���]eh �.�,l � **T��X�t^�_R���m�����X�D��"Kcf1��5��X��*��7bSo+l�
6|.�|Nq%�,/�e��*y�TB4[@�PBQ����vc��IA��=�ZIZ��zD��'݂�Z�r��:��6� ����'Տ��@)y�O��o��p� ��i��YHmq5��]Ì:eH�ȚK��8����y��_��֖We���P���)��*�Z���o���J
3)�)������ݎ�g�`qv�MV�:���NL����X�>�X@5�Bvc�߅/��a��-R��-f�FV���~ׯ���-a����G� C[zn�;B�=�J����>'��0���d~��y8\n|�����HAx��9|���%7����b��E��`4ABU3H��7�M��pe^R�H�85@a3Ž��)������֓�n���L�:u
�ؽ{������C�&�zx������f��7��������Y+%���Gw#>���ç�+E+�F,.����5�_��w=�(�����%������k_Gs�T�z�Gr���IZ�ִv.��9�417oL���e��A�n��ߍ��s��~�7�����m��3����;�����S6�|l�dDr*Xs@B*��j������:�L��%�qI+.�(�H�-	
Zo�����f����	❤�za,~�Y�/Y)�0Lf
�a�1�Ps��G�+�ք�Q�H�t�z�Ѹ� f�v���%�~ueW�\y��@҂h^@ڠF�؆	�!�)Ww.�v��M߷��/��ǿ�ށ.L���jCP�V���_�ѯ��?�-�yx |��ؽm ��v���w�򮵥�:�{�����5>.�������x��ް����B����V	�
^w���ۀ�72�������$to��F�0�g��YmR��6R���o ��l�X�õs�����B�[JJ;P��7�I�;�2de�%�"�%}AQX@���Ǉ�|?>����S1��1�-�p:��K�e���!���xSK"�C|����SBUU�~�%$�9�I����5'������:u�/\��僦{O(䪀#������F��G��LN�iU�e�E^w�aw9�&�'�����Ɍ�,�-"��"���Ysb,�Pm��M���ŧ���$��
s�G_��i
7�*<P��*^�ɳ�i��`�=�{�|����ani^uN,I��] 29N��Y�"H''�=:)�h�X��u'?�~���+�Z�M�ӕ�������9��� ���1�Ӊf�6���S���Q�M�B46�ZJ��	\��)t*��'�3���8�c���2p�x,�bٙʗd�0s�l���^��7�U;|�f8t�Xyr��܃"h��.47z��K}��6�@��ۂ�~-ȥK�D����1@cS>��f���a�+�v���	�Ss�z})X�~:�K�	�k�.��g��M�2 ��"�̋K�ةga$y��n�B4��������m��z�f	�ǩ	Q���ƀ���ft��ఔ��m�%�T�1�ű�a���W/�����N������j!�q�D���R\t�H*9��
؈ƐHa�t�%A��:v:�Bw�2LV3Lv)����Y��t��6��~�i!�ϥ٨�?��`O'6�ke�v`ۖ>�mBn'I��-�J#�P^It�r�D��D��&eڹu� ZZ�V��*"@7��xO�_K��L�:p��U�<s�}��-ފ�Z1��8�6���W+�Z*���h��pe즈����&�9�GW�nU:�5>bkȂ��rR㤼�u���|	��-~�&�1��nf�H�gb�2.]�� �h6Q�n����n�1��@K�.M$J(��h��i�Ն2��U �7�64	:q�2W���U��U���0׭�F+�2%�"����&�������=�9��~��<��/���|Φ��_r	ja�B�ʬ�TO"����.v�^G��ʽKi��+�I��Ƭ�L*{�!���r�ҰH@��QhʪZ3KC^]Ew�BΝ8�%fq��L"�����7dz�h�5'*r�9���!Ż�ߏ?��Ǳg�4�l��kx��g1qu^��� ������%ҠB�h�(/�oJ�&�oU�Kr���>5uK��V������������^x�~�U����~@h�Z���8N�>K5��i�*֬���sq{҄v�	?���"Q�+_����Ōp$��'N�P�'��7l��\LI b-��>�֨~��P�<u��&���LD�)S�����<�?x�aqv$��<���<��_���O
}���?ڻ�P��J�4�BSs��]�8X�],�6A��:�)s�8���\���\8��%�@A&�+�x�
����c��4������l���VX2I���QI�`6
�z��iQ����`s:�`��*Ӽ�a$�ð��I�[,�]�����c��pf"̄Z�3C9Rcx�ȽSӬ���H�j�yIa^6P.����v�j׋K�Y�ح��XsZ�Ь(5��y�A8w��~t�,�.D�59�#���@�C �5<����V�CZEH��D�����4��WR����3��۟|�W�}����Ԇ���/�����G���lx����A%���~�^~�e8t/�/�Z�����C8r����:>���8x`/�\�N\��"�!���S�T��B��w#m.�g��9�k�x����³1���S��PM6=6�ukZ%;�X]����U��+(&�Q�FᲒs�D��P�X*ʐ���<�Z�`�gϛ�X�b#����>����W�����L:)�}^��d�SS��$3)8��<p�����i׮8p��hm��S=ͮ6^��/��I"$�N.�=xz�z��7����_A<C/p;L� �+���ك��$��pZC��*�U�.Z���!�06q�ষ:��TxH��BF�x���f�wGT��*�Hl}TP���G˯��������e�wy&��	C���~�#�zt�/͋�!���dZ���l��8�:�jx�(?��QRة	�F�*1�|�W\křp	%��LB�k��,E��#�����$�N�����-:$�,��qk�����&�ځlM�:���v�ʉ��$���d��2-H�N5~��7�ڱ3�Z��І�� l˱�*����5:����2�S��Ť�㚬X��b-���r��8������Z�s������3������2�:�X�[ZC"U�f�"�50��.<tIc6JH���wZ��{����A�.6���j�N���"���5Z��{�6����ŉ�0qkmD=��b�(�a1���Ղ�C�z̰kU8��5�
%�aa���z2��/t!�k�Q�b�2	��vw`���|��U1�7w.�]��a���.^C*Y���|�C�6����%�ښŐA �T�Aa:V"I��t]tF�	��UF�eY��\XD4�⾔���f���v�b��W�O/u�r�8��<n��#�t�9�� �/N��g�J�m�0v��u��o-��_�p�W�;"	�.N���q0^���DcK��~{��zBpZIǣ�M-��jC���d�`9�����!(�ȶa�t�%䂩��('�<��D��Ŗ	[�"� �d��������:��)E>��6'�-����j�F��S�cz.M�8��[�`��[�W��B�G�F䋳r�YP�¸JՒ	E��biÂ��(~��Y��SB�"�kG<��|*#bP
L����(��I-E�����۩��uu-�Lj�=;*A��+���=�S}@��U4(5dS�bc����\���x��P��*I����,LcqAHR�z�z�	�';CBk��|"���z[��[p��c��uK���LP6�|=��m��hҩ�F�4h&n�%��C���<�];7IA�.������K�t�������A�B�Z�4��E���@,�y~"����-C�XX����cضm��G,��4Ν����G�C�9	G֑���]��	����Fd�D]H<��<Ɋ0kJ;R�J�@'����k�b���?�m���[�Ù3g���Ol
��ء����v����#��SqU�Ĳ8ya����+�,�&���F	�!;>�����O�K�*N�٠q�|��W���/�#MO��:d����4Ї��n9_#�ƨ �kvuU�33��(4���=�]�����	��}ۆTPX�Yh�b��;՜�[ǳ��>ν�&lv���ž�>��,H�,���V�kt�TP6���n�ƒf*��i�	�s�*��Pցp8)�|��a73�E!�l���Ux��gn757J�������P�Lc>�uQ��>4ː��.5DꙥSfl�������u�_:��z%"ž �N/r�	E6��!����ƺLC�(�L����ZՊtx9}�涿����懶ne��~��7��w~��ߜ<��7?������	�L������,*U�>54|���Ͻ�
~�ӟ��o ����:`�h4��@��7/�"�Uq�c��5Ͽ6�g��� \�M�h.��j"�5�h&����a�
�-pj%d�k���6�o��XF9�]RV9�O��$�A1������	�*	���#������~��x�?$ԆHtU�+�+�qMn*6�WEN8t�8Y����ohp3z{����!�iR@k������z�*�S7.�[��	Wo��V�Z�}�:�����a�f`@��a���ix
p"��d�#�ֆ��Y2�"�1�Nʤ��� Cv�kX��U���PbB1�j�ڒ���f�`61E��,�n�=ʵn�BBm���\�$�L�;�	��)�RA��m��?oȇ��yq��R�S+6C�r�aW]#@!h�iD�_5� 7���nt�..�=}�q��O^nE,B�VS���ؿ}��,ԯ��ۓ�"g��M.���[H��Ȗ����p8N��Jk��b�rqA.��)�:�V��,�;t�n̈^���Ic�t�(22�:؅ݣhkp���d�zd��tyE$9����sW��G��T8'.W��da��ڀ᭛��݌��������#Ҵ���E��=��D�3��^^���F��A*��=�?Z�����l��ldo/!����Yi�x\�̸:���Gޒ:l��35�bM[N����x��uª���T+lv/`�`n)�߾y�q�y�^U���%�h
�9�Ek�)FM>�iQH���n٤!g�JX�D165�����:����o˩M0�AO_+��[����xE���1�f\��Ǎ�Y��6�J�����^�,ત��T�V6��REw;�`��~�����Keu��"�H��qz����vwv`S_v�lŦM~Anx��I����n�3V�~��L̮�br���fq��M�K���c��SvSE��4��UD2e\�1���q��d�1�C��#�M�m��M+éSԭ()�Ë|�
��s�x|k6�T�T�8��ͧ�-$H)'q<WԜD�9�u�2��X��� �it�}Vtu�0�݄�'�L�� ��� ������WQ�Hϳ�����uN�+j�t�K	.���L'�X_[����իrX\0Q�dxI�-��]R\��iy�u����x�����S�kw���<���sJ�P[�����ӄ��2���dH�eKڐ8�V�acCD�j�(��",#�D��s����籶�,A�Z�7�X:���`/�
#�Sʦ��XŽ;����ǱwǠ���*Kf����-�9�p�o���U����+�`=+��cJw�{8�}�"v�L&��E��}����j�#W����S����+��^J��͉q�U�}7Cػw�8��!�Â��<��ዛ7o�fu=��%�hmi���{�3��$���-���+�XZZ��褱��`":�]%�K�
Ai��aF<c������K��P�#G�U6/aoA��~�>|�=�JK`nՙb�}�M�p���/�ɤf�1�~at���۔�B�YDFI�(�^Y���1�=+�����:"�7���Q�un
�2���,�<z'^}-&�1�C�!��ad�W�%�4�R9��0�*�v�;G���q:p.��$���5��wa�.�-�&����_�Bf.�y�(>�0Ѳ���h/>q��3(�ƺP}!��94�N� ��N�l
�J�Jۜ�x�(��з���^��N㯿�,T-��	���b�!3�_��܂�*���(3��(
�;�XK<�}�k{��?���T0/Կ|��ϼ��[�}�=�>����o��B��X�N/�P�2t�˹"�]����Y,���hᔵ��x��{�}����]g �ZLy�����~�L��]�~~I# �o&��t�H�ݟJ���&b���"M(��[{�$���d7�r�%�t��bwH�oHRi�'��ȌT6#c0��N�߳S�z�7�7�ӟ�#Y�J���]����!�"�y����Y� ��c�֌؋�#G$�X�.���ŀ_\h�,�8x��-�M���*����������~�#o���� C�d�c`h'��� ��V\�YD�bÖ�[~�sO2�P|Hzh�('#���$��Y���X�Y��U mHd�=Ey�+ꄺiH��� =���&`*#BM0��N��VT�"�
���HC�kJCMf����*�>I>e�B-m��3����ԂZۄ�ɪ�2�ޔ�P8���-�72i ��6S	[�[q`�ft6�`)P��.�M�f;9`baק���!���I�
��a�]    IDAT��T��V�asW�ݹ=�~8,��P�U��F��D����~�"�x�,���ymZM�X4\�>ԃ��F�\R��U}���M"m�쥛8r��oV75��"7�\�B�T���GGk=]����PpL_q�G01$�c6\����I����e/s�X��`GH��}�pjE���8��3�C�	���Åp2�sWn���+(t�hE�i��k$E<�Ex�:6�����d�Y���'��O����o����f�.���h�J[6�`��t6pZ`3�-̡��!��	��7�p��,G�0����f�o{ؗJ�)L���D__+�6w"�g�H�y�{ND�E�q�*�ߜ����铜	>���c&�1�$��"��PF�������F�v�;E�+�sGa�I�I�pkn��]����\�>�vwb��0Z�9���!}��	���=�T�6��.(nD%#���-�س}P]���S ^4�-�qe|�/�@4U�ߓi15`�:�B�æ�f�6���V��t	t:�'���.�ss+z���Me�](�����\�J�M-3�]��� �` �C,E+�,R�vܿg+�t ��D�*|$"4\�9���X�,�޹��M����̴��2i�!@B��&�������'N3�lFʐU�b�̉��T�=��s��u��kR�	�7	����,����瓺�s]? �TC!u�H6)C,`i��d_��`��4���[���n�����
�(�n�43�Ks�����t��aҋ��:hl$"��uu	b�]�#�4���>��Ǳ�ͽ��XY������k�%w4����(�|w ��p�Z_GE2��B���l�166&nDx��ڜ��Zd�9����oavv{���'?�ii:�9��G� �}��8~���d��G�8{�,�9"ַO?�����u��-�G_��/S6R##[�/}	{v�������`�B,vAPD[�3]�z<�!g���M���e���I�ꕣ0Ln��S*�F��ؿ�w�v	x�s�5�;��;�C�yU��M��ep��G�Z�&�T��ƺ���0�iBt��@j�8í�#�IciyS�3X]\��
t����^�$�@ �P���l��/��/ ���[o_A��@�MGvi�D��*��)8,(�6W�eh3�Hm��eC {��J*+��DT�$D �t�b6��*A���X�d��At�Tr
���h�L���ᦲQ'�tPi\�w����b�� CB���C��� E�a�`��%��kJ��D�i����������G�.�ח�a"��a���o�j�j��P��z�x�m����
Y�8lK����������;���^y�Ͻ�#��i}�����@UDO8�������Jt	�?=�=LN�I���WՄw�����B1��,v[<Q�[%�8m���o.�'ϟA�������r�!੪7V���@�*,�$�Ƥ!H,N���
E|�:�EĂ�BH]��5	�X,�JC��7�Ê�e����;�=��l�y�U�-�����Qn�L6[����ĲkeiY<99�{Gww��&����^:O��)����.'>����F��������?�`�Q�Q5���ҋ�{D[�0�֢H����`T��	*I�������"b9�UG6����,6QN��Dڕ��}���7k�I�4+3C2����Ȇ@6!aQ���0/|ޥq31�&>���	�{G�?����L��#S��gY�&vѴ�#�Qi ���
����!���OP����:�~Gl��'�v��Uib��T���ׂ�;�r+��T3IfXuˑ������e���,��(�ch��,g1�݄������Z��.if̯$p��$N_��7B��/ݜ��bd��Ў�z��H����X\M���k8ui��_�LXY��Mr)A�3�~6��a�� B�TT�A���͋\фT8v��\�@��{T���!Hn���cþ��ؿ}nk	f#���%b9���AD��
�l��z'߾*(����ۈ�A'$L�&�g�V��lK��U�e_iG�lťks8}aL�74Zh9k���Fk���?�[�t� �A�P�*��`�9���i�tE���v8m>h�B�؅3K��x"����`P������%ߟ��B8a�ͳqkv��$,E<�q��C�/��䓲�*���2�m7a��#[���Hqj���,Xل�-��(���1�=��4]�&C��ؾ} ��_���
"fs�l����I���S��i�ɰ�
\��:��D�ژ�C��};EoU-ӫ��V�:�����g� _քf��xUs�I	:�Fb�H���{l2�+�2>'֥�d�\��زeɍ���D�.�E�[����	��\�9����X<�$�+0U3�=҇w�݆޶�&�n�))�9�+TNqi|�/�#B�*��/$Ǘ�"6p\ɹ�^U��V��*v�|�B��ͽ������R/��ڑ�'�u���̀4Luה'X��6��hV�������8eV����I����&�m��;��@B��ѱr(�@:ZB��	�Y� ��:t�&ǁ7�$�|�&��Ne���"�)>�N�	��[hphx���}�~�B�
����̹sغy#[E�����ZO&���A�b�(��:��ɤ�D2���E�vب|�������-�-�СC"^���z��/_����Ͽ����K���O}�����mH!Oz��=��^ý��+T$~0����C��(��<v�w������p`�>����,aiaQ��Ĥ�FG�j�Rr­���c�'&�L���D8|�"~���Z�(Rɸ���z����x���R��,��h/�r'N�D{{��Al߶��ZH�L�����+/��+b&1�u��މ��.�|�80���\�(��ff�<?�D8,�y6S��5����l�"��N��yud�x�b7n��ϣ��L�W�r�p����@�sq����Nd7��X#��*�9[D9EK�b�"�,C"~��1���B�j����=�t5݂��F���+{(k�P���Z���Er[�Z�^g�V䰎�*
�H��GQN�H�1�V6�;^٪#F�]g#\���e�Ø1l����א��Prd:H��4p4�͢���U%��(g���&���������o?��C���|��S���W������ں[w�܎���V�+�.�"�&�_�W3.ܸ��(�M���x��*��;:�v���n��+��� @��q�ˇdՄ�^�/_~�f['4�/�q	���yr����f� �2A�
H�Mcy�f�/#�>0w���k�4�Z��+�N&u�7K����2����ۆ���"Vzss��YܽwC�9>.�Ȏ�jqJ%���♓�NkO�|�af���Id��W.����*���$� �{{��jD'#��Qc�,I�V8�>���x�����ah>�B�:��bp���E$�E�q��Қ��4-��������s���H`zl�E%�Sr��8u�Ee�l�9�.�S�$.\8�a�ؔ�J�'�eH����U�ze�?������������'f��F�H�������zC@�`�!P�r�7 bz�����SmڂJ�8���L	�IY��<k5���f��Ak�	�]q��U���qƁ��"��uc��Q��ՃB����#ڠD�vs�;!h�Q �O[�n���"N�����e�,*E������h����t��	g��i6?E:�)
�ba%�k7�pki��]�,6�意��9�Lw���ɋ{vmFw�F.�Y�>X��r±"�^���c���F�@��T� ��c.c�`7��=
�����߭����Y�������q-�����6>�B�b�h,=���f�¯��j���1`C�G�/Is�����.�M���fA�\��e�H��	ފ�6l�*\6M<�I�sy��Z�k�Q�v�,��@�:�����6C/^e��G!Eow�nߊ��6iN� 3P���+�Y
�l�
B��Mx��AP��P�W~M�qR�.D�8�M�VŦ�fܻwTِ�+��� 1���0�&�'�t�O��AI ��@��-C����ǜ�����Ya�=(�-�X�o�<�\�.�G3a��f�aTs�x�`�A$c��u��@%3��p��k0@6;|^/��ҋt9��}��6���� �0���x��+8uaL�S���3\.7Z[PHe}Ld�(W
��jǁ�{���*V��Dc7�q�Ҹ؏����f���)�hp���waǖ^UT��Z���X�&������^����O�	&���F��Ų#�H��9%��p�Ά��hXf�e��Ÿ#���u���~���������X-��6�o�"(�*��մ
��c�sU%�������� /�|��2�b�*T��2O"�t�
,:���0rYh�B��=.�N�:>�m�z�d�\���!KAj*)ÜL6/\{� ��G�����'��][�� V��Ϝ�񓧱{�N�O�%{���C��������%`n~^����ߝ[\M�Sx{v푠���*^=�~����^��҄O��"�}�7���](*�'_�{y/���]���{���p��a)�yNZZZ��3�H�ꍛc�ɏ�����@�ğ�����\lɗ�ŝ�C����^�|Hvy��pe�Ia1�u�c%U�/��sGN��n4���4�~~������dkkzyϽ��_|����#=���EK63�X�f�����_;�x2�` ��"z��4(Z���.�+�lf16a�a,�*s �*՜)�C��P��-hkhA��D5�-��¹K�?�64�1e3p2�/����5���m�1e�E>G2�!�&ASY�2J�F���\����&����MS�T��5 S-��󠥳]���I��ӝ�3��"m8�����F������K�_��h+O&Y3���ќ"��6�� ��Mh��\#������C�c.�C�f|��#���Ͱ�^����z+�(�'"��#}��<�s����������[y�����P-gd�a1IN`WV����u/Vc	l$�By��r�����ڌ��Vl��@�Gx� ��<:MM�.D���ǯ��×-x`�Z`��n7u"E�\��p8Lh�2:���4s��0�@1��6�)�����+n�lv�ȝ�E}.�,悒J���P?z���Z��;/0#�ޞ�nI���?�p��1
)ٵ��b���Q��oD��������v�g'Z�1>~���hnlAg�KP&�����ݺK|����boC4Y~�"���3���M�ҹ�	u`������/�W$�C"[^9E��Q�]�Զ��	���#��:���"�ڀY6��N_,�*
ʍ�*n�/�(P|�ȁB1��QB^�ǩ�g�J�A
�Y曤!�ǘݻ��?�1�MN���)��(��@ؿ�-�C�������Vx񦾫ؿ3ySڎ�F}��,4 ѕ �ii8�e�ta� ��:\�?
��C���p����c�Hӝ���@:�,�D�~��x�v��Bw�_�	�)S'@��d����8{�nN����%lx�{FH�q��g6�%>�t�0'|j3+XK�!�&)�:�&sfW�nF���l��;7���MTH�To�@��N����_����h�0��
i�����Q��8��8ԐZ@��4ҙ�����d����(�ܘ��F.o�Ь≬y��P�z;[��ф�&7B~�Ej_�(V$R._����*L](L����;z�w�_lFy�r��c�N��X�څ��+�̕�876�X�+��ph� �A�B��f�qD7��Æc��<���*XZ�ҍI�-GP2�k��$�3]��ǸY9��T�4LP.�n�(�����[�r�JȺ�&T��Ao�ML^}�$�\��!�|o;08�*Bۀ���DFYZ�z-�.���061�������Q��yp��z��e
�"�4��|��Wq��5�"���ɱ�Ԅo[���^�����̈́â�KJ,a`f1����t�r�Q�`�Iʳ��ߌR5�|)����7�2�@-p��,ο}�\Y�W
�=l*E������v��]Є�S��jE&���Z4����qL.D��Z�\`�]�Ю��2��u��u7Q�KZ)����,��07/�_���wB��k��:�>�]m�����j�=�?Y�׬!�+���k�sR�b���"�BQR_h�-�i��fhMM�4H��Ƃ�(��k?�̭[2�ټe�;�TC�@8��D2)	�d�`���k0e6���_������B���ͷN�C�%,�]>���NY���F����c�H�0O� KKXXZT��\��By���'���m[}]X�ǡC��g?��؀S��/��q��|����l*�/|�x��GI�x�"�z�)l�:�cǎ�'?�	旄����~����������}\�zEb<�_����SO
�oea3���K�h	�j����2}Pī������P�F
������//�����i���!ې��j�����+��|�*���Q�^���Çq��u<���xp�A����hV��Jd�t'�>��gO��VW[;��~��n��0��bA����^���Z.#�-�4���0Hŧ�B�z�
�V],���
bӷ�~�&2��@4�B,*5���,��̡��	���SG1�B1�����gOf��RJN�"u��6�-(q�v鰺ݪ�-�%�(�ϣ������`��*�;���T�΁^� �~&�Bv���-�%��	ape�1�8AQ�@�"�[����-u	�ي�݊�߁|S��܇����t���|'.Oa&�D���@�6�f��q/`��Z�z��֪�Lt5�{�������_���!�Y������_9����U���+�Ų���ӁͰ0��N �wMfX\.YD)��koŖ�NV4:ut41|�S)�!�6Q���&�x��4�,Eo���H\+�F�B�S}FE�\Z�:*��\=���K����iX�?��;H��<|���u���y0�  "$� �"%K�hR�,˫��v�۽��=W���Y�뵵�h˲�`�E*�""g�`0���t��u���릱�������TM0��~��}�'��ȣR�A�3��(�	v����hvg��g�͂P��-ؽs;���#�3��%��k?����R�wtw���IFG�p9=F1�dׯ��������]2�(0��Ԇz���KF�!��\>	�al6ń��6S��1E���\�1�^�Ŀ��nN�J��B�l�Н��o�І���e1���@ʩ�`!Yg"9�HK㳈�,�M(�,lւl��bZ,�ذ����"�����H�[���	��)��a�+�˴٪I	(��Q	.$�؉g>�	��L�͊� hn
9�sL5DB}�T9�5��*e��x�[���M�Ws�m����� ȆM�OI��R��]=80H��Š�#'��1����y�N��$F���E�����L[���ף�����d�%~V�ŉD���\���RT�|��9�Un*��΃�;���݀��
��.�<p�&e9*&3�bx��U�.���T�<A+QҗY�F��sP�� ���j�bW_;�������	�l�ye֤[��m�xc�F'��X��X8�e�M[���6�-�źU��wy.�a�!D���6d�e$s�.m`=���S��f���<"�1�)���7d�B��ҼpaOf*�g0=��D�(��N�(=/Ԡ}�]����d=�6��[.j�d+�{1���Z�'Ocv-w]=T�"#�Y̛a5٥����}AB�,z^�ʇ��Ag{���ͯ�blj�k[����d�ߧ��cⶤjV�dEpωYɘ$����04�Mr	H-c��+L��iiZŊ�p
o�wK�Q��A0��8��������+"j6��eJ�X��F����)����P=A��I�v:�2h�p��~tw6�ZO�1���u�h�h��x�<�X� 3��Ϡ�k��n���    IDATFo���y��ͬ�)Hg-،�p����g�q�_x�tL��!��/#WLK�4�ͻ�;ѳmb�Μ���#���
��Rʕ��!���>�u�_�\I4KrV�" �9����u�F�(1���B�@�(��YK��y)�48������Y(D���1�ŵ��3��*^&���I��%6�����Iem�@���	����j���I�q��~�@�yH C@��&Re��� ?�K�IM%�r��uY{͜>�����5.�U�Fg�CJ&�D,,{Q�����4����4���2��Sh�a�[��`#]2á���o~���da��wN�����4Yy�CطsP�`iTĞ6#�ߠs$��O�D�ˆ��x<G"�#�&���ԇ���FN���ʞ���$�ߗ��e|�S���s���ߐ�ɧ^�$�����01>)+�����?{]�}�3��}��'��_|Q�ǆC`�������Z�Al��anj�tn��
\��U�B�u'4��}�I��:�k���-|��7�ʻ��U|��=Bq)�#���x����ǿ��&�y�=N�E��[�`qs�}�q��oC*
��-H�3:v�lE��Ib��Ǐ���6������2��0�u��Տ���B�L�;-���MFERA\
n[>5����O���%����G(]M��i���/B|���S(�ҰS�+����1��#��Ƥ�"3`x�p���
�B��SN���<�Z���i��. x	���dz2���ӊ\k�����z"-Bs�i�hh7M���j���d:-�i���
{���Of�V3N+�~�w��{aھ�^�+���scSȚ�0��`Ai��9݂����1�&��+��d8qx��������7M,�����_LMy���~�'g�f����2;;r�xA��'=c8���L8;^�1(���M(d�ho����@g;���p��\�]eqB�P�ۦb3U�{Wf��Ϯ`=e�2$(�I7�E܄�|r��58�
vq�>���k�GWyd�r���md��J�����OA0ř����s����g�N�u�a:<�Ӂt!�w���p%7�<5��ͭhhh��9�!�&+���Ȩ�ɻ<p`v���u���~��u?�ۘ�	��hٜxs����.F>��&��8�����x����k�`u3]���Ѕ�w܋m�ara�[q��n�T7lVC�hT�eTL%��t(&�	��-"�� D7a.�a�`V�(��m��+5�7Gx��*D�l����.��&S3�e
L�})�Y
�K(�!PM��?��?��43���f��@�>���E�l4V�����r��!�I1x���@���Do������IFIC&�����.��68�eT�� ;&�ɌQ�_���FEFN��ڄ�E���MA9�CGOk �-q,� �ת�P��`~-�K��1�F�bL�<.�k�6�1�ӌ�z'T+}�F�bw��eF�Q�-�\���\�V<�'��e��|At+���0�TF�931��,zZ���ӌ����i%�Hg��h(����V\���Vb)XL6���N�TH����߆F�CB�h-���5C*'y �o]Tt���D%�)"_�be=�KWF���	��'E&|�wbGOTGE삉�Db,�ű��o}6ʺ���)/Ͻ��G�v�(Y/��	�R��ݴ����W'��{�,�li�ٮ�� Q|�����.�4�[�L�#���*�6G��bh�\�c��>6��p6�q�ղ.��GWD�De��6q"�d��K��#��b��.��э�05�w��Ya����;?"�|��/�L:��5���h�[נ�H�U%���	[���Q�:%���#�1%Z�V
�m���{��+2���Y���k�@8Uƻ��F$��D�
���	��x�����"V�D���&�6$����UI�.Z��)QDS	�S�UL
KJ ^�L����f8��Wo@��$��au��IJC����[	��5��C;Q�J��$	�*���L�8<)ӮH��;��'�v��(UOr6����H���,E"A.�bE)��b�(E�L`oK�Mk��6���O)���S�k4��:���"�m-Ь���A��E0ς�v��S	)��Dt����l.W}βP0e��ײ4c�r�z|��o�KNk����361)_�z�ۤQb�'v�EL&
[>���z��gǑ�;�2��5�w���7�m�x�cOc��>��6;�I�ϭh�j��}�	�QD#�x܃A�� ��!�����w��7�|�hT�r_��o᳟���}��!-�/|w����2�eZ@0���o
���=��G�����6,<nԲ<��x�ÿ��ۍ�Ʀd6�8C�����0-�5x�&3Lv;��y|�>���E�Ã�s���+o��gG+��;Ĳ��CE�?u?���|
LF����ޭ�u���/1M�؉�j���1\8wׯ_���
t����&?q��P��-��ԣ���Q��'�b��A��8>����ni�$u��2W��L��STR9�Z���ΟG|j�H^���&�#�si|�_;�����DL�ي"	�G�I��=ё����(n��nCA]s#lM�@�G�ILR�ayz�Dݻw�]w���H�T40?�u6]��7]\AauӸoB8�~�L�.ag#T( ��Axj��!�a���bE�$m��������q��a2���8�w��D�k�
L%6����,�4jM@VS9K9;q���}�����3zc���>��������k��ڭ��s&#L"<2Rj��hV��kb�S��e��+�B�iV��{��]���"�d�4��P��3O\,�KC@Q�J�\�.�J|�瞣?jXܠ��ݮ�(2^����X�E97�q�&D�Q"�Œ��E�iw��eK,�uSs=:;�q���9~��R,������6<,����/X���x}��/���a�Ӷf�@d�TBsK#�]��p8,�Gc �fxS��8qP�V��r��(����$�D��?N�ngQ��/�|�EL̮CKW`u`����8���D�X�^+%	�2�2��.�TԄ۷������ڄ���՜�4���pť�b2&��B<�Y�#mM�R��Rj\����V)ƈ��BX��OXw��94��~��"T�Y���7q�TA��6%��?G�^uBPv�m��[�G-3��{�i��jn�R��J�T�bC@W��EcЉcw	���x�NjTΠ�8\�5>��K�S،��p.�6i�XPZl`9������Q���&�{m�U�].�KV�,*6"Y\�v7&�Y1!�q�5��z�7���
Ķ��p"W2c=��������� �fw�6'�n�l8!�n&%gt�Gw�{�ڤ����I����q��ȕ�ι��^��Z4��#��IF�2���A��7ë*0SP8=bG�U������v"ON<��y��ztbW��a}#
�נ�1Hl�`���)2�瓈���XX� �,��pI�Ŧ�뵉�ضF�꼒�@���~�t�ҭp���s�����$���
��p
����P]���h���(B� �Pȥ�K'd��mk���>٠nN�!�Z��jL�#8J(p�a2�G:{0��G��1U��v�w�;���3�&v�V�-.9��\���،�k��3Y�)o�p��B��t�H97�\M�*6+N_�z8.�L��N E��m�Ю>(
�FUI.V0���释�oL!���,��2J�,"�kh	9��Ç%�^&�"T�
�hFV�!�S���a�35�J�U�Jp;=�d9	*d��:�:���)v�`3���F��G�9��x�f*IC��َ� ؁���!,&xU����
.^����"re��q/���6�wp�fQD�ς/OJ��� ��[6R|��J��9�q�k�@MOR+�k~�RēҐ�!Y��y;��Fz�~V�Ԛ�?e-�m!����42��������ȟ�^4�G��ݧ��)`��̣M���WJ����'�fjnN�I���F3@*�b��!_{J���R81ԏ��q�&z>���7�g�����x쑇�P�C" �Ev�X� N�y�T�[&��C�_��1t�h�;֖�F<��#��c�1��w�F܂�<��}�w�>�����w����ٟ	�ǩ�=w�-����M|���{�w��������g�CGG^}��x���f�l��!b\N��^����A[Sr�	yR;�
E%��D���Ť���M흀�8��0���|��}mF�=b̑�/��ц��_���`a�h�{����K�������4tt�s,�Έ~� '�%-��w��/<��m=bLJ%�2�$��<�>;�ӗ�bzn��*v�u�3�x�;��ہ��5a5�Û���lhFС�Ò�!7?���'��[��PD��/�!���x�9�!}�a�'�'�E1�Fbe�Ur1\�&"&���}���ɤ��g�W��duM�`
�,�+(3G&Bѯ"NѲ8*��U8�d`�P=N�8]��y�:�Qt�� ;z>>ǢQ�@K6ln ���ld�\�dvN7��X,"C`�����:ǞX3���o]���	�狈��H�,J��,2�L��X�MF�!vߑ������������xC�_��㯝���͒+h���B7��I� A�[s���y��h�CA�B�*�&c�p���+�}-�mnB@��-T�nhm�310۝�$9�Z�_~�M\]G}�^iXd�a�,�bf(��2 ա���qi��3�RaiH���cwR,��p�l�;$ʼ��}�{����N%173�υ|�1<�����h��x��ױ�4��LNR��:����'�}�$F�]7�jZZea�C�D���8r����+H$�%vh����֌v�j�J�G�� 2!�Ƀ�LL�b+�BCk7z��`x"��������d�
���������+�|�depGg�۫��P�v�b���G�H��c��(]�͜A�EY�П i
��9 ;Om�œ@��,l%%��!ŖUX�V�
��CAC��3�;���~R�
זl:�h%ES���!�P���ZLP���x-�M(���>ݒ�I��*G��)����7^�%�f��p��9�-A:�~�'��I0��)|�h�dV�f�]Լ~��wc�8l%�u5�Cy�u~/�Ad�r����0��%���U����qذ��	C=�k�	'T�d��
(3}Ru!�W�����z���0��%V�F��r���H��11�@ո�J�,TKQ\�����~�Y��"x*(ea��qitF��k:MyP�g`�q���m��S�\��qv J�Z��'S c�E޵V6����VãS����# �0�w�]ی�R+eE���ƍ�3X^Kʤ�E���@c��]M����"���Q,��v���J�υ뷰��@*_���X�ՎR��1��`�i�¤XѨdPP�VB!��C1�Zĉh�X@���-vn��0k���RPh�&Tҙ�%3K(Ilko�m�uh�M�d����c��ZK[��ES9��.�����R�����ط�]��x���OB�����02���~yZ,~��z#m�jE��Į�64s���n� ���o6�ܚƹ+7���%N\�2�R�lm�!��ɇah�Kh�i#D�+t�p`t<��SX�$��	ba�ˉ>��NhI��xU�dsi)����&�Z�2ĬR*IR+�%�R��e�1�Y'>��!�49�(
5)lDs�^���s��ȗ�~Eq��i|-F;�/U֙�͈���N����o��C���TA��zJG����$���6<L�Th���NI�%F&#��n$��d���g���!Z�C��D�H�%������F�A[�~Wg�4460!�ڀP�$�F�T���&R�8Mgc,��ٴ����u��Hr��m��報7��������mB��x����3O���.��>{����	�N�B/�05=-��������:���EP,��퉈t� V�,�:ۛ���`�;T���ɛ���'���՗�(�⟽���/�B�Q��=����ocjbR4N�%t!���@Pd���cڃ���x�I'z��'pǞ=h�0;6��[c����X&-�A�I�45�d�����咯�P�� �n,n�/�~~a	�YC.�{L�$��|�G��c�¥�������?��WǱ��
5�H�&"PF��z1�;�8�/񷰧ǏD
����܂L�n��av3��H\�Xˢ�͏}��I�_<{
��⧈����܀{��CwE�b������k�9��5x���f��`�b��`^��N���4f�#��'�ͅ�H-@���AG1��l|�3�k��H��3O!�P��hW��̈́�^FN�_JQ���E�Mg;��G�68N�;{$�SDK[]�ׇt
��u�Ӏ�df�j?�u�8qw����@��q$<!�v�~z�
V�D4`#�GI�Ca�,M"H��2���+91H������+��o���]C���ɟ��{�h4��^�d���ĉ"W��33EX��RB!O���8�7�����@>�Svm�Ů�^�Ȑ�2� ��W���ؼ�o��[�xsCrt�[Dŵ"���T)����~Cp��[Hl�@c�V�!0��y�fp1Ul�	�⤣
�H��.�s�������������E]�!����~�㗑/dQ�� � [�L&+:���� /^��q�˩��$�D")j��:
:556�$�\D�P�F�����a���p��ゴ2����+8{�2|�-8������~�?��I�*��!4u�F��!�6��dSy�ilPU��BI���,�|Nڅ�N�a��5諳0�(<��R�eZ]�9��	�n R" #�dc����!/Q�Vl�*BN]�FǣA�����q�~<���pxT�//�S��4��X�0ʼ����J�������FvSx�O��ڄ����6���j�_���0L��.�CCh��a�+'+eC�N'f[�,��N`|v	�D6;��jp�D�g`5�"�mo����E�=��$E`p&E�JD���-�u������ց�V�DRR�1�6�ْ��2F'Wp��-$��m�$�0d\���MJ�i�vŠ>���f�{�۰��u.��w�`�� �T�y��<:���MY�d�@��ӊw�G{��� ��Py�S��/uA��Y!�ɰ8��l:�a+����
&g���{+�	R���9�F���jL�UK19�&������~�6���8Iᰉ����F:����qA�9f�6�K�$D�D'�Rt͒]u���~�,f�0� #%��mX-yL)��� uI�U3/�1���� �ƥ�%<Q��s���Q���`/��;Q�"G?)c<����h�	��v�dAha�6�F�s[����+$��R.�hd�dn��&q�9}�"�����C�PE�IZ
�ʒ�A�QU�������[�E!��FѸI6�|&�T2��?=�{�;��r�K7:R�ؔY1<��#Xڊ��&�j3�>x��I�Dx�������WdB��Qp�h�������ht-�������}t^��|Foj���ln�ob�֢�E����4U�Y��p!�ÄH8���MYc$���Ⓣ��S�3g)����r&�e@V���fQ��jr)�ǀ��'����}zdբ�F�	��܁��i��sJ$b���]]�g� 1A׋�x�Ō���ګS5r�(��')w��l��Kpi{�PT��ۼN$c��1,̪�����p����w⷟}w���A��/�Ͼ�q�;z�iF��193-4@������rQ��ghV�g�F�]55��}x�>:| �s�sb�������2Ƽ�'>�A���[��׾&������3�<#�13��k��8{����@�������^��$0��b��婧���}�r��~�n\���;U�8��ѭ&/TJ^?.�_�-��li��Ҏ��A�\K�ş��k�F�ѽ"*�DE���N�G=���q�hP%z,r    IDAT24צ��~�_�A���[Z�R/H[�lZ4!��]��>���{��ZJ����*�����5�.� 7a5�q��a|������k��#�L����G������@iq��X����&�`7)��6����V'�ȲPQL��x�"KKp�e��U,�ZIsn���[�p�S�fmWd����T�U+�P]n�%?�kr��V�,�Cm=����+E�2ӂ�����V�Kt�bj2Y�:<�~�S!/4:�7m��=b�bF�jA��B���h��!��o^��߿}7W�X����
3�Bk�@��؂�L5`J)�k��?���o~��W��h���~��^�Y�o�a��nǪ����U���Aie���F��,S��Fس���y���|�E���{���S6���̴cs��ZQ� ��Ƥ!�XοLƆ@lF͆�Q~A;M��ç�2!~��FC�	�� *tE��&�"M�tv�-�y���u�c+���c[o>��s�����5R���<^��Kk��܌B����M� ��y��{�ލ)�@�͆����X��'�w�^�n߸���7���K&���;��C�J�7�d,.�����d�r`p�1�r&��7q��,2,p��Zйc�,"���4�Q�l�+(������еfFưx���I(H�(P��bJ��e�O4���1�j�,�! �KA�b�b��2�Iڬ.�&� �n��8<b��9����T<�8�Lΰ4+��0J��,��o�2�O�	T�kH����ͷF�}Bp;��Y�|�Z���� �{w��=�������bC�d�����5�<ܞ����D����q��΍�ۊ�/z�\L�$=�h�re#��.�`|a.wP�h�Ә����u4��EL�~NY�L�r
.^���Ü��n�5(�m.�Ɔ@��P�x5W�E6v���ی��-2!h��ol2EH�4d�fl$��82���E�+�1"��9��]���%���av
�I�O����)wc���G���6;Q�Z�d��f�W0��%����{qh�Nt���Gg,���-��<��eR�hu�#T������kAO��&D��<��#cڕ-��\����'To6�[
%e�H
#���p95��mYoH� U��7�S|JN��J*+(�	�&���b#ː=&AKfVɠ���x�+�rPIÆ�4�݇z��J!c���]�;�q	����6�Q��`h�=���N�S�)�L����)�����[Z��i�A�>�BW[�dU��Y�f<���9ܚZ��V���U:�)EG������2�y螽��q:��`�m����Z�ijE�1�0QdN;\�5��@Wo�H�����8u����L�t�]����d�����3�"�֠����ݒM�����Q:_"S�T�+�T�`�q	:bآ�1��q�ɔ��t�!��t6RE�5!�^�Hv���-bm����$��j}���=��Z��f�?'������&0�ю��f7rj��l&%nr$�B��tZ>'�*�#�6���p�D+F��JYl�Im%}���F��	�)�Y#�xF�a1kx����ۿ���蒢2�/���+��������	�ǭ"��a=�eP�vI>&��|'^��H�tR�_"�}��@��z:q���{�	i~H?b�ط��[�'@�.��=��[�я~$I��|�s���� L��/�Ka<���x�t�N�>��#,`��<�����'����{�5+�~�.�:�R*��.�?K�";�I1��0�d�b���jES�LG�����s��*~8\~b�<��%|�ރ��'���:5M1�����^��g�#I����baZ��QD[��a����to�#됉��lN��� Y�T�t��A��1�Me\<w�t^����8<ЇG�A��Bdl��א��B%��5_�E�L�"�o�(}�І������H �����:z	n��QO���)Ф� �Dv�|Fv��W�
�WF�,�$UZ\��Y��
�M!��4H! Y"��ʀ49^uD�-
�ZIN+ٜ�f�r��Ow@���F�����`udt ��P���{��?t������?����Zi�,����D�d�1����*���=ۿ��?����Z5�?}��O���}j#��S�~Rmk���wɫ;+��E������ؘ(I1�E��{3S2Y�������X]�ՋQ����Νh��!"���
��ٌ7ޛ����$63*��>I*�!Q�+[�Y�O��knHC^��ȩ@|m��&�%�JJh ��2T���v�ai�G�.�Ć@�;R�ޱ�}�Y�n,�$��q��i�rC�f
2�'��ر��o�.�ꓓS�F⨫ɢǋ{hh�9�Â3g�㭷ޒ�Y��@K�O~�1l�ކ����el�#�/�[���&f��`pl$Q��̊�UO�:Ѿ}�d��M�&���+��UQ����]n�@,MLcs�ʛs0��E���H�uf�P|��ʎ,��"��11��V�6;�,F+f�L.Xl�?���p$��b	�RF�ѽ��ouM��]��*��y��1���%�¾TE�D�i����ܔ	��q�B�@&�(XUGp;�6t���^�qw[��wnÎ�:qB>c؏�aF0��)Mh��$ʠ�G�R����t�l��Hl��s�(x.��ؠ8�،��Oadr._ N�!�����h���4�-�)9(&M����9݅�x'���Ց)�s,
\$�R޿�w$��I�1��,���N`����w���A))*f�M���p��(��Z@��-
4UD�zd� ����
���czfN�A���G�]�]�*5D��d�Ε������6Sb��
�����v���MA���e\�X|���lp5�׹�s�{�;�2�TH�*�5���d�o��
C�&0�E��YQ*[��#ݑy,�t8�v)��|I�Ȧ2�ςR.'�i�U� &�,�����LDpǩ@��S
Aխ�u'97bJŝ� -�^L���mx�{P�t��e����U�.�g*�5+���T_:ښ$�E%��
f�y�%	�7��fq�ʰX��h���C�l�#�	���r`bnU�	+a�ͤY���)�$D�����u���C�򋑩���E(��q>֕�Jf$��0� e��J����n�DGG��-.o��L�.	N���$��,~��^���~1��� �D_gr�8L���ְL7e��KNx=��&�K�Ҷ$��[�Aw��.�x,)�)Z/�YF�/~YX�}M�*�RP�*M���p��T���W&�"�7����5����j� A����W?k���.�����Z+��K�}S�8��J���bX!Z�����pɒ&��M��
��'��Ϧ���L`��!Ј!/4Ҍ��z�����'�o=���!�O���3��᏾�Uq�ڽKlf���Pf�MI�T&+��Ԕ�X�)����#H�b�A� �*��u��=��C�eO%����/~�Ν����@��P��̌L>X�?t����a����N�<)�|����񜛛Õ+Wd�g0'�c��ă>�m]]p��ũI\<{+�3�|�I��n���Zb���M��ƚ���P<�}��������cЬ>X])賙-4�<����3O�M����f�������1~��I	6��]���~k�Z��V�e�%�Km���9�4��w�h����<�bZ(�A��{�BS}�Ъ�+�Cuh��ޢ��ㄿ\Ajv
�W�YX��"c]��j�@X9��"����]�>�E�VP�
C��O���&Db�e:D-!u>r��_�^��PrX��aR8�9��A����5��c7�"�4�P��~ev�jC�\@<���#Ќ��2��*�.�:\^����������.i��hn���~ J� �M��{o����ͪJ�&i��f�$�J�!�Y��������_�̯������m��Ͽ���x��/���qܱ�7.������azj&�P|�(}&�Γ�5�R���W��X>��G0?7���a�>ڳ�u��:U�|%h���*�<5���"�� `iEYq
�^K*�PkT�	^8-�4��N#�<�l�	��"o�QA>�p`m6��t�u������)<��	<�����B$� �1�R������<�@{{�L��,^�`����-\�tEf��&���I;t��~�ϟ7,�v���!�D���=w�=��F��aiaQD�MM-P=^(3�k��K�>tQw�3��RV����h����h4݊"}�eC�%��E*c�sy���-�ckn
���� J���3�&'Q�,��V��1J��Fl��Jż��|��=�t*[aW\PLv�M(��͆-�Z%tڅO}�shhm���*7ո���&I{[)��@m3����jeA��O�m����� �vn�j.C��4U����������V��Th!iA�l�}RZ��oV�:�ϗ��LA��6+��["�U3�|n�RȪ�8�X����Oalvv�GVA�ݱ]��e\����p���6��5a|~�/���rX]�3���� q�+�������	$I�3��S���F���!�F�[��)�L����K�42�L�,�� �z'�܋��(z��>#�)���8��� ��ߏ��>�U�o8��![/|�JNͯ�������C�����A�K�iW:1��+#ӈ���$ ��z'�����m��ʰrC�N�$��T7
��i��6���4�"p�9�D�ͩT"5��tyx*B�~���z�l��nA�"����0eچdQC�X�}n�)�Y�B=%:-�5�]6}�%�]+�ٰ^���Դ8LZ{��ăw��g��2łx� �����J�x���jhDoO�h.ZC>i�	��T'��4�bVqsb��\���.�)�Ю	�#-���lM˥�X�J�� =N�R6��~KC���kCW�>Ә3�Z}���z=����e�rE$�	�$R�P���^�_�����N�5׮�ĩ�W�/�P�Ԇ��E�wy� �c�n��#��K�`>�iA��t�ter1&��V\C��oj�D\��Q84��H%�K�c�A��dR����gI�g�,i�Db�\�ŧf1Z�*�&|�����6	�(cՑ�v��Rh\�մ�ꤏS,I�L���Oy�e�]�M9�,���c6Kc��$��K��g�N�h����Rƍ��X[[1�M"�l�t�&�%&��|kV�DO�&.-ӻ�~�����i%�Ű4>s�
~�+��X����nGGgv��#�pT���%l�����(#�B:����	0h�I���>�I4SP.f\�|���wp��e���yc�����>�s��.'�Լ�8a����v���k�J2�c��C���������jG2��ӧp����1����b(�J���x�u���'X�:����pk%�������YuIÕτ���_��OੇN�Z,���`jq���o��*R���rH1$�.�<g�sKe*A&��،r���EĽ� ���$d���.<�����'I�4vq�v��,��F�^YD�Պ�^Bx�
2�s�d��2g�6����X���t���8���"�����ȭm@���Z%���|^���CqA�%
������Z�P�Y�� c�� S�^�.�a���u)f�y�%���q�<2٭�5HfҒf�sA4>7��ꀛ�C�3#���>d��r�T_�����nt����ݸ4���~�oN A�9�f�,	�jeTh�O�m1g8饶�����w���������_�	�wϜ�����7��p����[Oݎ
S2�:%��F�,����)��f���*�W������=�k�/���5�vv���!��=n�0tB)��p'���h}u�C7�H���HS�D^#�����X*ii�ǯ!�<�tl�F�y�T�k0YHwQ`W��b�x��O[[S�p8*���1<��}�=�]��ٳ������"��o.����/�!�e���~����Y\�6,h������嬊�g$ҜE���
67V��hlb�P��������M.>���Ǧ�*����f��x��T��L�_]�w��l%rBI�IY�P�͛����V�P��@)�Ef3���[(E��n4�yf9de���g\���F��mٸ��v���O��B��?ʌ鶹���ì[�b �n7���n<��O��)�����o	�D�)_.JC��	��v̾���d
@�&�������Z�_���n�D����k�����B��:B���ok�iaqU���ņ�fE�#�)�sI"�A!jjg�5EA����"S�a�'<�2v�� �8甁��ő[X
�$�|�z�O���y�%��xQp�
�t6ܘZõ[��H���r��K�oI��J���b�.�!�R�Оmm�D�O.�B���V��ƍD�'16�&5��\*���G�C�-HǢ���T6���M\�>*��΁��j��c��e���㓦(�)�&6�Y\�5��5T�I�$��> �m,��j8���SH$)H-��e����у�Wu�i��:[q��$��M��y3�Q(6�.#���㢶`����W�u��{{o�`�(/1Z�!0ie�Ҫ/�� ��f4�l䰰���=����2=�y� B�/A�,IE(Oĕ���8v`@�Œ���&&�V8��Q4�Xي��w�`naIև��^������ȭg���{lJ����3�|uѭ���-�ދP���Hќ[�`xbK�a�4E�����P�(M��İ�.�CC;���m-�X ���I�L^G�Ӵl�2�
����u�A�2�e:�5��[����. �)p3���i*���\Gok O�{{w�����e�v�`R�Rk3��צ�E�*k'l�$g���]��<�w�g�,����	5���f�WD��5�&L�cٰC���5���.k�mf�C����I��-����L���ƅ�1>���� P6.�D��D��"[N�ʒ!n�f�����Y(r�Μ���<��r�t��v2٘YB�4r�au&��z^x�)��'���ES�O���?��W�Ʊ����ƾ�{�F����Uq����C4����u���E�=�H?��Ɔz=t��tw����<�^}�U�N����1�{���!'y<��ukQ��������d$횅<�26Y�M�˹���űc���`��vD�6��o�����M&$���&�R������|��9dR4��jF]� ��,�ۯ���zC�(��fSb�g�6|�+_��w��"<6fR s�Q|�{/���>R9j9-b	�����BOW'��L��[ayO4D��bU����=�T{eND˕v�o��>�;�R Y7U�4fcq��
f�\B����8����<�3���
�X����!�4�k���B{[����cH,-é��w:��5 �{���C1�5�,v��:��]�<q�z�8>���9he�ܗ��9�
J�"ss�2m��Hڝk��S����n��Kb�m&���`�<gZ�;y8��`�ƥ�e:�|'��Z�@0������}�)(݃�8����>��nLbK+#V(���I�+��Ć��R��E<�����8�������׋2��w����o~�
f�}�>��ك�S�����pcr?��{�69-"#3���^8aC��	�����N��s'q���܉����Gt��B��=�]bO�橛����HC�	���H@-��R�����Xa.�[��/M���0lGi�h��*A&D�dto���6�^�C����z7�����#��{�n���t��\�$c����pt�T^�tw�
-�7���{���%se+,)ih�{��%�N�LQ^[������2<."�n������v�i��[�s8s�:F�����J�~�^I{݊`qԡwp�4,��YUج�?�ÁU��F�.�@��l$�6�!�Da.G��rB�&VP�qR@n)on��-1N��0    IDATW}�A��9������&;�'J�
l�:�wl�{�d4pQw��86���������p�i3HZbě�.��Q��+�h �D�ǪkF���x;'���ZC��b����r#�2K��d��&%S�`zaE܆
NO� =6&aq4*�h҅TYd�~��@e����:�Vd�)�&gW$L.���`F1W�z��C܉��UiB	[G2�F��#��1����|�[Y��S�!�q�-�֌�fNY�� "df",i '@ؿE8L%�ؿ�C;:�%��t�,S���Z����֢L6�yW��hP�IC�o�Z..�$�����#���vw

H��eG��1��t-s�b�#�c���Els�:��gg/|~�ei���%\�>�~C�4�:;<��v?�E_YY���PkS�(�L/���W��J8��^�8�d�6��@�հ�"ݦ�яޮFt�7H��3�V�;`*���ʗ�x!�	�q��4,.G�ڒ͠�0،Z�����P%�.�O��&���L�J��E���pt�_�b��ٞb�p�h���p׮ݒ�Ng�}h�w��Ή��O��y�-X��Fz��\3�����2|v���A�
�ςH����G1<>�X� ����`D!L�}��
�t/�������e+��f���r#��,�Rv��̈ ��#)Ye8�N	��f�7����@�|�.����a	�S^��~y~!*VV
HF6��шG�>�����5x\4�6��j$�S��qyde�G(���Z'&�	��5r��TC��ɤ��,�Y,��QJ�Q�p�[�>��5q9��b��gm:p;0���4�:�kj�5��Ť�xG�-�@.5��hM��x�O���+i҈J<dCd�F�@�o�SDP*���I�cgN����l��1(��/ـs����*�__:F�Wŧ��0>����-$tԼ������ݿ���:��[p��c8q�=օ��5?����	��o���{6eZ1/�<Q�,mGu�A��5����8��Ȇd�>}Z>�[����ԟx]n���`"� A/�ך�_kv�<Gy
���4_�C8�/|����c�����?��_�*����S���!t���㢓�q���jj�A{�^ܘY�_��
�>se�UE��E6����~y�\��(�!�K݋�|�[�C�~��fQCKk>�O���E]�# P,�%��5Nɾ`p�@SC��}�-�������ׇ��f4Ndl-�c��i����r�`g:�hDjY����F��^��5���i"����!�Arn
��J��;�⎤�E��+��t�����e4�@���Z��O�b!�����6�	��sH��b���̭����TF�CE¯�R�U
ԏUPd�E����)^,�9q�yfsB`Z�����7�h^�!8v�F�cZ����E���e���Z&��d����#���4�_-�ȧ����{}��������_�EmG����������V����:���V�3�;{B��e:���I���Y\��Ս���Z�^�S1Q�?���8��^��֦f<x���4B^��<*D$-e9�,pN]���^����C����!��,"xB�:�E����&n����3o#�2	�� ��Q9�y �8��^����D[k3C!�4գ��G��¡C{DD4�0�x���w2?�!cL�0;v�X���đ�a/���,�
q��
n��D�!G��}�XtS��G:�siI�o�u����䩱Xf(��k����XZKb+Aj��f��$5i�����ӏH2+�+'"���S\�.d��t�b[K����@ۚ�j.H�EI"�5�TtUn".@��6�_:s��ǆ@�w�bL��܊��;`��s:�&�������yq�r4����觞��eǍ[�Pl*�����L���&f]☎(�!��M�p�\��V2��
�۹�5��f�����jb�Q�Ru�4׹$��|d�u3۰��p��hW�`����S�ÊT:+HBc��\
�t��-�nA�[Dk@>����������El�X4�r������ػ�]M����P͈gRиx[�X��06����5D"9��Ɔ,���i�*c�+%g����I-iy$�����ݞ4>���Q��Lg�<�b#�|6�E���`o3�W�+1�[���Fn��x�ǡ��YB��(LW�aX��@Ew7N[4�GF1?;���:��&��|�,�R��\�D&kԨ��k��Gv��QA!�����"���16�Y�'����Ī���&T"������*��	�at-�^�w��% 7�J��ur�s�M�3UԐ,�qk~c3��������<�E�={f��0�  ��"V5��$۲��qY��ز�z����NVrn~�fݛ����%��*�q/�U˲$��؉F�����^�z�o�������\K�9 f�������>�XNy�<]��UU�+G�j��ƺ���b�#h^qw�@6�hx����H��qu��Á�h[�4�ֱ��%`_:��8-�j���e�N?~N��8 �mau�'�0?� ��oQ25Y|&V�vqebs�Q��0՗֟��ZU�+f����R\.�1�ׁ�'G򐎙�K�VO&se9�9Xn���g�8=h:��-e��6��XO��^�4
���7,��Z&֊��\�<_�p�9:$.�Ԅy��r;6w�x��C`xZ���Pf^��|R*e
�Z���ޱ��t�{�I�!�1���NU��D��㿛�V$�����H����̈́�\������>|O,����X�s�M�$݇�r�z����ɜd�7�=���i,x�����=�GkSH�^:/r�ܟ
H&b@&I���
�X�F�:�*��]V���߉����a�'�2�"O<�,��/�;�V�܃���f�߇t*#V��s�H$�b@�����H#����b�X�e�x�o}��N��]f�����5��:�笀w�~誱4��n��6ߜ��۠��kED�Ik��y�	�����'1�/�F���Ǟ��¼�b<t�����9V��ft����q;�b_�)]sk;��}����o��x���(jttt"�ˈȷ�����r=�!`eP& 	���͇���p�Y)������g����7��,��׹��Tzz���<�T��(�wd7�W�i���_8�/}�2-�t��I�[+c/�r��y�ݰ�c�T-�VHWT@ �x�֫��P ����%�3i���#%��'���ȴ@��<Z�����҂�o�Fs36���۬�x`���KX����~�2l;I4���)�5T��)}��Z���J��Q�� ��M�M��9��M�>��M�~6&��6��>Ԛ��KG����w��^�xu������o`i'��WU�'V�E�A+U�(UU�1s��rz����O������0���׆��ϼ�����W���l�ۻ{�z��;p��w�#D��nn����Kx�Wg1����߰����䱛𶷽�'Fq��y47�q��M800(�˰� ��@�h��(~}q�,�e�O��%�5�Pr�u�6�X��.���^?��їPOn :��8v���yn��W�����EKs^��{�9�{�x
��~�|^x�y�}�<��a��1&����N��7�`(,�>��iJzo��3ʕ���L�䡠ƕ.q?X[ݐ��)���0*
�2I%�<v�P��.Ҷtjq��N`ayۉ<.�΢\�-�.�q,�9��7w�f�"ǿ��ȗ,� �Ak{n;Q��\6��97���*t-��44�O_���a�S<U�tLaS�1���]B40��`B���G8�	���$�Q�`�\�� ����pelR��8!�����H��MhD�\4F�\"fa+.!^mE5���W��(�#{S�g��9~f��m��^�����%�� �ӹq�l���?�d����FM#M��i�t�Z��_�u��Ў�{��!�m���)�&��x����u\_�v�&���&��D�8q` {��ඔ��6��b�C�⒆���2��-"������T�FV�&Xhv�����W�Y	M�i�����#��S��RPJz�1��zc�<{[�
�VE� G��Z��r:m �[䫯�������)$�8{{:1��=a�4�%4�AA���V���$"x8��:t��`���'c<S��j
�M
m�����$���-� *����Tkr���(�.#]Ա������X�J�fw�����")5� ��W�#�nG�BuN��7�Ǳ�0��L�� \�nE�X��m��_���k��G�=-s%�]<q�׬
/��Lɸ&Y��9e�Ih��ƽ㍷K�5QX�W��<�6iܘ[��VT����[$P/rK·�^����?�p��Y�[��-HS������hmk��D�-#͆���M΋n�y�]���p����:�~�t1�o���#8u|^��
�n�:jQ8� E�\���K�:��+�t�<�>���|�׸t}.�`��i��^R���X��JI�9y���KgPQJh$</�^3��L�^�:�WF�ETnp�@Ђ�1fO��IZV��W�be7�}�@a�7����녟��c�7�&��Z A�Y�H�(A����:>�B��4�����yfހ����JM��*���; ֤�ڴ'5ir�~I݀N1=��r	m-M"J�t��C�"�hwg�T6�Ns�M���@��\�2r�8�Z~�=���ɤ�9t�z�ٳ���"��MH���a��ǝg�H�)2�����҈e�9��c��4��>MN��`#��z-҅8��� ��T:��F�������(�L��I��2Ch6��� �a��4����'���&���3X]]�07��ׇ����N47�i�s!��}EZZ��aj~�����/���A��B1���Z�\x����g>��9�i�_�8��}�a���m����6���Ͼ��p�� ��.�CX�����U#@j.�t�v�_�!�f���bŹsW���_/�-���GO��SC�ni���F�ˎ`�WU��5��!�H�]-�cN��L�RA깞�Nx,:vQI%j��Yg-��{@@��X�ޫב&5��D�5��U�n<��J	��~��;e���mѱ;1��W�T!����\Ar�X�����cс��K� l�����Ks�
�
�S�n�TI�(��Z�(���w�ZN�;��%����0:/����!����4F�sW�V+�^L��>v�S���g~�����_��n�z&��&x_o'�Go[��vb�?BGU�y��-������!��`ycs�KȤ�hk�`��N�U�ae�w�5�'r00����_Y��lK%�u�$Y��:ڰz�al��2�t{�J�ޜ����ؘ��
�̉���אLa�Bn�>�Ve�����Ǜ�p
���x������ ��,ҶH�Ѕ2�"Ξ=/�E[����f���%�)v�E
�L�W�P��������s��cJ��6�V�nɦv���̗��+Xߊcbjk��6�X\��X�7{��Q8}-���ԎtcD_՜r���`s@�9�ÂB.�f�b�S�!(m��RM����������,@�fQ��B
㎩�hxY��!;�3��Цi�*t�`�>o�ע�&�&��}�Ň?� ��\�T\k���
�t1i4n���S�2֧�s^������n�&�'�LÆ�_�f@�p~g�E)Ď�Ş�&�]6T�(J�����v�=K�Hdi9HW{#D�"�ݰ��J�C���=�"���c��Q���|��x���6��p���ZEgK@������"5.�΂�RR�ay7���\�X��r��##]6��G�܀(8��W-����Fe_��=����ge���65��6P��2���^�Z����߃PRan�ž�6�_�(T*�n�191��5fl�u�-5D���#�fP�����ʼ�l�JȦw䙥�fu����(SK;�]�n*�L6�VDww�vC{[�Ҍꁝ��h+(5d�6l%˸:��˓�!����DGCTT��< lB%`3V+gE��е[�����
P�^I�E[?�H��kӸ��2qK�8��Y�&Q��E�t��@�q�X8x�7�X�ZM�Q���{1���a�Ņ��a+����9�^����p��4���xl�@���,J�2
�2��e����U�./"�A_/*�t:zխ�Y������9�l��,���#���S(zB��4n?1�7�>�N�ȜX�9],Bh�W�Zt�_�Jck;.c,�(f޿��Mp���B,V�K/_���)9Dm.����dY,viR'Q�Ġ׳��Λq|'�6.�h�`��2M8]JdK�\�F�F�<�2��]EDܻ�c�-��0��s�7p��4�m��k�J��c��g��e�G&�X%��ј�(����R��Q�6�?��攀A�����fC���ϯ���*NR���Ig�zM&��.._|�(l�M��9��'wQϧ���c��&�4�ɡ�W�NK�����>����6��ٓ�<���C���jj˴}_���/66�8[\Y��2�'�Ż��eym�aQ>���,���@� D-���˹�Hv�>).��~�d#��n�B���r�.����p� [5e+��E�@V#��Z+�P3@�(����6�pz������G��Iݹ|e_������kp���;���6���c����;��e�����}�a���!S(�v��N!�Ӊ�|�x��߉ps@���nLBN;Z��ȉ�E�ynGҀQS���kF�Zr��_�������ʵ1)ֹ�v:u������"Z	m�>;�ݵ&M4A�2A�_�Zxݻ:��'���bb�lv�I"u��!�m�&�A�"Y�J��Mg$՘���+{���@+�躵�%��ő���d�P���n�{>)���	Ҁt��/U�՚h^�^7JBu�>�7k������==�>
��c�[x��I����^���9P�(s��U���4��t�����ۏ�|�����VM��˳�������;i�E�6*��D^������#�+����Z̃�g�]�%ːd̩���tE��y� �e]��^�Z1��Ǔ�Oa|>���u�'Gk�=�+�="X4��UE9����/ �4�J�:3�6D�>r&��9h#"��M������ܧph����B����Ol>�$�)�"f����	���
8x�0N�|���L���RǾ}{���ӆ�v6qG {Î�ְ��+�F���*c��n�v��T�˫؎��-h����#�I�Ӎ�e�M���mA��Q�Z���HN���� �"/����Vo�*��-����l�Ϡ�D-�˨�a�P�o����VL�Z�H%��Q7Nk������M�o�
5B��C���P��anmDQ�����ӆ�ۏ��<A?F''��(v"��vc��c:��Eu�ǚ�!v��Ў�R�]��81(��OC��ڑ��$P�,��2�N.{��qpoZ��bZ��͎f ��bfq���	�����zV���R�Bv��ְ�m��@��6fD�X��p"_�19��_��RL|޹.9��l����nF��
'��Hȕ��nՂ�Tӫ��\��fV�)�h���{!�1����%���K���0�ۆc�a��^�[�����q��B��kbٹ�(�J]��e�59q�@?��D���i�g.���
&'�����B���'oFWG�L*�Ud���I�R��r1#�,�RjV�EsLd�_A<��(�R>)S��G�q��C��O�8�qʔK3�SG�jC�����y��:�D��/��P�sD�')6ጲ3��7��V?^w��K��Qc��i��V��ynEi��6�2�KT+',�6�i��y�a!�_< ��CV�d9�:������6�rdH&�*��X�H7���.2�w���p�ll�cn~Z��{���R(K�7m�3�2�����]���    IDATmB�����jŵK��^�n�"'�dUЫ�T��������x�-�s�W��I*G�U��el(���F'f���I��ʲ4o>y#���#������O#�,�v�WJ�-�%d�b�{�mG0��Ex���!�4`�|U v�9i��X��@wx�!�R&6�04�9�x��,�̉ ��Y��4���"� 4����{LD��͇i|�ߥ �TD���l~��Zy.�iKCXlNȁ�{
��r�8���6:�5���t��� �!������w�%��ڕK؍��n��dCP�e$k�Ω�P�y�Y��dP��nG|�=x��C__��N�~������T5�N�K�9Jf(d^�@�d���(Ia��d��GiH��/
h�Lq_u��*��HA=�X��<��DZL��2M��/H4MG��K��[���nX6�>p���SY1p�=�&Pc��ּ��y�Z�V��A5�x]2��{�x��@8Ԅ`�I�ǳs�x���cqm/Cr�;kh���~�x����)H�ʸ6:���oቧ����9B��G�X�[�}#��>���}����s�_���hdd��v"���19���zF�Xk(���x��w���W�L�?zO��E��9�S�W
Ջ�	�HW;��<\�-t��pW4X8)���������mB#�=cC���a���5$�W�<��(�`�v���D��"ת�B��@��$R��8goX��nC��S4�BQ 2�����xLjjd�4��)}�M����󒅿2`�V��=�!�Z�rU�E�p"�����#�Qh��X4�_����Ϗc7��bs!G�:m`I�yܘ��aC`���[����'����>�[�|�g{��_��ŝě���1-��j��ӊV�{�;1�ߏ�������D�Y.s�J�����F,���U�2t��#��΋�f�9ѝ�l���m���K�ߨ�ji��b��X�6�=����S�AGu�Cv�-EL��cP�]U��j:�f� �FÎpk�z:%�7�ؖ���������x�G������.=z�p�qp3&���h�$ǘylE㘙��B��⾁A�t�MH�bX^^D.��ͷ�"�0�6���)�#n��r�����>�N%�m���;N��j'����<����܁��v,,mblb�3�_ڀ��g��v�cm'%�x�P�D�+ڐe�IcP��-�V(ccf	s�^�P+%�٭�V�P�������g�*�Re���@>h�`����f�n'|�7MV$b	�<�� |��I���%�|n~^�Da�$=E!5��!�/sJ �3��PS|'E~�!0G����ޫ�-�D�j�uX�����n�i�5g���Eй�8k6�6��0��2q�R8�~��i��	�q��=�
�TnC�*�Nl�c3�x��E̬���ElJ�GgX
�}]ax�
L�6��dU�v�&	�W�汽C6�::4)[X
��Z�y�rC�I�T�RB��@O{��:��'���*A~l(�����0��0>'(y��hW�?:�+M�ӡڒ����&�S+�f�ߡS�D�a?���>4S�M�1��s���%�K��� 8C��F�7qe|NRk��Jꖒ���w�@[�)�������"L'А�/^���K�H�i��i&�tҫ��]��D��K�]�e=}�n9���Y0��,�kH�ʈ�s�_��ձ9l%
��-�D�`1LA<�2�@j�6�vHq��N'HWr�j��7��+���~7�>˰5�\��t��i7,�l���Ʌ,�.`jjRF�tu�n��&c<Q��iL-���psHh l��&titS��H�	򨃔��
�#�R�+��8�L
��8s��V��V���D(j�%�~3��׍�I�& ¦�����f�JE�fG2�����oLc'��4ךn:7�PS��കpx�G	���E��ҍ"K��o�R�<��k(Y�2!`�#����fI�nXx�{��	(�d�+�D�)�l
�יȼY��y�ŭ���ee{)Emc�mR�^�G�W���J
�FSi�G"��}Jօr12~?�5�m���yM�Ś�Թ:V+��(&�ǑL���Ag��G��J	:��Ւ8��:rP���$����|胿'�w�E�~�������%�(������/)���C�7�?�"�������sE�������NTR8iɼ�{l4mfC��3x��7�4���hU5aJ�&5�! ���/�j��72$�.��lP7����4�dC`��0;�[�^4Vl�4�Y*�D��\l��P,a#�Z�'��J����:�N|�#�?��b�AЈ�s�/�_��M<���p{<8q�A�nL�����/��7���O>��<��Ʈ�{=}�|�ӟ�������=�0&&&�ͧq���O>�_12t?�����o}�+Qq,$[í��.g��u�PG3ڬ54�3�p�`��0j�>/j��>&O����� ��+{ufc��0�tF#��֞@��l^%���݆���	U�6�s�r���,�l
;�Ԟ�$��1�4y]<��Ə{iT�z�	LЉR��4(i��eC A�bP���	��9*҆��}p�|��g����iL�&Pѽ��t�I���B`QQ�U�!R	��f�˷9�ɧ�����V5߽8��7��^�Z����M�NQ|sL�Hs�MG��B�ߋ��vq���+h�"�1ar�BMH�rXZ\�n���%�/� ju8\����1�p��
���������J�J<D��A$Sv�%N��#��߁�k���sO"�I���Y&
�u#%Gv�z�H�؝Q���@��n��>�[������]Sc�H�X�Q�J.�����/בL01>���5����;�o�>X���]	=��SBb����8��k7�H���ݐ<v��뫢O��w�[����M\�2���8��6q#�-�26���Mܘ^��N�@�����#�"Z-Rl�Ɏ�b�'�n��E8ɼ�b[s+X���VL��
�J�Fd� �F_�������a7��(��-����qRzȏ+����ڼZ��ΣN?d��.<s3������sc}s�ݴ|fA��;���e����@&Dj�U�]Ù��`4���@ ��?���l�4��)�:z�B88ЉވG8��V���o~�����݄��]å��YN��9qC!ǰX�o��Տ��fi�`�\v���Ai�$�{bn	Ϟ����� �llZ=mM8q`/��#8��X��`7`w���7��Wbx��$����E$�S-��Dv��4�,�*�,\�a?:���4)u�a�\��B���LO>	��k�\A�9Q\X)f�	�i��G�D���E,���n�qDc����'�B6KU��#��I3�Z�`��z�)�y)H�����M���Y)�-���W���h�]�8�mMAi�
��4#�jv�e=��5)L�t�;�G+�k��,��ͥP�{F.�^�mG�q����2}�����wMe��0�M�ܥq̮D��]p�!�S��8�<`���
�)N�x4��J�-�A\KF�����ێ�'Bs�#dD��?lt�kN}�%��m�I����L9[[�p��wc��KZ�<6��\�ݘxm��H��L�$=��+�XX��T#�����#6��t({�*Ŭ`����߆;����ఫ��\�#��#G�G����.\��	��NG�JG���t��	�Ҫ�P*�$tmfaۻ	.Z�e��烳�"*��:�i���0�6�$Es�l�X�/�O������V��؜�Ś]��p?`�b
~y̂�L�IGT���W]}���Wѿ�1�=Lj��b-S�BAM��2��kMj�9}�F�P9.B됴aUD�X"��i����1݅hy+�g#dޤxr͙{�4f�y�ei�Ѫ2���k��g���� �J���a%͌C!�+�<�lj���>�>����@gGg�=�������[1Y�<��PN>>;}�ϣ�&��7T���+Ey^)�e$׎�皲�pTM��L��F�rT����❮��ޱ ��V`��V�uI�j�t%gAǦ�ֹ���Uc��,��Q�J3FGU5���4M� �J�n(m'5�._Pi�i$��t�� ����Z��!x��g���~���%؝��u����=���B�^�?�~7�x�	|��_��R6���8���˿���0���/�����>��f��a�������W����!�@�\�>�������A/���x�&KF��n�F<4Q)fs{C�#�%b�e��ڂ��X�y�ז�\Z��iC�Z*�W������8�1�N�k0��j~�9#�BlЙ?�hЄ�W�#��	��M��H?���FѡE#kA�k��P6�V��ۅA�`��vt9	��l�]8;����M���b����ZP5�H �a/6�I���Ttu�ԑ�O=����5!��׍�<��{��د�>QӃVo EڼQtS+��[��ڊ�f	{��\�n|YP�hq뱛p�-7c'����G$����U��T�!�Q������V��</���#)�ұ�p%r�w,v8����~�]H,��쓿@tu
��3������H�z�w8��=ݰhl�lH��_~�s��ԭ��r�����˯�sA{W�x$�+�M��œ(x`�1uc7��UB�Mm�p���ر#�7��h?�0�]�.�5~"<��w�d����%"T�>t�{���L�����bl|�NOW旷���������2�ַ��=�=C�`�6��%Qk�2�<*L���8��^��@>G{C+�R;�kX��@-�K-�Z��S6��V�?9t�tZ��h�͑�]��-Ɔ��/O���Qm��y�#U����ێ�]�/</V7��y���;r���߀����Mᗊ����k�����(�Y�u&���Ex��(�5�]-������˶�,n<@se�܆�J���Wqybe�2KC�R�i�ǀ+�K�"�Y���$ٗ�,��I�U]Ǎ�U<aK�EI2�Zj�t�'���.�8Q�V�m�!�[VdJ���.^|�F'�asx_}�X��Ƃh��l1���ي�H3�ۚ�) բţ}��]�(]��?��EL-m#[�A��h��Z�¨gpdd��c�NY��\	kIܘY�v� �w�����8�pw˱�h	Zu�R� �//��&9դ�!�߈��+Ӹ4:+�Dr�lZ-!�8<��� �+|C�?Qu���"_�Å���dP'M7�!P4D�v+�$*EحUXk�me�rx?�8q�$������(kp|H��Ϗ���[�Ҭ�u�4�����P�aO)6���D�
��C�3��<5dQxlU?�_,p{ښ��(��ҝ�"I��ʘ��D`'�Ƶ�Q�|�Z�M�ݷ�C=]�K����ړ��l�yֹ�5L/l��$�J)@s���6�4�i��Ui>Ģ�T}C�e�ءh�<F�()',v���uDw��J������D^r�=>�ʖ��&a8Ծ�zĊ�����&v�)褫؝�w,����@%������!�dաiE�ҹ]v����rO�0�����L�H�`C�� �],֤�&�����M����4��NL����7�@5f�b
��I��T!�n�8�-�)L�[��I��\/.��:��Q��?e��o6��)2���5�����J�\�:�)+��鰢%B"��/����*<�І�h�!p2��-�4<�lT�%d�1��|������ކ��&�eaj�Kc���:&nL��16|$L+TS�mo�a28�e�����sr��{�}=��XR�I�cW�B�ٸol:vJ���5�����(?_5�j��h3MZcU�Kڤq&p�,�U5�}Z�Sc��!y�rOc�B@����dA���i�j�"V N�u	�$�A�>Ț����=����|��#0�-�g?����q�긤;H=A�5�������×��O�@/q��-����7���E|�k_S��l�����_`p`��?���}J�r���xum;w�#b�����Mm^�Ji��:$�F�\��t!w@&I�lJ�H�Zh�Nǝ\۫˨��� e���Uq253j�d��55�3^W��4q����=�F�RQ�:�9E����'j>%"��Qڨj�#\�8��	��n�Qa�
�����Ձ��~4��3�禗��i\Z^�B,�T����t��dt�f��iiOt4�ѥ��������G>�����/~�&|3_~f��_�֏��O�XCM�3���A*�����w�������W��6#�N~����r3�����򕋈nn��[O����*���ؗ>亠�u�钆��7���?�ո���|rh�����
ɃV�f)�)�����a���83�2�Ņ]X,E�ZI�Y�-S@jw�E�_*�%��}��.����uZeBp��E�n�<�p� �L��M��N�a6��p��(���`�4`��}����ؿP�l�/\�#�<"	%	����E:>>*���Ȱxs��74�w��]��f���1Vע��?�x�$��wX����Ģ�k�����ٱ��D��<u
���%��8%��l�jY�U$W6�6;�Rb(1��Թ�2�Pč�,&8�'�BgA��$�T!�\�,�fW^*�j� �)^cC�s�L<?旗��s3f3P%�&>�
��P/5��tܐ1��H��kx�e6�$l�O�k�y� 2�4�.�4tЉ��l��A��F�I�Pډ��:�勸1�&����E���p�t��b3tb_;F:�b#�i�$Hk��@��.m���l�V�!pU�\]���ώ��q�� �j�����t�1�ڎ��]���u�άBMg
�� �#�LU(����>t���n;��Y8݁B݊�DO�xI��d��C�dI�W3�i���'�N�H�I�K�6:���eѲ�Wh-:�����h�p����*5䎲�v�b����95/�ps�1<q3+QT,N9���M$�5��f�+�������y�,5�\�Ն�63+1L/mbq#�T���8�P<h1l��hrW�p��pZ��u�e���!�I~l��3��½�llϽt�O�uc���л�eb1��4�\�C6<��lT����Z�	�����]jz�B[�R"�R�F���E"�UD�el��������
���{��ގV�%gZ6iXe��*�G�t��\vqr�46+�m;tsх���*
���Ng����b�#�w��[nB_O@lS���=��R|�������z��)�l'�M��F�[�t��~���as�aw��f<��c�#]:*�3g�K��<�����80B5���b�g�*�\�#S�!��blnc3+�g�B�����#�HD,�/�8U�o�G���'� �����8�~������3E�f�n"Ȧ�P@��������6iD�qHM�UEI���B̀9Qc���L�M�	b��b�T��6�U��Ё��� ���t��J
�K/����:|?v��J��d��HgT*-�&��?�BS����~�=����]�^�4]�.]���
����Y����J��'��oUy�,5v�gΉ�餣��b���'I��(��s*�#��aeuKkt+ʡ�hE��t��� R�x�%�J\�j"��������)�kf��CuNYZӪ�SE��_�T�r	o@����&D9Ԫ����!���)6�k��i�������AW4 ����'�����.^E2��Ɠ�5Ҍ��y|����P�+_���|�n�;�/���q��!|�K_¿��6��)=y_�c��������1q��vڢ�V����ƙ#�WQ�X��N?��<R{i�L��Ep�,	�Lx��'i7���\n�=�0ܚ���ui6뜢p��^(�j��fJ:�F�����������I���׉�T�?� ��/�Pu@C��1�f��4l,�1(�B��Z g�z8���^Dat�a���G/\�������W��U�vN88��c���f�8iܕ,J���]'�|�ѿX㕆    IDAT���V5uǏ.�����g���)y��m(Y-�ۈ�%%?�^��Z~Álz�X����D���Gុ����+K˸�����$؇��<����T=�����[���~��Vw7O�x�s,Hq7�����GE	n��hqZ�4uӣ��:�vam��bo(�B��U8�DZ���Q.fqhd���qӁ!��yLN�!���L!�������'G-�.*��T������t� �����b5������g?}��կ$ ����-S 8@ǿ׮]���S����U��]xǻ~�]}x���pcf�`�ݏ����܋�����,�5�����'ʝtZB�(��9}e�x�*Z�l�0�kHml#�4���&jE�!`~CVh4�M��(�Ħa��͍O��PNJ%*�)?�+�Ft��+b���@���p���7������Ej��T\��h[�����%�!m�p��8��A�L�@н���~�^�5�ֈ�0B���#���_�?�V%�f�5���צ�x��_cv9
�p#��b�紆��r~�a{��oOA/زh(�bC�.U���Չ%̬f��KV��k���f�PVn=2�=s���P�L=�l�2BY�6��b�e�&�����æ�,�����=G���fw���h���R^l
Oi��ӓ���Zނf�
M�W���R�p�� <vH�͵H����^x�*��9��؈�j�bVɧ%���3�HS�pP>�V!u�ߋ�5qz`*3u��-`#����.*5�O{�ˀ�Z�,���49`��E�+;�`7[���2�O3�/SНFg���8)U��9�%qb:����~t���Պ(�7Ft�M/{&�����KX�eP�8��F���4t�j䨨S�dD<װ��T2f�ci��,e�u�����)���C&.���τz�X��*�$�Y����YL�O������N쉰P��Vd�f�EA�j`�̮��\�����
�w�H�JpR���O틙�M
F��fPͧ�����'�o�v�(�\��ܦ�+�f���UL/mIA*�Q9�Ȥ�cA2ʞ�JڌM��L.&��JwC�5h0QD)CG��y�=�0e��t|K�dyH}~Tk���u\����9q�bv�R�!�} (�2a;'��q2�v�3b�K���ߤ���5����|=���t�p7��r^i�̟e����6��q���#?\4h�� �,�ޤ�Q%Vf����)n;kWixh�)�V�ü:�1���cm���f��1�*��	�>����8�Z.�b:-|mK�*�!B���8��wߋ�ϛ�o_JE�qJ�US�*��L�kO��<Hh��P����W���'�'?'��j��Ns��3��rQ���R�MyՂ��(�~�9<��_c;���*wFN��h��k�Y1r�*��f� �#�$�: �e��J&�#J��ƃ,
[�3W-׃I��A}������&|���9a"�q�P�J�BA7�t�����!�P>4�8w�e|�1��"{O�Z���ui�~�wކO|�c21x衇��g#�����7���$G��������~]�7>[��~>�'��޽���W��Ǐ�~�&]�`�
�{:�޷�	LBڝ��+EĮ#d�Ò/�V$�a�M-�]�A�OѾ�%��1	$����B�x\�Qg�"\�oj�_�+�g��V�Z��2<L�v���2Ǆ� �	���Ȓ�� C�Y*l�${��↽*ݷd��u�;��R�ӭ��Bٰ"л��6��"�ׇ���_��O_���|i݁Dł����BɪK�	�#�MNK̆@�VQ%�]L��s��O��/>��oUC��K[��������܇�@+���퉬)g��t��%5��9�� �#���؁�����𝇿���9���o�]����i;��_cq0Ά�ŁsW�񝟞�����U��Ƀ'\ݐ	A]����O�^��V?v7�1;qk�㨥��������ZXD߬��m
�r؅����+���p Kk�x��XY]���D�[��˘��~�+X]��Pd�x�,=�Q�����D	�s��fp��9�'�h��>��X�@?y򸈏�6@~���n��4�tϽ�[X�<����t#����؊����>�مuqL9|�F�Sy$���p�K�kkHAme��K:��n��2�m��΢��!�T�q:���h�T����D*�8���R�����(7c�%}I�>>Pr��a![`�f}�o�{?��2�0'q����ϗ��/6f�Xc�ȵ h?��|�t^c��?��!S�g����p���O�HW�#䴢�Ń�Mhy% �16,.b�*�7�=?���<�͝(�X�1�Ԟ��I�����v<�Z^R �q�.D�z;�ù�70�D1��LJ9%|N]�GO�<�����">�tk`�U(հ��J͕�u$�5�K�,'G�.8BZ�QTO=��^]�.�vrma�P�X��ᔰ���D���3˘Y�#]Ԡ^u��ޗ3�Z����0��袡Id<��[;i\�6����%#C��_'hK�RNp�݂H��}=�ӥ2*YA���ށxU�R4�W�永�@"S�]��5����ky��r*y:;Zdr �Rp�*�Uo���x� ���p�°'��Ws�9���ΰ�N@W$((!7tRlt��L	�N�0|7W���s`�B�L���|v� k�X��:-�Pʧa��?���C�D��1���~�P�2ټh���QḼ`|f
��$::[q��C��B�n�VIK"��j�ՠ���f��__��/\DZ��~T�6�Dq�� B�ڐ��H��\^CC�Ê�8<�%�"m:s�����ƕ9��i�ZG��u_��l��U���h�7]�8��	��r"�L��as�a� [GG�o}�)�4b~�A�`B!/�gn�v��dY4$g/�a7WS9jq�<p��϶)��,�Mߜ*�}l� AĽ�@�����#�M�l"���6��@MT�*�Hi*����������	 �҂$� +�
�y�8S�����uռ�!P?�a����!�2d�'x+�ɮ���ͦ<㤔�x�Υ�.J�������?�t$��ӥ���߉�}�hk�K�@�=9�<ӕY�o>Ol�mB�20'W�PJd��x��S {�*ֈ6��HR��Z��D��^	�g�
�;����=�09Y ]��y,"y���_�lB î�f���w�w��V�v�&��T�g�M�q2��ƫqޑ���
��MGcm����4����Ib6S�%^� CNI������!4(^�n [.���x��"��I A�K�.�X(�ԩSx�����!��O~(@���Ɖ�O���CϞ^|��ÿ����w�)�p�uw�����>���9|�arz�\A�Hs��to���mV��L��4�Ztz&�Ӗ|Nr�+e�6���j��ކ��[ص:�6.�u(�3rVqz@	s.x�����RVV��	����f5%��$�f�ƎBB��Ui��tZA�5A&�R6�fSF�U�7j��T���%���	ks3����<4��˃+K[�����E����V_3
�U�u�K��=T�觨�e�q��v��s��G����?�[�|�����o}mv#q�'�{ $�,�t�kL��x:=�keAuY@��u��-G�7�?��c}mw��N�r���!:��NrS5i�_�Q��Vg�:�u��Xl���'c� �7\�vK�
�����q�\��bb�Զ$��,8�mxN��Hʩ8�~�gn;����N<4�xb3���*^������"l}m�|^OH��D*�d:���i:8�e3�hPPu�����+X_ߔ��)5##C8xhmA����Ii<����#�܆��y/_Gk�^���nkN|��O�W/\@Mw�gϠ4	8ϕ�+�Q���ؐU�8mJ��p;�}ri�U�$�7�>;�r**(�P��3k�lŝYPz6
�'/��pM�ł����#��(�R6p�,4�Ҵ�q���ɂ�3��w?p��WV��j��@��!��b�!��k��X�MC�j�������B��W��Xԑ/f�s[%Dlog3��=�tx�M@�����`']�j4���Mcqm��XA��ڑy�r����12؅&�Ulp��+�t�܌e��+c�^J���R	���X�ED�n������<<H�R|s�N�~rg��Y\^\��N�,���ȁ5�ቨ[��D��;�t�����C{��2�|j�y��Hayc�Ӌ�Y�F�b���*"D����8yx?�"!xi&������D���$m��*�u8�)���˹Z��a��`x��Mn�(��%����6vp}v�+Q��5XXR�I�F�"J)��铤^�׀æheb\�)AM��z�L`bz��怲Ŭq_S��]g\`��X�lǑ�>�%��Yy��=�h�0�:6���%��^���CRl�aP��Z��&E%��U�x��$3�ɮ����G�(�ZHȄ��B�n�L�R���Ņ��<^�>���9q���4�v����8��.+��,z6�Sh	5z��NIs~���y�22e�l���<Z�卜:Q|,.PE&ǔ��e�4���(.�:�sb7\�Cr2�K!�Ս�ՐÙf���M����<�ץ���}px��Mdd߭�֐��|W}�!��t����F��LZ��,��N��.���kS���B���?	�X�ˁ|A�)T��M34)C�w���?��Q�Wh�IR�&��`����q tN=���*�	T��B�mR�(�������-g�#N@�
�bE}i��`b62;%�B��w;���4b��vv�uy��g������t�).�4J�4G04\���I�/�U��-�����{���،��@]���8%�I�;�il
��C�Ah"|6%����2t�ө��Ԑ)���*�A������B�������#��M�����|��QW?KC(�(�8vt��ԃ���M��)�$�*i^Ho�{4�i��F���{5�2�Vnz԰�ɛo�#�'�'k�H�f�Jn]�(�t
K+�H%3X67������2R��ؚ��/뉍��䤸%B{W�����5\}��ͧ��ۍ�G��#Ҏh4�������fg�J�1��z���M���mkkׯ#:=�*S���3Z���nB�	�-�X`��+��А���"vE���J�PR#)�e%����<!��gE96��ƓBa	��������7Y$܏9!P?Z�$%Y�����I��S���Uؐqbn�wO�FB�`lu�����-"g� ���	�d� ]��hs��� �h�x�{+!��45�}�:�sw�z����O�V5��ԯ���?�[۹ʭVw�K%�L����:��e졂�*r�݆!�z1�3��ě�p^|�E�<p {��"�P�rN�$؜t�HƎWƢx��g1���v8|-���K�&`"��T�.����||��W�]��q8�T���0S�x:#�͆�Ca���7�o}�.��.n�N���+p{t��KwLG!���N/�B-�y��pƒ)\�zW�^��N��`�'����șT� ����G$��������������҉�=�_���r�@=���-|��?��nvw�{�o�F���I�2�jN����M�U]���J*���l�Ϣ�	a*6����*gI {
��P�X�s�B�"J0�࡭d;R���Do�.�?}oyϻD���C�.�!�07~D�v�ߏ�� ��Ϧ6]���!��	���!�D��'���j�=�
iq��׉{;�t�C>�]m6,`8!���2!�2���h��.T*TA�1FE�������� �7���Q��dS�X�"H^���s/^��|n_+<D��y�V��8��u�8�{{#"�#�;�)��2&6v���I,�F�����KN݁V)	��7ľ��Z=�j����g��C��y�$V7��ϖQ�y��"�FJ �S���8rp��1���#��cay�&f��̣��D�*����Rϒ�%�Imi��	M~�n�"�3�;hyL���\ܐ@>�;�1iv�P��4:���i.����r�ŔnКӅ�TW��qy|ۻXlXlnE�euK�b
�\�=-��u'��ύ�vFP{N�2���]����]���4N6gP���b�����k��2�J��[��BnY5�YY5,�8M����C��P�'`�I��0�?�~�����^�2���(Ju��'e�rbd �OD$d�d�T-���H�s���0��Q��g��s�>9W���չ[�j����`K6� ��af���,00s����{��� <���`��IN�,Y9��
-u��r����<���e���./���������{��IҾ�=<��e<w����䀸�}v�v@ �o�3����v��za��w��E���	�"��3�O1����K�?� ��c2j`�!�p8�N�-������/=��OPÌӧ.bu5�f�&����D�����A�~�L��!`�.'~^_ =w�bS9t9�z#����P8,'50���C��4��Ʊ�+�/m����S�8��&�v0"���g�︡��hQo�s&�W�Ҵ����Q�kh��*P����F�4g[v�g�6�ݬG6����v۸�Ps���Obm}E�3��t���V��^��v��>��݀������8pp>����n�P��~��I� �u��Jl�a�D���E��y�b�F�6t���	ٰ�h �kȔ\�����s�o�<��2=��W�ß�"f���`E�2Ma1�{�Ɣ3H~�f���o;�����[��فs�I���W�&�P#;+�����{40u�&����}B����H�8v�#i)���~al���T��/j-�l;0����ќ��L;6uRu����2(�Ij�Z���'5�R�����������_�/���8��Ѓ�51�N�w��P�y�y�~��X m�B�V�&�t�#��te�J�X�-���b0יV�����G{8?��x�����ә�k� +D.��x�ɪ�bb�"��P��0�E���@MNj��)�`}ɫA���5>R�c���"�{bӻ��u������=�".�7�I���8��#������%��a6=��,�Z��\4���ӭ��sd�o��������Ϟ|r������s߼������jx���::����<�T�I��B4�0�m\�/<�Ks3X_�ʫ?Ob���Vø.�\�Sk1����[����#/��\m�����+E�G�4�hUj�ynO>&�z[�*�����+e��KOc���@�����06��;�P0�D,�V��;n;�_��q��.�庶���_~�/��Б1�۷����6����z@��u�L2�+��SO�@��䤦?\�[�N��8���O�B�V�D����X,���\�<'����)M+0��p����-���ć`���#�:�\}4�mM��w󡡘'�����H�/���f�:3�vfID�.Ć���c	IA���f��� pG�ſ6����,�-�(�;	���c������R�?Z�	ǆ�5����r�q��!pE�.d�kop�(��Z�����z;kU"@�ნKV�ty�<m�ݶG�Ė���qr�����a�E� U�ӗ��Z@�o�c�4�"=�Kk�^AOcCQ��9���iD�}Yű)�)F�k��ŕ�%<��I�,�T��C�Ĵ�\Й��ȴ.=��G`��-Z@�I��T��\�]^�~��r+W3���u�#1����`L9 ;0�u� �mK|\��ౢ(Vk8s�2�:}�����-��tX1�׬bl0���7�vZ�l��3�.cfq]�7���#Y-rzi(�b��A,�H*�S���F,�}%{�R���~u���^?�s3Kz��4�A�)�*��Ɔ�طg;vL�(�V+H�L3+A����R���0��C��@���s#��G7��\lH�z�1=G%W�¨Rkb�PW0}�O��E��/��%*?+�!$�p�    IDAT͆@�W�kClH54�|U��d�L��T!Kw�z�Gѭg���[��X4���Jm�����3Q�vᥕc�<�n߂����D�n:� 
Q�����Z/��ř�%Ѽ���iLUk z�C����J;�\�FA���{�kkޞ��d�@�ւ��1.������E̯�s	Ei��C�CD�������f�%��HЇ��al�:�x:�Fx���xaV�%����9�+a�DJ�t[��!h�kBؔ5:���x�7q����!`SI"�P�N�5� �'n
�R3g_��v
�,�A_���Hn�9�E�=��D[�F��G���I�uQfA�ZJ��j}�����r�>Â�_tk�L��_�4>�׵ڰ�D�?�T,�����E���rHz2�{DHv��h��hW���xF����J���vރɉ�����S�L��j��[a�tj3p��d �=��t�_s�HC%�ۧ��X��y��J�M���X�� �{��+�q�����w�����-O#��IĊ������P�R�b|�����{�혞Jh��}Go"/�NK`LG!�N��.c1I��s�C���Kp�S�I6u�v�1�Q�+̉�!�	ʫ"�J!�4:���xF�}'�/�ZJ�ak3x&��?��Ԁ1������Em6�!O>����G������!ٷ�VŅE��\9�:ξ�
�kX��W�hW�
u��H�FB��Q�Bc���}��ͨ^.�Q.�����@kv�wDH���0�O�?ۮ���p�����؈��2�d��FB�<���tI�	E�Ə����\p�H��#22�ԶiDw��Cxkq�<�"�8��V�Ӹ�λE"Z;��G��B�DZ�����n_�~}W-/�{{��Vssw���G��o�x��������S{#��?�kš��@�E�ih���	�C	�p3����U�³^ɨ_;)�/]�5����`bH�"�==���ҵ���KU�÷^ƙ��4����05z�
ʖ�"�mvC@���c�h
;�GQX�����:.�xE�!�C����g�dC�D�ʥ5$�!��}������b��1=o�����㨕˸���|�&ټɝ���imH�P�zI�����*���66"S�;DbwJ>���H!�t"�?R�:��(�#����y.�?���x�Y��	"cHn�)/��P���+�A�a�l"�0"���/n
���=�T�X�p˗/����)�Nd�l�S(O��/��&gq&�*�3�s�����o&�ȶ�c�����~��Ҏ�{ 6���Q|���Ɖ���M6l9:�q،ln G��tNSO9�$��ݫK���-Ca���TxK;+�Zۍ��x��斳h�9�6��F�f�6[z�]ۇ1�#���i��':Pot�����ˋx��re�X��L�d�`&��F~_��'��&�%f�a�֐���D�Y\er�,��7W�+y��j�&Ǳ��c���x���Xoci�.z��Wf�/W%���:����&g�nI�=zxұ :�:���G����WpavA�
���a@}6���Ω$�������Ug$C,��A.-���
R}N��E��E(�Ԕ����v�~��s��߳�i�h3G�L^�LCmt�-50�����e����hv�&U�V�9��d؏�Q�MOP�ܓ�'�28+mTi�:��������欓bh�8e�k(���y��+����'����n�M)��x����~GN�!��k�`���s�y�v�
N_����|p"�>�n�������5:� :=?�W�8q�
^>5�R�����'�����²T)�T���hY�:#���[0=���T3
�^����t\xC���St��pˣb��Dg ݎ�C��L�chh}��kE�__�t�VW�L#���jd (jގ�q��p���P��k1�ǟ?�+�Y�cC�y�Fh4�\��q�q��5Q�>&d�F��nsa�4	N���8wh(Π�A�d�i�~;C�k��Jw�!`q+'�m�k�������L�{�QbgO41<FOf6J�H9�-l::D�A	�k�2�y�)ds�GtRx M>�	#=�RF�J)ò�	u�C�v�L|t�|n�g��i�j�jقF�P���$����1�y-��f�b��q(9B�]����<][�6�,��������g:|&[���38�(���9��x���v�>T��m��n������C�ݍ#��KP]�TЪ�Œ ����ءrBM[_0ͥfҮ�\�tXG���&^c;J�D:�I!kJ���XM��md29Q��ȼs�.�޽Cף'3�>��6¡ F��߀�,��A��S�z�Á.B�����i���~5��k�S0�g�{O<����n����Pb����
UW��<W��0���UTYu:�z���14����B��A-�����F��Ok.��o�usYt�#���Oq~��R./t҇IՒ��X�6�-�'��An�L�G�o�E\[�ZSk��Q�_��LDy�������[�"�SHON"26���R��7���ko����x�g���_G��ħ��Kx���(�=�F���Ā���v��^�Z�����&��w��[���>��M���	T�g����g�z����'�x8K����?�ƽ����MA�DS�dd�i�߆����S:3�P�z���,f��h2�����D�-&h�U��ZƗ�y�g�hb@7L�c�)EŜ
�v���@�݂7�Ŷ�lIE�*dq���p�سX�9��]|��fA��@��^A̤�Ѓ�XZ���Q����z�~��4��fV�E[Q4'^��x��9j^?je�E����ӧ�o}�/_���68p��c�a��#ڐN3|���O6yq�]& ���C�|����?�,�כ�&���I ��@<9�������A�zN*Z�"�R�����1��M̝9��gO��@M W����pP ��n�&�B_��	`�����k���P��?�1_Q�8x0q�ux�?�P,�"T�n�}#��{'�٣��h�9��N�b{�4����C���*]�gC�5�MatdÃIAÞ^M����� ���!��'ܞ Z=�ke,,�Eʗ����Z׃ɔ�ϡD[�bt�"�,OS�x�9ג��enA�J�f�pqv	kk%���=m���z�x0�19>���wb��V}@�ҒƁ��?�Z9��&G���]^s؉H�hĤo�aȋ�Uf���N_�����le�I����x���.RQ�pp7�m�E*7� \��F˫���C��u�ɳ}r�� �=Z�����I#�617&�RL�9�����`����,�Փ�E��Y��A�����Vp7ѪD�ڹ}vMbd(����c&\�I��\�w��p��P7Q攳�E��>�Ncz�(vNcb0��.,T�-��}t���WKu	��Vr(䉦�Thp��|]��^��% �r��ܰ�4�/%ɵr�@o�� n;�.N�˴S�$�Ax!^�]�s��ą�EcI�����Q�d2��n=�]�)��eT��`a艠��cvn�^;�7/�#���V�9�4n)���FE��pc(�R�r������w�q�M�)!V
��ƻ��Z����\�ɳ�(�u��`�;-DCA�S1��-u8G�!�1�N`p0���|��ӧgx�������&�b'�o!���C�qp�V9��+U��-x��]k���g�)�J�*	�G��n�|b;�p�m���V�� �1�Po����wc߱o��v�$�	p�=c-���h��wRm7��&���=�������~�~���c��4J�n�7��D<���4���}�i��Y�~�Ay[t��E��6�P��AD͚����.�PXBmmѨe�,�C�ȅ�ڲ]�((fdk�L�e�A������m~��E���5��ϔ��_+d�tQ稤[��-y�MN�}A$�i���j�dR)�lʤ�Y����GċF�h��� 또衵bYg	�$�$�g����t�ph�I�u6��|�{�R�'v��s�PX��;�T�����1a���t##CI#����_��v���������'��c�=�3o߾=��۱cz�\�?�8.���F��ӻ�qǝw�=q��9d2Y�KU\��E�VŖ-cL&ЪT�_\���<<�&��>�Z��ɠ��(g��V+H�����81>$�x~m��e�YQ�R��RI$�Q�Q��+�g�ٲ�>bXl<��ˣ^%��\7R���w���&S�~� l0��r���Ve�D\%5�b��޶���Y�LF`KDeF��(�5}n)��ky�[-୙E\-V0�g/~�����^Ժ������سX�4P�yP�V�%V�P��R@]���>"4�,e������������?}868t��?���3�a>�����FQ]M�^����΀��o,����)0�k�P�e�T��\�U����n/^=���������*��7҄����{]n�|6e��)�C~�-�
+8��8�Ƌ���ş��1�>'Ђ��Pb!᣺
��;�q�������C�pÑ��y#/���X$d
-{b�iD�\��N�_���믿��~�{�K޶���	��Ƌ��U>X�'�L��1�	.^:1�Z\]Z��/-��g^ų�N�4��!=�ՖO�!�?nh
n7Ztm�[9����F�~M�Zj���`��\>�&�ͨ!ཥ{�l��^�>�l��#�3��J�{0��������Z�X@��w��O�
 ��d��aG$H�n���M����؎�̵�&�rz_��Ά�p���o����mc�|�ۜ��0�"匱)hfL���s�Q�[JÅ�\+��lh����[��2�S[0�"u��b�U��Հ�G��	�aC����	t��8��)h��@�͉�s�Ӆ��J%��3"w�ϗ��S��i	�D��X�R��֟d�A۶�#��ϭ7 ,�v��W$$�0�!/�tJɎ���D�HX�!��XtO��`yh�i����QC�аfe�@V[��_��ª��VH0~~�͑��ST[F$l�W3��h��M\^Z�[�g������LD�i��裎V���4���q��>�t,��DD� ZO��������ui~^�%��R$cH���u�Ɩ�ۖa�Q�2��r�X��q���2f��(0��O.���{���`�f�7V�b�Ԅx�\Ԉ���8�E�ܰ
�^?-�P�V��C��'�r8}�*�:�2�҃H��B㪹$=-�{�a<t�~ԫ*z=_��Wf�����TI���B�6�ۑ#��f��F�"�d<"�F���Pԋw�u��"ȩ0�9��Q����N_�Õ�����^��,ko!�A<yŹ^���H���D���\Z]��W�`-���X(�@����*�%��]�:OO��e�gE�\��m���)/���+�:�V͞[�!�&Ҷ8E��	�r��"�LeM��Ї��i
�}�G�q���_��ۺ��h�ӌ�$�{��蝜�o�{���� 9e��|���ޝ�B`S07^��?e�L��f�0��8
�,^~�%Y�Fcaqۙ���9A�P0�����?�
G��y0�Qk���A�h�`��Y)E�t���u@ɱ����9�O�u)@m���=ƵK�R��{��f� �<��U��d���L�_T�P��k6�D[R��]��i�����ф��H��db�!��-J�}r�e����G���ߩ�P��*cSʟw� ���1br��I��>��q#j�AP��x��Z�� ҵ�]o�����_���|���_}�/T���a<��;�K���J~����~�RQ�mw܊���oK���>�'�|Z{q&W�`V�N����D}&��H������z�/�y��~���	=$�5�_}�6*+k�-]ՠ#�em�p:�8'����Dq�J��j�2�N��D�\A�Rٸf\��R�>pݐ�f�:6�2����y,Fl.�*��+h��#6�T#�aJ4�p2	w$��7�+�".�q~%��L�H�o������=۰���׾���ԋ�t=(�,�Tj���rh�#���Y�a�y�f~��>�����'�w�����'��ԁ���?��@"q讻ߦM��z�^nBl�ItQ'���� �
���$��Pz �N�W3�}�.��y-rf]]%�z��4�hy�8v*���.\m�g�L	~e��9Tp���5�v���������dv(�^%�%�qh��[@�.q�oP�����ӂaC���-�����D�[�p���p���e�N�16:��dRi�T�+y��f�+g�Bh.�)E�/��j��}�~\�����(�,�����0�������|���Ɨ�>.�f��$�M 9�Go��u$t�S(G��b�g�'�*�맩�ϭ�>NK9���j.��P�jg�3�6S`��������m�����96F�AKZ664�Y7aV
�zmxRQ��F��=�Z���w����l��L�K��	!Dȃդ�f�Nt ~����g
�;>��JEל4��;�c�/�5z�W	���Zp�i�Ǣ���69�a��-��XY+`��Uܲ�طk��\W���c��%��ioIj�������)����%��0�l��6}�e�kփ��Us�uQ�����(�L�@<A��{��H�RC���M[_=ģ1]C¥�JK�P+@�M����̕�87��r�I�9!���=�G�H&��twL�3%�@�S���g[]
y��E�b�]��uhW��(�Z��v��F3/�Ͼ�;096��D�<��.�-bna�
� |� �tQbz�b����TZr�aS��ae#)��:��'�6�	���ԑ3S�RG ��@Tk�K
 �Lϔղ	"�P�t�.�����X`�V��l����oB|�wnv�b�%�0�֕v�F���6Q6p�z���F8�g�wO��eH�g���#�k����![i"�Ji��*g��p��}x�}7�R)�֨�����%���v��?�N����m���F��T��mY����ØJ��7ioK��ۥ!��zA��:��.�\����*�u1��Y��#a�¤K@���p\�[ę��X[���F��'04��֩A,̝��oz���F�����Z&�'1���O*��֧��!�A�
I�%�����9��3�yS���Q������	�)6-�]���;�e���4D�6֎��d7�_VS��&�tc�#��L����@���oTJ��H�Q���ꫯ��N���U=�S8�,�N��@9�ux6���b���Q�ca�8]�_D.W��m ���D��B96=ܧX�K{�1�K� [StҕE�2�q�N��r��{�5E���t��vP�Yu�1���Rp�a�K_�Q�@*����DC*��k��>K�a��]dz��k�g�3�rG��P�t�-��)�L��)j��p��!��dd�9��ٷ*n�): QN�k���?���×���_�;�m��A|�#����ӟ�|�_Ԛ����7�!�s�_���x���f��y���r!߿�h!��b<��x$��hq�;�-x:R*��L�RC�c���^��c��$,ҟ�Σ�YA�Z���Ha�f+��h'�n�R)��=���B�B��d����e@��@=�=�j�z���Q6����<Ȧ�B0ArhHZ�e!����,)"XA�X�vG��bǍ��6.�P�������w"0���������K_}�fVPuQ�%"�}���-RBe�n�M��iVμ�mw|���ÿ}�Ǫ!��o<s�>������C����g��`����=��6�Pf߃H,��h�jc�~�}���m�x���a��
n��NL�ڃj��D�N*MX����1�y�u|��Oaf�Wxnz���Fٷ�6/��yhq.N=8��|�I�$3��ma��[���q�� U�-M�h�����%�������?���j
c[�1<���p
{�Mc��-H�⽱�S�+�I�-S&�u�a�z�5|�������;��7�`�mX��P47uN.����6��'��4X    IDATTZ(W��Ǟ���gp�r#<�c�7`xb��c9��
��X��}��-&�Rsa͘���k�أ�����ʅ,�;���f�I��^C�Q�e�)�v<0�va'q7��'0�&8�um���ڦ�=�ƽ�y7�!�4|����
؜Iq_�Zl�w�ɺM`��6�mذճ5LT��j: m��ٜ������@��͇�`d�!��,�C�IwO�:���]�Ut{�Z-+�b��ٙ��/jJ��I뱡!��E��GC���{M<�A���IAy:��(�\XX�ayuM�'�� &@ٿ(��n|xiy��:��ϩU:����qL� �-R-�p��QA�h�������OJJ�RM:���dJ��^�ciPS�\,J���nI�s�v�@*a��]6�nS�(n�B�.Ԥ��u,g
�_\G&_TC�X�	Q"
��秸�S�����7>2���&�J�f��x�Ξ��B8�'/֍�/**���DpP���G
(,H�0>6��-CH����d�n�g�C����
����tx
�u�U���U�E�t�r���ǩ3qu5��7��N�7�Y����gv&�δ���J�f�´�9��ZJ�C�����A�|dF�Ӂ�8�s�gq��<.���"�����γ� ��3���8�~�!�E8E�����Wp��U\],��
ˉ�SNY"�a��R���-Q��D�~9ME"^��:��T��@݀�.�\����f��9������z��^D!�K���30;��z��'����
Z�>�� �I�x�>��X^�E�	���m)Q8N}����X"�/-�����Zn?����p�%��@���8zg�QaB������k��k�nNc���O�^���%;��h�F#a#��k� �k��db�V�|��׆��C51�C��c�'H�B��(J�eC�u�8J�"�?�\!o���4j�>��B��6��\�\}�EQ>ʭ�'�~v�[�m�ԶI�o���ŲN�9Q7<y��d$�@ ��6���B��dêtk�F�^0I�ױ�|Ea�	�s�x�ו�?��Dar�;�l�'p�����m�>s����fq2N:#�1���|���&bFiNb
S�Ƙ��T`~��:�����h�,W��s���Z�����E�UD*��J�v���!��+��:4*i�P̮�C�����������#_{DV�|��r~�~S��������zDZ�R����}>���\�̧�Ǐ���pS�I�VU��#�c�\�>?��I�'�HG��z�f)��ׅ^��z� 7�+�n�h������ j�
k+X[�*w!�p�5��azjB��B�R�rE�/��#��A�׋�*-ݙ��4�����Õ3�[���	��a�щ\DХM�!�@�D�݇;D�ӗ���!G���r����?��]���ƣ�L������b_}�	{��V�
&�7�h�k�e�Yc�b��tZ�YJ�f��{�~�G��{���UC�'�z���٧����u��qT�}UJ����?�Dr&�I��L
L-�e�I�߾�'qh�.��O���9:|7�t�����v��{GѴ�'^Z�_~�	\�zJm��1�������B����4
�YI�`sb�-�+���P �R��9��y,�K	�^R��E���⮹i�c,4B:��ō�E��Ci$RQ'059������G02�@�]f��"u��F<`n��]8�8z��޳S�~���sgRc��B7T×��A�_;�?����ﾈ��^����SX��Piӥ)��,���/�M�t����&0��Jh�藩{������Ϡ8;��zP�0��ף�6U0,�9qv@(�Y	��&��ZC`����٥�u���;[����<D_4���jL3p�!��p?g�ƢcA�����h�bY�1�����D�|(��,���EG�@79(���g�ɮ
꥾�ORAX���nB1�-R �r�,�j:Rq���<jx~��O�A�TR�p?�K%mb�r����=�g!&������ghQ�I�:m;q��A�%È�L�'T>+&`��2�9c��'<�+U�|�es(U�H���ġk�6nN����i��&��`�t2�F��:q�>D�1��1��b���]͉�_op��7<��_p�iA��p��FØ���萊h'�:�����[Q�Q�{��5L��:t�`�g� C��~K�
x�X®�ea�	�I�Ɔ���8�˩�@���.\ҫ�E��fQ��� �Ei*������|��A��M��Xtj!T��LC���gq�ڔ���p7^��'R���^�3%�y�D�ي+�RO�?�h��,��16ǭ�^�T�..,��(�8u�<�\YB�B���\�L1y�z�9)��:��w߾HDج呈�1��b(`Ic�s�U���x.W�*$t�����r�����<2�ZI�,n|�F�!������
�z�����o�#=91��w�+�V��i5�s�U�Z3D}��P�UW�֔��7��4��L�,ę_D&�Y%2dx"�lr��^dL���iL��â��Ź��q����Z8E���� ��Ҵ+!��6��ͦ�*;��S�;(���M�a��|]5�N�gGtFx]��݅����g�U�Z�s���EMq��H�(ѭ7E�3	�&o��e��Bj0.�7�˗/��P�0��nCNF�줍y��*�;J��--�I��i�p3.�.�5����I����z8��#�/���
`�z	I�١bB8��^Ϥ�6�H�����.6l�ȳo�yZ��~t[]9�M��_�Qw(�L�)�.Rgi�KD����lv�D]x��SC�� ��Pc��YB�,B�y
��w5��(��p�������m�x�|�S��׿�u�c<�n��V|����(C���G���R}����w�w~��5t���k����WDVI�k)�Y
���m��X���H�����tЏ0�z-�uk��'�k�5�rںe�۶b � y�H��
��<��>/&G��$��QN'9�'p������W�S�T6�=���?�=�I-��C Zw0��
G��3�{d;�P\v�j0��pG��R��@�l�ky�Ã�>����!�c5ˍ���x��sx�/���%d+��J;��
�P��n��e`M���1<��{��_��_��B��������|��j�����$\ͺ�Xg�8�l.j�����0ȉԶQ|�����x�����k���u���{PkU�jW�e")_+���{~���R
":8-�C�f
M.�_����X�p.v��,9ODC�3X��@iu/?�.�A�Yj%mJdC�!�i�0���Z�ŉ��<��z4 T��p:���Sسs+F����4��)5S�z�����(泘ޱL:4�M����4��+�9��:�%GvN]�����{x���HN�ǎ�c��ë�/��"�L�Y� �1K���(q��b�K���8�Ǵ���+X=w��EX�ڍ��T>�?ѡ�O�k�7wX��.C܊�!�x�Lk�UCJ�����)��=t�Q��އ����[W���Z�3��1�99͞�{�J�����_�4���}l���7'�6��"̞�qs�&�k�099��"�� �]��`�
i�Oz�H���V�XK�]ȞF�ӱ�#	��yH%+�~�F�h����z��f۫D_�!Y��;� �5[X̓Q0�)�X�󳓊�1�L���DCj��[(R�Ԑ�Z~5[h�rexش�5���;B,M�!�.�?�#�`��?/Ұ�$���������Xi [�
�eȕ,Y�$k6�r�Ն�괴��[b1�R�7�$��2(���ax=!�xh+,�e�}�:�d%~1�9�o�ը�ݬ!��ar��G�h�5��Z�x͖[�j�Y:q��M9Da���X[����s��]P�����Q;���r
5�n���Y�*$m����.7�6יT�:�e���Ά �a��V��1�T�6����N�>���"���珙�/��9u�6d���ƽ{����� �	�_(��c�c~n>?Ù"�B�Y��Ec��^$��_(�š��e��DZ��LqN��6|�9A�됷��!V��y�zq�T�A�������-9й��s�?��W�"�+#�i�P��v��\���55 �ǣ�=�`i���j4�.P(����K������U�/��3��*)ņ�Z����j�ۚSp;�}�����A��懄�P�":��:���%���k���i,d�n�r�W���5v���KT��y��%ҧ��&��Ҥ�SuN�����L%�X����o���ـ��0�Hi6��4ѭ��rPǜ���`��֤��`:�b�{H���(�'�+l����}*:�ϭ�r�g�9�����ý7��D��Z���/��iL���%|]f!)��E$��?��<���S��b(ML�&EZ�F��	�κ�д[�j Hg<f�,�iT���Z6�>B��&�<w��xF�y�k�?΀66���n6�.DU�^9�l�{5<K�/,�����Q��h5����=��G>����.�O��|�ߐ<��;�����ɿ�k<�oJ����S��)���>�` ������G5L�~W�+hZ�*e�x�]X�2nR� B�3�j��+%Q�9���h��5�[��� vL�a"�Bq}�|���C�RA�U�����b@a2?���Btz*�Ir�7�ܢN��L���-�\P�H�_}�(i���<l���:3�z7�.DFR������7�^����"4�C; �}��A,�w��{O=�㯟Ʃ���Zh��@���VWNFހAvi���m�iHf^C�������?����7_8�����UC0:��lt*a0����9�7�_��C�ڐ�w<a��q�ﾻq����t�
�|�$Fp���h������4�#���A���s�/�ӟWs�c��@WaE�_-�"�g+m"]mi�o���aaі�?�U�s���S���^x�;�@;RZ�lЯ��]�+	��Z@�v�jI��T:�P��!mq�#A�~����)LOOcr|�x�v�F�c�<��K��1�=�v�J�W�:7lt��Wѵ)KWM��<�Z��ssx��E�b(��87��\����	u�m�RTı�����! _�'-�(p���V^�`���s�p���6*�V=�)���'�f�jN�lm�G�' �0��@��VZ��攚��ǃ�������$����hr��ٱ�sH�.�G�?�BK�l�|���@�Y�kA���<�,i���^+��ÇɎ<pk�q��$
�(M?�czd�L�9i�磆�O{��i�	�D�wP��&� ���H�N�rS����J�Ɛ�
v�=i�Y=I�g��������!���H���ÐT8�{��m�<*�ɝ��1�J�}�sIZ�2�Ic���z��#U����S�C�HK��ɍ�g!��m�R��Zk*������,$䳭��N3h uD�����ę�v[6?���~Q�������sȠ t"��6jբ�nʵ͵��M�I<����1Fl�}���bmmM�|��=����%Z����QL���*������=�u�ϝ��\�����m���j);��u�mNa�����^]\��jmX�4��}��I�6��%TjY�A:| {voמt��
��t�L�� �~>�"+_;��r}�>�64:��� ��.��aj< �TK���
;��h���0BK~�`8�h� .��ȬgU��v0FZ!�) .^�ًW�J�^ϭ��&������ۄ���`�L���'��f�\��م�[}DÈ![�`~iU�qf|N��������T�������_,86ڛ~�>�9����w��ym�b��(�|��E�JT�?ژ8M�66LZu�.���i��7͉��$?�<mj�$�1�2�j����l4��<\�n��i7ѪT��G]��{����GMa�;wMa��	Y���&�� ��L����C�����÷w�!����.
WWHQ"GG��D����?;;��0�/����������n؋J�����5��64�Ȑ�x<�}����u��z�ͬ���u���%��:Zg��셹�=�"��E�P]��&��_y��#�NP�D�23#�d<�l&��Z�h�z]d���u�1�|14�h�_C�����A��/���Ͼ���N^���>*g"�N�Ft�=wȁ��O<��'O����&�s�=ǳ/��/��/���+rW�!C�� K?�!A�s�h�Ҭ#�c8J�Џ�4��Х�F�uN����hM*��2Q}A"�ԔQG����i��YGne�b�3DlD"յO2���3�P쮍��CP5�t�j�^�2MAzpY^�,�jZڌF	�q�{md�%�[}�b)D�	x�f�j�j�6�k
ض�����L(��@��:��}�1��-c=WG�� VXa�e&۳q�]4�o�Ԍ����<O5��O��=�~䋿���6�����!������-�����I�U�qJ�B�Dg-$�.[SD��
".�RCp�mסWf/.��+bppP~���ʷ,��������<�����R���d�9�1^�t�PC���5.j��.$?y����vTK����o��μv�䟐���M�pʊ�1�|����A������+QgW��*�r�������j�}�y�hB�� �i!`��1�r��߷S�Ҟ6�.\�>z>n
$Pз%(KJ6�/=r
o�[F��B���|���]����ot@������x��G��-ѓ�<fO����3�W�J�U����D�����3�(ͦ�( R�@��Ŭ��m6��x����N�q��[���LCpumm;Q�PH���֕s����-Z��>�γb�w��2@�4����s`���Np�������;�~�<p|�up�!���vp�sTh�9超����j����M��c/�i<�~�k�g�O!3����r�����]�E�3&>��Ιr���+:m��o��^�𾈊d�٩S :����4�g��Si����>qܔ6ayiK�-�¼W��#Wӆ�IQ���^ۮh�a���''��s6��S�}pȔp���ҫp�.�~�>�5>�@�S+Q-LpC�14f���2�ev�#��d^����$��pLa5�>��sr�Ϧ炰�M%�L��(��a�E��d6��2�ʙ�I�1�6��gC�f���Z�EoǬQQ%xo�A5_D)(��ǵ�9j`Zuԫyt{5���a�]\�<��匚�h4�)8���7���/:��R9�=�{��P�����m�(�汴�h(!���䗅$���59�޴_�ǒ(W+������&�&0�e�XTڎ��%�/-I�BZ�2������M7�M7�0i�Bz�RD�Ҡ� �Á��"2�%,�籴�A�ц7��Y��|M�x����8�2ǭD��Xn>��P���恄s�9���%��I���{�f'#���}�F�4t��Wg_s�x���GyM�;S#V5��� 3�U�T���a���d��U����J����S�cmyA�d�P�J�,���EL&���f�T�DD|��_����.��'�!��v���WHI%e�L����I�醳���m���8�;��u����Kp�u���h(�͘vB~\�]�?}����w�@��B<9�ip��������k�ݦC��0�އ��y+n��0҉�PG��y}B�1�G����q#b��ba��l���q�"�9Tkh3���&%@����C��k�����cnv	1�������f�k�~�w~�x�v��$71��^X!&����3j'�X1h6�o��c���~'N��/���B�n��x���B�`���Ǎ�?��P �mC��s���X\�}��s�B���<ڭ��YXC<�G��G:5�~��e�W�U'9} #7a�D�6ٌ�A��o3 ݠ�fXi�Y��Z�<�15�'<+��{-,�����#�Jcxh��4��0���k�B4�s7Fv�C/1�~j��'/���'�ǋ�^C��W>M��4������8~^b��    IDATc�ϳ�::j�H�%�F��n�����}�����b��?|��hC𧏼|������\����D�\L
�x�:�b�9}�t�� �e;ǒx�����[�����&��qs)ReC@�;k:��{�|�����<�1�^�`1�ž��=�Q�ȀN'�DP�h��T.��_��=I`��l�N��^����x�<@>�Bi��7�^ZŸ(��aE#r�`S�~�D!=�;6�g�m�Fd`09NS��v�Ѩ�U�#��!7؉����m�8��m�M ��S21))���_^x=��}������/O ��@$�/L4�"d/�L��H�.�X�x,�>YBa���+�"�AHn4�%5s�O�_b07%�z�&u�T*�S���̦�>��l�ٜw<�ʙ� ��)Z~5�NDq�=�n ��! ��1/b᭿��&�׏6�D�ݙ@r3 ��M���I��D��{x�8S�%S�U؉�>Ŀg5`0�s�"j��|��ۈ	?�C���M"v�F$��B���(�א<YM#Y �I�lN6Q8�g��i��i��-CVv���E�f\rM�5uDߢ���tz���g�n��|s�ߘ|k
Kʘ�۫�н67l�0n��7!���h�,)�j�fN�g���?C�Y���<�w5|��Y(̣SQM�"S����tS��1'Eͦ�M�mG��޿YC����Zu�T:<r�?���hj���ϝ�RO���b(�{����I���c�G�'�����9lN�7ܖ��6( )�>e��ى�3N��IPI���3
)�.�y�>��j�|Q�@8���
TsWl;a)���z<Ba���2� ��-"���Y�X"�����T������R;ʵ��e~NR��=�J��6@T8�z���EMȎ�#�#�vU����a!9�֧N�ѳǴ��z^�^�# @��a���@�n$���}���ZW�\��ᗹ�5�Ú-��|
o�8"X���cCp�b�������&R��.d���zQڌ8?���k;T$�z�<�����i6$�Vrﵟ�P��`:���%�%Q��DH?\[*0�Jb����8w�
�
�t�
�P��Ѩ�p��C��G~����q�S�)��ك؀�i�glz��G�٤b��[4����C�<;�?�=�h�I��@���M�����|/��=�U<^���h�FE�/�>�3?����6�xx?�4/�QN'��d��p���&�kC%�?�����h�**�a<�3wXg��h��d �>��0���|�<�«�-�Q)1p���e�p� ���;����M>�	�8�\Y5J��Z��h�<��H��-lm�@4:����Q<�w_�Z��V
ylsߕً�fY��[��!\�k'RJ+�M&�k��Ye֖q��9d�W�����߇X ��dt
dmZ�SP\D�hJ��Z&HJ"�U04�D:!��YeQ6M��m�}S��A��Q�;�d6\=d����ʨFrx�d�XWV:�����jǅ�zg�p��9�~�<��`���� ._�f����|?ls�V�\��q�SD��x�}������?�yo�����hC���|�����|�Գ��F��$�	!w.sj)Y��m��qc�� ~�����Ƅ�_ZE�TV��S�@���+���s����(C�����'�#���h�tKv}�ЍK��K�	�7����H-b� ���x�]B,�C<�Bu}�?�$.�8�Zf���[���DI~���#M�b=�G4G<�ւc'JGA�#L��G/f#��D������`*r(k��r�!<�нؿo���1Ӆ���Vn���ᱧO��L�kMdJ.�"i$��55�D���ϵ���ߚ00M�'{t� /�Ԑ���)��,������.��KJ-a��������"��7����z����Hx�X��DRrM{�hC�XG��Fܘ__Cop;g�Psl�"Ûw�h�@s��7�y��s eN�w�h5�9h��F�V�o��Й�I�����Z�qMɩ�\�!�k���j�ɟ	�Ѽ�1�[t.1��-����o��D�v{FwD��Ԑ��i4TH'|.���257.1*�mk\��P�VE���F����'즀�
�k9��UG���p�L����.5�j���b�)���6�L���kſsP����E����P+�i���0���-j�B�LPfo��ȧ�ܦ����x�w�9EU�a6���R�d&Nא�����;�J�MɰΔ֡��&��R�)��arl'9Ø���Fw�v��㇛6���f�#'�_j,l���)״g��� �i"�$�e�X9���O�<݂��e��Ws�k�� �:�:h4���Xt�"�ד�����4Xκ�wS�K�g��Q�LU8���c�;D��Ա�`A�$A^O�Z��%��ѱI�ܹ[� \���8`��zx�D�4�r������A�[���;q��.]�7޸��.���ĵh�k��c�s-c@͍��4�,W���#^c�\\[7��b	T�R�0�4���ݔ����+�cf��5���h8�����?҂�#'�������_x�\�@ >6�ժ&�a��vlZ�0k�=gl:m���q��7���p���R�F}����6�M��m�A����}S&��D�m�E��K�ى���l"�+�z���!=�l��/}�[���:2��\{>�N���}��	m!��<ʥ,��/����ߏC���̊�.��z����{��O����)\�~��^'C���W>�.���lL�-��7-��4��R�������7é7����+]��#��W~���mo�Ig:,����:�H���<��������U�����ￌ�����y�d������=t9جЭ��jԐp��}x[�i4�9�l���I%cj
.�?���3r,#e�Oξ�':P���«i �P�'�d�k��tl��yr�����e������j��:���¹�^E�>T'���bhp�X�h�tV"+�!2:
w:�\ߥ`���\��󗰚)�W����j�Z�IC=�Oȸ�1�X�D��e�`��j(h�t7_��}w�S��K��&`����6��/����ߖz�����}3Y���%�2��D�.m0���*a��m#I�����ۑ_X��S�0O�ྜྷ�E�]e�7�<`7�������/�Ņ&ڞt=t���&2S"v�|�X>u���-3���Ð�>��<�u���X�.< �y�+%��Vp�Q^�L�,��S�k[Z���WZ��P����h�RIŊ(Mz^w	��b�DtM�p�H�aNB���C�Q@,������wb���������ե&.\Y��/��ϣ܊�o%a��Ix*ΫF*���=s�ІO�;7Szޓ�ۍ%��k�~�Ds+X�0���˨/�ʩ)#�0��R)g�������3�s67z�sj �<hh���K�4Rg�poj:>7泫h�<zP��Ξ�+s��7��fm ��YC�����#T�cy�b�<M���tж����Lµnl�9�Y|sh�����ms5̤���G)���iI ͢�43��j��6	S�f�(	�	�S\pZ��:�	C�Ź� ��g��5�5Ź�*~�`hk1t�i�j>�S�N�É?�]�l�����7L����s;���r*��ڻm�Cw�N�vҚ����;M�S\���,' S0�гiT�S�fϦ|yY(����~2u���6į����_ܾ�<�L���k��L�c�nNa�8�8��:D� =\lE6e<08hq4.
3�ٶ�,1h�,q%�p4�hV�ۙ۸D��i4ύy?���bR�I�`�_6��Nb[.r!M�˺���FM�V6��>�咬�����(�^���@�/l<6:"Tz�$��B����8�LZ+,��d�ZZ¶�T�9�a�?s�e�}]����4� ؛XDR{�DQ"EQ�-�O���l�qދ^b-/�8~�q�$�K,YT�Z$�E�I��@t0 �o����������<-��Y�̝{�����>��w:�D2��K`͚u�Ӈ�ʒ�gP�6�L��/�u޿�T�ꠇ*VOM��K.��T{������Q���i��+�f�hVx�<�zO4 �����:t�L�6�s���W��Y��`s�@l{��#�L�^���p*Ӡ*y�D�GI�!傒ƹB�׮V���'Cu~��t*k(fݽ^�#��2�����eT��p�-���~��᪫.Qv�Z�NZ�)�	�2��1�e5&�8�Rɽ�R�ܿ9ߵ)*��Vș���O|`�hʬ��!	����w�����������Q�cT���>'g[V�c�,.��+^��~�}�����Bł'�:�h��,9-@�:�;�*���(7?x�!��9O�'~eI-��� ��Ro�?|�{�ع}�Dˋ�J�G��k���w�"���F�S��g���$'x&pX���##�3�SK��K���>�:,sG:�sQ�I�d����"��&R�l51�L�3�۩S����0Y���-�cu1���c�?z
I�bK�vJ��RX:vL���N��J0���s٬��t~��h�.�II~4Z��5�{�*���b^���(���L��126�3�<GeLR��8V�!51��-�a|��.��ܞ�x��,�Ul�;-����*I�֛m5犣��Tbs2���3�BZ�,���a@��5���7}��?z������~��W��?��?o�F�/�یr�E�	�����j�Ь�D*F�D��֏0�N�>7/����]���}��݆����t�5N�p`��/k^zmˍ�Nb��I���j.\�) q�]t�-�si�Y�c�9}�;$�˥%,/�����߲n��w��<��xs��[�R2���T��[)�/ 72���ˌ>m�{NXnd�pHSbS $�E��@�e��eՊ#Y�s����w�k֌�*i{�/��_ū{��|�u*�!S\$hD�E<fTWwI�C=�Wv��2F�:X�I�p,d��d:���
J��K��^���νX:2�����+��Sw��ryI%|>v��ؚ��{��O�B���agƝ�$�d���?>����
׿�6�i,2��h�j�x<04�B��Z¢bDx��z�CMf,���Ohf�Z�{#����vp�l���\>�x�����~ ��m���|�������р�KM�ZHIS0��d�E)3qS&��:� G\���C��q^����^�[�#��2�*z��sɵ�*�^�f�����+>s��A���!�McCr©�Ōs�4�GOz�oo�t�st<Np�V������:�I�avЛf�lЇC�4(~��h�+�Rx���FIX(�����܊����AU��^��4�a�`�5�Gz08Ol���޶�	��{s0�U8� c��ϟb�H*�g�Ǫ �'��h6N7�A�{I�#fr�3�+LRP1�z;.��;��k�.���e�y����5Z�Hؾ#3���,c���ۺn��P�D4Z,j��h,��k����,C�\>4|���S�6�"��̑#GP)W퉽>���''T��&Q=����*��[bÂG���K�f�{x���iY;S�� ��_���u�Iq%B�Y��b��	J�Ze�2Iyw��N`�Gu�L�h�G�)��r	I�Al��t��_RB�^�M7]�_�ŏIΙ���l`v����߰w*Ẉ'E���):������mdh�HF�+��c��W�AF�%E���~��n�~�\bro��Q|�����|Dҳ��6�8>i ���lZ�����(���,^w�9x�o��/�9�y��a���0弑f��W���x&�Y�G�c�"���P/ӛ��)d"����.&G�'���A���\���<�8>�ůa����Y	��I]�j�m\�vR	��ʲ�Xm���S�O���C�-Fֆ��◑����i��G���<I���T!`���"�*f��X��>+�&�EQ���D]^F�R¦U�p�i�o�Q^�W�p�6����=Y1lw��T�a�R���E���Zd����ϣ��z��RI�g?��"���0�U��
��#EU8ټ�錳�.�Ig��l���"91�5睅v����"v9��z{�b��<��Q�(z@�,V�y�3��j$�+����3##�.R��f�L2�c�%�z�8FR�g��;~�|���hd��ݟj��?~㉫�3��%��ݰM�7t3X��<��l��Zm"֮�[YF���vW�w>>���5���F�"7X_4,��	�����.>�����9�Zĳ�Z�#��F�{�q���q���=Yrǻ@��B�N:�n
�&���eeF�i�f3X75!��~��g�p|z���K'��S[^��'%�W|>R`x�$�Q��2����3�s�Z'.��4T��S�^A�^�E�_����7n��ޱc�8H��gFO��է33���h,oʕr�2�7�K=��$�<7�LJ�9v�+��*���mT�e4��X:8������2tk�����p��^�2�q�18r�����D��Ӕ�m�[=�+n�VA'��������eR�H��QMf#HN�NS���
b�H��xpC�Ö��4c*5G�G���ɗZ�T@(41��g��4���Nм&���\y�(������Ɍ�"rMʠ�0�3ޤ1�@E������$$z,�JQǵ�{J4(����P ���.�f9aK�����D�wݣl0`Q��d��E'eXD3�a�.F]���b �2�r�M���D�-��*c�kI���A���=��qg��R��>��e@+ȥjZX �4%�b�P��^	���xt�\
��g�nܾ��
��<K:�ty�5�Ɔ����K�\��y�yo�5���Zp� N�fLiSֲ th���aŘ���C�@s�W�3�~�tٗ�?t��3u��G��Qw�(L�>:�L	����5r*�d�W�(�y��Z�FG�����ʞa��oJƚ��{��{�����&:�S�z���@���[\���*?�+=^��*�������,{�u�6���粞�'.\�4�%�2����u�6��������@�۪qe�llԗ��Oca��49͓f��N����U
sؤ�\�^:WЪ�p�W��~���K57���-�~�o���/*+�yE�+s0���~<��>���,k��HqN0��g�=>A���)�%��5'?2����#ǰm��9xTՁ���D�0�R��D�ɛg2�F��&��F�Y\t�Y8��3�\���P���y�0��elJE�{eɟ�'���O��Z�RG�TU�y�Tv�gp����3�2�r&�R���<���s_���#!�W&4�6��*j�E%Q)��UT(u�!Hn��5����3�A`/e�R��}���E���9��Yc�]�9ߪ�8��C���F��n���#yd)�@��n�J=���C�X�R��H�u��K��]�uN.�	�/�M��bE�%d��r���b?A�Mڭ�����-r'׭Q� ��F���踒Ӊ�1��I,��8Z)�G��~;��2��FV��Kcvn�rMU�|��&�@����կ@�Ca���*;4#U:�X��W����g���7}��?q�s'm�?�~�����������?_i'�/n:=���}���w�pZY/�O��֞d��N��~���X�_v)��N\~�Z�V�4W����}�L����E|��cǁ
j�1$����Ry���X"E�R�d�JH��~�b�\`�=������Z֩�h�Zg�e�Xb��i�)]���֮�S*ce�N�?��ݻp|�>�F5ₛj	����5�X:J��W�@eJ@�t#n����v�ȌOb�gb��3��\��̔C:7�~��X	�0ӓN2m��*J�%F�l**:��L�/������ټm�q�1Kj�q��3�W�X9>�:�ҩ�2o��T1AGN�,�G��YbL���1�8����e���F�AWz����Utpp���Jj���%���t�m��7    IDATӤp�Ų{;zD2�^) =����OV�5"?���a4�MƲ��"9 ��{��$�πJ"���� �|�6f���2���v�@A�����H�;n*>�-���$c5

`L��><�L�ga�gȲ(����";�E������^|R-�l4P�&UЂS7��5Ǒ/Xf�i6����2������e��^j��?�E�4�v���v-#��e~ך��q� <�z�9�3�=(�2v����)���Ѓ E&5�M�Zs6��U��Ï�z <�$��Ж9����>��;�����.5� $@ۿ�z�ϝ0�{ʚ9����(T����k\dV�����5h��g�Ϝs�Ϝ��}�᜗�":�U������c���ps���]�Ic�~b=ދd��x��k�גyҰA� �~!T��ך?��9W�5;2��^�A�����υτc�����U���< �@x�w�5E2��x�bM�� MP�#,�h�&�4�N�M���ʶ�
�,,E��_��(���r���r~�@ݩ�K���2������	�@�lQ܀�#���=��w�?	%�������D�=�6�|�>/���&�TI�#_�����I
t��UVy�ڵ�D^X*aa�&��5p�����h�%��*0K�<�# �~�f�,VD�
՚�C����s�f����F=�(�>�3 �Z����܊)�ߪ1	G*��X��U�������{~l���w�xt�V��/|Ͽ���6&�+E���̪�H�|H�b���@���S	��1��k����Ϭ�ɢ�J����� �"��$��R�d?JW��
hXY*$c�0:"vu�&3)L�3�p��r�'b��Uj��3�2���T�SP�B*Р���qV�E���]z���� �ϩa���i[N�i��hn�9�c+%�,����Y��x����q	�<�������j�㨗[��9�>�:�khI>)�Q��F+�G��=Iբ�r榐IeP(d�j�@�S~杷_��>�sχ��'����7��������R;y�������0+cRB'�fr�S���:�XU��b���sq�o�EgN�U[F2�����q6g���G��Q���r��$z��� �&s��i��+��R�綍D>�V��z�j&\ɔI��%-j3�48����JiY��ѱ���($�X��a��:�Kx����ٷW�
sǎ�SZ6��h�Y)R$�9�X���0J��*n(�HԘ���Mظy2�Q��^�.�L�J�����E��B����}�����e=�hfe1d��$�J��	͊��jXN'g�Mz�r��4-�dmnz۞xG�����qU������Զ��DeȖz5�����%�hi�#�EUz��A�Qܸ���&\��۰�i`ϱ�heR �΍�{/��9f��ݬ,�0 ��e��xx��3m(l>��ឭ@
R�j��2��5vZ�س|�T�,x���(�?��`;�f�C�����@SP��x q�M���mt���@Nk �V#�=�;��J�ˋY**]*tp��W��V/4�9��ʹ�ENYp,ץ��W'|��5:�@�8�b,=���T43:�%Cω��"{V��!��~dc�Xʳg'���c��QT���Sdb���VC#+5�������"�5�%�	�D��3sE�Hc2��I�@Ф�B�u��l�(h�'�����)�f� ��i�e=g�Ư�
�*�<�~�M���eߊSc�|�(�=T�Bv�b&j8$���=��*�%UHsP�t=���f8ۡW�`�`�@UTCW+�>�gP��P@kn��+�x�
�,���w%�����m"�f`ߛ�*b����h"�i%��'��J���^�h�
M����耒�&zV�,�
A7�==+�gw��������2�d�P�Ut�T|91=��܂�űv�$����S��UE�S��7���K�UW^j ��ƾ��[����3/��l�fzt���0�)^'�g7�A�ߑ� ���cC��q�E��$rycxe��a�Z�۰^��r����T	�{1��cX�z��`N?��Ξҋ����ŪS\ �^cƹ!uD�i���i�8�J�~EU��UQ��GưR)�Y�Yi)�� 3�F
� �S=T�J�(�ܴ��x��L���n���>�.��O�:�L�j^iv�ǟ����ں�NRtY���*En�6�X�Ғ���W�[�,F��:m1JՊ�a��I=X!pW -��Ћ�)�<U�xN3QK�.ǫ�kJ��j�m1�Mc�1L
(�ۘȦp��5�85�$nu��X���B�j��ET��~��q,P��INJ��4ִ��{�\'�s�R��ʓV��}rM��i�3�w׮[��u�P�7��(�/a��1̔�HM�F~j����C#�Ś��R��}�d�jS���� -;��I�bB'�}�O;I˓�~��ݩ�V�G>�|�]o�����c���G�������������̟1q�Yht�J(Cڤ�S6�z���{)�G��Z=L$Ӹ��;n�y�&�o-#k#��]zZ*16�ā�>���ڋ����:�LW,!�	>l��\i(��S�J��J+���5��nM�Ծ�!C5�BZY�z��T��M�3S�����<���<\�e�$��)�о���SO���=�4�.�/�R*���j�5�p���(1���*����U�^��ι��4斀ٹ
L�����Pr�%R��L��h�pMsB�%�&�덂���r[l���C&���e8�l�^�����K��x�����]譜��͌���P���=א-7g���I��Д:��3-�&�;W~���3 ��M��ͷa�����Chgɷ�˚��1 ��Zڱ���7nj�iOW�	 �A�Ξ���(0�� �{So�-k$�	&fEl& `p-
����X�jieſ,���Y6��>�$�w'ne�)�+�����Y�2�D99�m�=:Pj�7��L2�1J����\���y��a����yp�\sn8�&�=s��&
�4/�3���4�a��[�p�,��7����蜉fs}�x *p'��Y�25$uP�
�z��V�������7&dB��� �^D��k�'��t$��u'������k�੒�5(N��*6���'�qSf��$��Mt�! �;u��ż<��t
9���H1���?��c��!���Bo�?	0�I��H:u'\u��%������C�?9��x��'�ao���uƤj= pRu#4���0�s�Nʈ�C���
MN����W0��`�-���x��X�X�J��i0g��֗A�sO�@�M��H�����bi��؈�g��F�%���gqp�n4���o���0��{/��
:͊T��r�����]x��0��>��K�7���4֬;�ݥ[���3;����q����<� >+�֯_���U���eq2Y�V˘�[�d:�G�C�R��F䍠�o�kT�bZ�ۄ5\�Y��f�I�n&0::�
m�^{����Ie����j�b�@�H���P��FM�ɞzE������z���&��
A�����t3���6m� U-k|g���7������̂X�]�R5ʨ��6*��Y�4i��\A��쑡�K�Mz�)����%m�oԱ��s��+���PO�W�������t�s�RF>C��b��Rq��}��a.��|��i�ԬJ���lUj���>��j��6f��2��b�8v*	A�4�驊EU��kg*^vo�W� ��x�t���J an�T�k3GQC
�USHQ)��Z68oX/ED�w���R	ե%�L�r|H5d_U��Ud�����N�J�Id�	l��ј����֟�?�;�{�?���ӟ����������
�7��߂*Cxq�-*Zq�6Rb�!�ٶ'a�R�R����*�w�M8k]��
���3�,�р����/e��,/l@vtR`Cґ������y��b�NҲ�A��	Ө"��j>�2�H�hqQg��h���C��fe�^�L���L�q��I�}7;`~vIe,Vfh���*ڤ�v*U �1ڭ�d��$�����S��@���J����B�T^��Z��T����d��lyp�%������Nl�"��`�)n[���<�H��uQ���h��0��n���
��GE�2�L[��(p�3L7j�r��ɔ!r����l��,�fzhƖ]�W�~+nx��(u��ulʡ�䯪H��w	:H�a�d��A}�:��v��YW��t��0x��Pu�L$�.Ff6�l�[�Z����n8h����E�����_ `@G	}=<$Y������ �v�l�����/ dȃ���E�"��iX���R`43SR��_&_�Sde�g`f8��)gN�ч��Tq�X�U^<{-��S�^���@b�K�?d���$x���g��CҬ����PAhҶ��A�A������@5;�0ʨ�<� �
թ*}�Y���T��:$@�QQ�Ɛ�&�o  ׽pG�>�Hf$-X�n�lB�+r�b)f�$�hN�J�!e�c���|o�\��v&df�>e4^��h��@E^W��jM�������1�Ɛ@{,�$p�~,���{ (qܡ�fB�?:�ˀ0f �e��6�9n�r�������_�|sJ��'��G3�>w5����/��CN����(p��s:��y�� �jT]V�8��V3��;bjbeB�����~��fm�^O�-�kaϮ��k�NL�[�[��O?��݃�KKK�?4������'���o3,K8����mw�	�x������D����[�_�q��,��QbYuaO�V�ʈ�m��2�+d~61�J�F�Z�
�揋D0\���9�K	��yy�Yg��.PUb߾�8zlN� ��"4�LJ�6�dU����s��(	��Ϟ��D�� ��Q�����H�d�;)Rs�����)9��d�0�B�
7���b�~�u��O�slܰ
4%_iv�Ҿ=�����Cx���p(P(%�&i)�;:�e�cb�����^�4 ^�S��b�}�z>��C�6�_<�H|	��Mn�L���F�L$PV�> ���?�vkFGq�y��+^/%DVV�PZX��	A�g"���q%�Yɨ�k��}���d�Z3d��T!e���lު?T;cS|�b�VAf��x���F]<Ɠ8tb���QdWM"�z5��+I�Q%~d�k����
ZՊ�S��[�(!�(��t}�����(ɝ��ۦ�UF�q�Ve�|�[�����G���O* ��?��=���_��~a��������7����@���+�+���q�v�Mt*u��Ҹ���p�m7�u#��K���R�aV��g�W;�W^;����s�5͞��
D���أh��ή&{�,(۹ɫ���O��I���"B���]��p�Z��%��c #�H�\ZU{�q���� ��P�ʕ�]��&&УT_�I�V�r��5�r4�T���F�d�M �����<M~?��R�^��:ԣMۆ�d�[Щ���-��(��N{fK����&u�A>`�dZY���B�WA�F�	��j��H$i3:��X���{��6T���o�8:�Mdyi�z�Hd��0�^����4uӖs;�إ2����V�kp�����܎r��׎B���J�����L<�S�ԕ��#¹��ȳ�C}w�Qn�oZ�(4�&�����R+�I�4����D�?�BU؜H�(4�w�P�����>�ܘ)��@���N�t�?�q��*8pl�j�6�!ޗ@����*�]KI �=*�|8F��Ź�'����fH���'���9����Y��̜���w��4T^P��=(�=�{�oe��+e���`�4�;��h �
Q�Ș�����Z�7r.,P�%���S�-ЋɝX��@{���~ŋ��J�{���k�3ն*�2��5z���ԃ2z��
�T�B��ԦT9
���r�r6(4��h�$��x(`�qt*ؓ��ҟl�7J�St��T�"�ۘsx?\�*���RA�#�"߿�+�R]ܚ�ɵ�����!�p{O�<���d �zBk,TD7���7��� yH�1řA�R��<��������ak�j�
��SQY1�R�_	��%���ʔ&��� E��
��.֏0�I`����S��x�ݷ����ѹY�x
�;�`�K�o���0q�e��*#k�-w܀O~�ø��T-f������[���cؽ� K���_�ɉq��<��:|� e2�h�Z�S���&�����v9������2���YUje�&b���Kq�e�I���Wwb��Zp\��G����P�?��D�rIs�k�Y#(�a|d�h(�ϊ׳����\�a�V���p�{h65�|!(,�i��Cy��V�4�$U�Š �^Z<�x��w�u>������H�����Ͻ�Ǿ�^~i�i�$��굲L�.��\\~��(����jvu�����#E6���1 �S}��R�o8���ryE=�!�3�k��e3��@�bS��[��VuR���T�hV��������Y���M1I��f�e�Ӡb$)I�������5]hq�YRO�����yFA Ek��+��ԃ��g�j�E�'���@���R������SXi ّUHgF��+2���9,5k��H��	^�T�V,y*�x��3 ��Eܜ̒	y H�����x���f}���S?��;?�ǿ�3��(C���/��}�ڹ����Ӥr�m�ٚ��Cߝk���܉n�X���y���뺫p��Q���d�Čx��c%�n<�m���ٯ=�=3�����2�I�q(�S��c�j��o��:&�YiW���>#.L�_�d��a$?��}E�}ZY�F��(YfĻM��2���
*�%�c���KeU�[U�Ԫ�(/�P��vd|Cn@��'矍/lRZ*��\����`�@,��(���h�z��3��<;XLI�So�q��t���,��Ӏ�{�ֺl���8���/�#�Q��[A�5�0��?���c���|��؃riY��~(G(U����� I-��$5��VV��@z����V\��;��m㵙Chf���� ��D��$HN�1�L�󬇧�0��2����hCe �Q:	y�:p���ԒBs�5T��{��r>Z���Ã��^ga�5�q�1����B@�𣴟�A�,���5�Z�0_��mW+؉f�# ۲ ��B�����4o�Q�f��D����TDf?%S��@%�4������^ �r������%��U�N�B�'����r:���<,�Ȑ/�/}N��ړ��0T7B�i���Ԯ���QjR��d -<�5�ea�y�1C��`JN f�U��4}���Af���
:��uoTfb�E�t�ZH�ވ(h��`�i�(��RT�H[���z��){P���q��&C�ă8Ѭ�Lʿ��S�l�ƨD�W�5�h_��� Ga]*0�Z'a����C���}ݞ��D׌�s0�S9�>&Wl4k`�g�}-��PE�Vx���JV�b��s)�|���t��s8��	X��>���P����ҺjO��#�E�2ҰT%�*�1\%Jbw��:��D:��{�c�ӏ��ξ�
\w�ͨu:8|h�^��������\�Q<{����/�ͷ��F|���(�
	�_�{ �z'���o�����s����~N߼A��+�VM�t�pM�zbaǏ׿��9���&X_�~=n��Mz�t�޳g��0��)j�?~s�X�n�;�<я���ѣ�5^#�Q����2��ǉ��V��m��b_��t6m޼�s>�F
�s�>p�O�Zq��i�><3h"�WS���LNMa���Ԥ��3���wan��^,-9L��G��7q��oǧ~��X35&�J��������}O��K8t𸜿������F	�O[�_��w��[�E��6U    IDAT��L�V�H�rH0��f���^�KU��I�eOf� V8J�e��y��łƏ��?LR�4�
�s��qh���8���9tU1.�E�gS�>���n�Z��O�-���"�ϝ�H����I�Z=��.�*�G�W����7J�=*1,,�(�d`�^E4gm��f��S��u�Z�&�lD23�D��n:�x>���
b�rtU.��\Z�̡CA 64�7�.J��7!,³�B��	���:�y�S�g�}�M��_y�K'������S�!��������_��Nzb�����"A��ߏS����V�%P�vlJ)�NS�
'Y���W㎫��M�]���$FRT�hjsϏ�����K��4^�q���8VΡ�Z�J7i\0ʍ2��p�������e�ʁf&�Z��fMU������/���4�|F��r\v�K1�C<:f-�U�	�sQ0���@v����F���$�,Sqs�aT��X�0&���R�NJ�ȬSɀRY4�4��i���߾޷PȡQ�����
�ʫ�bQ	K�c�TBcv��YZ\�k۶����@m��E�1��{�.q�������N�>�̪M�D(Ys�O����[n�MoV��;�A1G���0 d�����CV�dL�Yvp�ˀn2u�8�����C}����Lф�g2�h�^L�=���`Y��u�<�sr����!�(���(�@h�� {��m΃�<��g0��/�+~��'WB��8T?
jHݞ+~b���L�gn���o���9�U$J�� ��LAA�!<�ISճ��4����fe��,lA{-��t@�Rnh��\�Nwwe�<Hl>�}��
NӧT��ЏQZI4������A?�0�0�>u�y�KT�@�a����JG��#�dR��g%�=r噅�P��/p��W����Rҿ�7)�h��,�C��@u�п%H5��Ȼ+x JΡ�ިJC�zL<!Wa0���{X�<�gә\ўK��BA��T�h*���Lz`bh��n��Y,��g��`���$Z=�k՘G��55��%�ϡ��]���B��Ẉ���Y�n�0&����n��1�����}N@��Ku:E���v�*����"�ڇ��y�n�]�z\{��(u�ؽ{/f�cn�4�/�_�#Ɋ4��4�c��7\q~��?�7^u	����2���G����G����o�[�z��ޟ�����ȋ�@��m��]XX�=�����Y>|XA��_�w��.l\�����#�<����,��@�0}�����,yfR=���r�|.l,^�n����P,..+���sߩW+J"���kar��k�ŭ7߂��ש�w���x��`���}�Y���˥,#υVO���W���8+!�Jm��
X�vJ{��Wv�k?��{����*�
D+���7�7��'�z5q)CM��_�����xjJ+ud���(��~�t7�r~����9g��e��� =���=9ڇĈ;,k.�������~#f�j�E.���Ϗ,�<��٬��M��p~�j�ш*K$��e1"ڕ:��2�k5�g��5Vl�Y,U˪n1�*ݶ;]��u4q�wT*W�J��`�?g�^�5(��g���s�����Mn@ft-:ǓÊ ��:m͟����f���_|�Z	ٴ)N1�#�#��	��zп�(��&�XB���&���릏���y�$0�����_}���W����8:~z��J_̀z@`<~f�J��7�j$,���])��vn��R\��8��H��T��IǸz7�.UyR1<������Ɖj��z�W;ʞ�3��!%��T\�g=V��G&��o�ۨ1⬛l�K��\���L��:��&�uX�a-
E�2&G�ef��L�'%�=5ɟ�r]Y��Q��Q �}3&�51��(.�S�e3�:f��C˃�\/���M�U��>#WՐ�v~.�:(���3M�6ҩ�&m*�C���2Yѓ��c�<���;w`f�.���Z
��L������*�l�:�0g��R-�}�64KIc������7߈����6��8����֠$�fn�y3��T\�(��E'1�?nCn�9ݲ���5@�kA�yW}�^�H<<��w�C�i�j:�ud�4��l��_��U��;0�<��k��u��!bWAN���E_b�8gP  ��J���C���Q�8N*'+h��E_�q��tMAJ2
���>�;Q ��
�=��8Y�ҁ� ܠR`��A�0*�载�c�He7>��Z�.r�N����$�����������F����������T��q��/��F]:P��!��]��J3��0 ����Av;PTLrZ���0�g.`x󪼅�`؃b|d�읪�*N��p��`Z�C�|��)�p��a�>)c�b��� ���������@A@O� y7kc2�ǭ�(�N�� �r�N���a��������6
��r����2��D�<���N�ճe%1��q'���2����a��s�oE�S�U�\��/{fV�L���q��?��|�z�f�϶�������������rӎ���w�],�T�w�~�3��{7x�;�<hj_�4.��L����t�������?�kټy���ࢋ.�SO?�/}�Kؽw���Y�\�����u��a��*
�Acw&���LI��Z���ܦ� ��L*e������:����pƖ-2�z��g�����jy_|1ι�\d�#jNN�����x���%�m�d{�$�_(�;�~
_y�;X�t��Qo���8�T��{����	#y�ڨ�;x�����*^ض[ƥRUH�i��iW�zUx�x��ލ�B����@��������L �n���_�%<}|/�\����Z_f��t�)�c� �Jۖ ��Н�x��n�j����+KR��ZmVZ���Ǳ�E��}ӇgQ_�l�By�ːݶ� �N���hdKV��rh�J*�E���- %p���Dt��1Lm8]t�J�#��>'T�ׯ]���?_�˯���C���`��؉̠K�;�X� ���;%T�pS�.��%��=��;������{^�	b��~��_}�-���_��F���0~:�1���X@ЍO�A��F���\<ifV���Jj )��8�&��sq��c�d��.
��8��,4�i ������>��s=�G7a�ƇM|\��#�F�]���u�ͬ���r�nD���:�8L.��a˗��:�Y�����X��u0Q6����e�&�uFÌz�WP�6U�'g�J�$�aMM�)k���6e��6V���������(�U5MMLh�Z���L�e���b-XF�t��J>���2C��N�/S���6: �Fž��c����ۿ�1Y�dL��Ǎ�Fn��{�~��3I3�����~4s�te�t��N���[oƭ�|�ʎvH��
%'C31�@R�@��#4���qP�2p�\P�-�4�3�T�(@��z|?PN,�f��APYz�̻te����=�y�)���� �d�ʸ钼b.��\���0 ������u�쵫 y���hU ��x�݁�߫!o4����t@��1v@��yRfT7\I#��?�(0>����v���g4�#�ۯϫH���:�!ȟs���ʯ/�J}��D�}�Q�&4����S�a ��(0P�8'Dz��K�N�S������7�ac�kr2U���M��B�!\OtD+�'�(���92��xuNk�A�@��di^��Y@1��G�*�&��e�5d�S%,��D���s4�����J��܇�D��y���M�����Eш�`,�d��ϑ�[ Y�y�9;$�Plߧd���0s�{�'P�z��"V��15���׶���>���W^�X1���Ә>t��%TfN Qj"٢�F[8ڍ*�e��ʋ�O}��|�~��������O��f�D��wގ_��wcl�<�����#>����XZ^m��O<��{�o��?�	\y�U��#�೟�,^پ+��5�j���?��n9n���ĥ'��}߰a�z�(O>:��$n��v�灟�کժ$=��G��7��NW_uν�\іFWM����L<���	�Y�J�lͧ��yf'��K�����4�1,,̡ߨ�]������IRڷ!Zѓ��ğ�ŗ��+��ɏK�V�"�c�C	S�
��O~��&�%�"-v�e�\�,�0^��r^p|Ȭ��V̄v[�ȕ��l��g�K������m�&�Zuʠ�M� 14���g�Cme�҂��v�$���%������m{��cOb�΃(��Dvl�U�왒.��g��h�!Ms�P�	G�����zp��>���Od�%ݻ0�����4� k��g�*��p�ƍ�2�����=J��8/4�Km�8��W4���R����T����Ҕ�O���ۯ��g>�3;�g�O��j@��/|����_��j'�9�j�(���^��^�l�챔�3�~������ll8W�s6Κ��Y��0��c�h
�\Z��&K���m`�t_��K���z�uh��$�:-��iЮ��0�|��L���6YPE���fO�C�Rs��߹�v���9V������2ҁ��" �9:V������R��0o�.���Ln��	<lr�c1��Rf(mS�P���byyI��f�9��U^^�ѣGU����f�ɚ�,�qm�;��S���>R�"6�s��0�RQ��l3sG�c׎�8qh?:���ǆM�AF�u� �����Pc9�e'	ތ���6И2нfɉQ\s���]�`!��ieJH��¡n8է"�˦3 ��:_9H,�(l��r����I�<�;�6����XB�CR�K��Zm�2��fU���?�A�Iy������V)Se󂊗�zB���G�P�C��ep�s�3IP����8�{@�����t�8m�k�E� v���e޼7@�$
�"����aC�1�5�Gʹ ������(EI���+
�e2(&↯�V1���O4C�A������B��&��ow�>5X:5p�Q���j�1��(���q��kX+[�4@�3��W�zj@��j�(�VU�����H��kũr�@%��8e��q`@`s�+�ޫcS#�L�����A`'*6�Cp�Lh�k5:7< �ߙ��9�<��l�!f��}���0���f�mmY`�ʳ���c� Fe����@M��p�y�KRD�����V�fѪ� ��a��8���Î�{U=�.���u�`��,i,٤�U��[n������+/F>C��£�{��7�=�����$�o܀�o�o���ذnV��ٗFi��cǎ)�$3�LJ&[�#X\���̌��;v�3��/��:�̳���_�2~����}&ɲ��4g[��<cyF���� �c�&Y��HqPae␉@j�s���"<R(���~7���2�����=�o|��׾�*\��K0�j�\^��Ջ��J!G`�N��jb�VA��D7��+;��G~�c�5 E���Q[:�{����D.M����N���g��M<��6��ZV:8?�.��8�x�����x�[n�!)�ʲ�TA)�1R,�ݭ�a��kC��������s��~�H�%=�� I�0���2�i,��JJB�j_}%9S���O�+䙡߫#�ĪH2��**�j���W���^܁t��$�0X�̤�S Z�F��KaJn�-�,2Y��K,d���"��i�q$ؐ�/������*�E��4/�	|O
6��W��L����g#�Jj���?�D1U�̿KL�^�~�'3�����>�[�ۮ������O5 ��_��m��Ͼ�߫�������Et�P�!�2 ��8�+�*E-[�/v�j
I$q֚���s��3N���ǑC#��X;��n"�F,�Cs����
����d� �U��vYv�/��� ��� ���уd3��i�F�)�q:�$bH�A30�1�W��!�[镁��5��R��Y�u繰:���k��o��r���D�Y	���H���P�::��s_�r�t�t$cciJ��_�W�13�߳R$f����N߂����<��΢��e~Dz�ˋK8�w?�Duz���k��C[�h��t �2C��@M��c����p4�Jŷ�N��x��A9$�
"��6���8<� $jhl��>_5������V��������FHPU��5��?��#i��.���U|�6�5Yʠ�������!��{�4�FA�'@����x�L�R���6nZ�oQv��sY��@�q
���A��5���Y?�ڽ�� (Z5��d0���K�Q�@�w��C��l�2d s��������W
N��H�p��-9}j�^��F�o4p����>5@8���!j�ʪ��#.���::_df�(��E�y?�E�	�i�)�a�f����������SA�n�}�g��e��2��������3�ȩ���3H�^�jw�<�ml#	�NV�@Pk�~����^���x���l�9�q���P��6�l��l6{�Ê%N�i�;� �ԜhuAUK�JUR">���o$&�d���6�ƥ�;��MbiyϽ�"���/���J���*��>R��f�H��@i�J#�$��v|����9�&n8���Wv����⩧_�=�4즛n�u�^���	�v�Ԩ�9�V73���14�5,/̣R)	̳y���4�;�|�=���>[�����������ܟ{�y{#~+'���)��s�&V.���l٢����Ǳ#3�t{z���~��~��{�������'�͇���٣���p�%a5��2��!�}�aO�,�f���[��M��m��`�+�Qa��0&@�����#�p㕯�o��b���{:�_�q_�ƣx~�~L�߂M�O7�g����,����߀���Ez��Ѩ��s�N�ܵ[~���}�}�/����D�A ߗ�f�F�\S�Ne������?L^��������Yk��i��D�K+JQ���hk֌�-��%�b�V	�^xa����aǮr�m1�O���W��=DK�cC�O_�$:!1L���/'TBZ�>���j�@�/Ic��9ؘL|H*�Щ����Y%E�>�{M��z*�Z�%H5�A8�ҴlIc�R���elX����o��c����v����5?Հ���������x��k�����-�p�xqvM��S��^t�we�F��FS�\v�x�-w଍�@��L���C����d�^{f���ן��?���$�����]�ͥ�Z<�m[��c���"� D�%�f_Bْ���Є��o@�2~��!�H); �0�c _.��;���3C�AzƸ��`��V"d9���.ҬC-��O�]sP��շ�Х�k����!���@@�2T�2E�t^�i쌳����s�����ѥ,�$�h�Z��w@��ʡ=��,H�Q��9[u%��+�
�"�H�Ǒn�$�7��w݁�'�u��.�j�sީ�{���c�C]+�Ԩ��+Þ
f"d�R7ڇ2�p빆��3�
�(7�  ��;�!
�¢��0MRM�����@�����4ό(xd@�>�< pz��U�+'N)jQ���6��s�nr���Q0����K̖m5�|n>���xM:=��(�M��Yց��7|��/�JD��6^��u�o�ωr�}O
���澃]+��~O��;h�&��(��o��`�5�c�:"��@��U�h0��g�i�T=-rW&:����`�1�r|?�fW]������Զ��zF��دك�`�5x��0�����O}>����ܪs�U"(��``�r�.��M��R1:�+`��f0H� �`?T'}.�\�3����{�|�_��<��~���  ��+���雯Y���g�7M�ȍ�ڦ�����i	�,p�y[�n�(N�ž}{D� (�Ek��kH�Sȧr3��Z�t    IDAT� �W�vr���{��<�͛֠Q[�<{��}������S��x�&�q�m����5����@i�a�RT2%������L2!v��4f�u��� �?�B�#����{��ź�p뭷J�����ضm�*�sn���q�
��ä���C(���7��Գp� }�Q��}� �Haw�}7��]8�s�4���g���������w7nZ���:��1t	4��1)�P���X =zz���v�s�B'WDfbR�k��,�O�������p��	5p�Zm<���x�k���
�cSX�q������+�X�=��.9z�;0UL!'� )@ֿ��3�<�/~�a<���ba\q�e�*󋀟ϙ��O��I.k=��{��߾�Y"ǒR���u���F�䛰ē�<�V�����j8���x�}w��ֳ.-�E����K���<�;��!�#�x"-�F�&cY]dRMUaJʃ)i�(���Ͷ�_���L
�d6�'e<�,165E�3�juT�a%3�U�|"ڣ'D?�$��3�>2�d�Z��:�]3ɪ>q��b�T�{��y�����b�����������?�dV�]�MFZT�P@@�8�G�H�bH�M;t�%el�"�,U���D��y6�{�}�`˨�&��&�9;HX����(�c�9]�C_}Om;&���Ȅ@�D.�3�F�_>�g��U���P?��<F�A�;P',�o ��ތ��{�TB�fǔ 0�Ճ�5'4f�c��.��	`�z|��\��('�2������N�XS�M,������� ���T1��A�Ar��1��͸���q��߈݇���)��l�f�1�� �oͣ�U��i6s|��7ʋ}ȸ�L2Aڇ^EP:P�1�:���T�bt�Z9_���<qL	�ȫ-A�;�3�����A�]Sh>#���L�� R����,��@M�Cv 2X�sH�zP0��ٚ�]�}��8�Ual����$y]!S�xs|4�6u�-dQ}����>�� U�@$B�1'�a��d-$�Dk�fzO��CE�(�q�س�|��=�qp����D�c�C*հ������q�P��"��r9�A3�Шˁ�_�v��<�*#���f����=(����Ų�C�S����� �:�'��̫a�8�X0�C��l�R��v~]���x����P�T��*��k�g{�'<�����R݆{�p^�ar��3>X�S�!��̽χ@�q�Qh����2�2�҇�������>��5����)(N�C�P�փj�N��q"PH����)z���(�\�9����>zᔀni���%���,�K}���Z���rh�*�B!C�_*G5Р�L������߆�gp�����Xc�ϼ���~[�D"�ӷl��o�7�|��b���۷++K��z�tZ�f�#9�����;3s���R��C����zTjU|��_����.�M�6�n��wީg�}�>��>���s�߇N��1�x�����O�Qk��nP��Aݭ���#��DPx��W����4Z����x��#�
I�@8�Mg���5���Q��$R�2��肜F;�Fi�Y�������}�gދ��Q]^Be7\r~��������(5[��_���=�^B'Y@:�S���Rr�{�E�v��/>�^�M �i!�ëx���?ܪ���uk%��*��,-
�z���F�$r�5�ù���������sa�@�b�#V��F'0�&�5�3Pe@������b�������y����\�blt�y�%|����g�َv�=�Eyh0@pO��{3��>AsGa�OA{��w��GTF� Y�CI6 �G'�Gn�&7nD'������5���Ń^�G��b��UM��k�*����=�k�	u��HJ�l�T��Z��������k����������Z!��?�ʻ���_�#�W�[�uNN��Rn���<zq��1��I$�%�֑��q��V��L?�D���#cxÅ��;���7�6u��@&c�G��N,�Z?��;��W���W����Bnb�ZW���i$�X�8�~�˘��,ОE<a����h02 ?�[w�@��3���X2���٬�P~�9 ��+Yv�XDS���#Enz�ܒ�c���5� �@f��>�N�Z@�_V�7#_��$�5�l�D$��T2�"��32���|&n���;�B�6}L:��zWҩ#�"f�ƞ�_@{��1�RU]8�e e�  ( ��x&ۮ��:J~���DM6��ȯ���܀7��V,�ۘY��l��?Z����+�^��$�7 Y���V��X� �@���h`ͫC?�( s�t*����!�j��s, P�},�d� ��B��%|�(4,�FmJ*2CB�fꐣ(�3�N4hg�������A��ݰ�ҞϏ�`B���*<�ςF��z<��`G��eC=H���{*�gN|z&I��H� ��v���O���p��P˟E�~���:\�3:tQP��G�<�9����ީ�= �A}'��>�B����D�B��d��5��|9�3��r��,�;Ѡ����cjOC#?�N��z��v���U3�D�<�(ষKt�G�D� �7'm�<�T��u}R�	}8�Ӈl^���S�����y��(��&L���Y3�)v	�g��7Wp�IR����oŀ�j���eu:z�C����i�
	��d�d��*�������s�����2���Ld�oT����8s}I�6ԗס1����ӋI�������2����|�C?�׽�l�����O��O��o��Kg���M7݄t.+jΎ�v�q�X�cRY�"Z�:F�yL�E����٣ؾ������>���{1�<��~���Cj<f� �D��G��׿�������ʆ?��������C�j��׽�BI�~经((au`|b��{/.��lݺ���K�teig�}>��K\��+1�Mb�3OcǓO"Ѩ#�
�X�y2cy$ٷ��{.)2�4'�JS�&�^��r/����S��ӻ�a���Ǚ��N�^w]s9>���cj$�t,��fS����l}~R�	ĲY�Z�u)��c-��|+>���ጩ�<Z;<x�������C�I�݄hT��F�����U_��J����TVA ��q:����)|�Fq�6>�j�� X����ZKKh4˸�����1\x�vf%Rx�����|�4�1d�􇠐��2��M%�e2'���Q݉XM��K��\��1����8�6��������g3X�k4{xz�)ٞB1�U@@�$bVU��+��� ���įg0A)}:=s�m��~"�����c��*��W��������ȯZ#6N��B,͛1��d7�d;����5��]�Ѩ.����N���#���+��{ގ�]�3�Iv��s.Ymm�1R9�����ކǞ;�fb��I�i���҈�g�����kO�@��d�"=r��Z�V:2��J����C��G�c�gSoD��E(�{m�J>޻�	����%(eH�P��>�t;�NV��I����Б�d@a�;�&���nh��� ������p���̎�.��o~;�S���14{��N�Yk#�Ob����
�l@j3jg�BG��F�(��}Eb58i�ׁ�������U�^�����+n���|�YgQ�,�vW`�,��}�T7 �Ҏ�6�5{,Ȱ��x��2�N* e��P.�S�V� ���#Vg�	��ß���U$(w�ʎ�T�O��D���cm���H�|�~iJʒv�5�7��f\j<��|�!�Mm<f� e 6O�]t}�9<>|xP=|���@l Lp����3`95X��d@�2��#���F�՝\�����:Z0O��]!�<8P\[h��VB���i4x�=G?o0�O1�6�?j�\�d���Y��Pɇ�K@ƿ�L�����ѨL�`lN�/E+7�����{�0��+K|=f(V��33�Qےc�Y��qp&�L��Lx�3��t�����q�̒�d1c�J*��ӽ�[����U���t:��O�
�w�^{-��������]#�Ҩ"�3H�̪~jj�>��zUЮ�4X8j'�25.�JVX@�	>O7:��)n��� ]A����[�;R'8^r��T�Uh-ZȀ���W��|�`�N�ҟG��P,Wq���\�z���u��)Ṣ���d�9��_U2����EN�.Q�U��\S��Z�޻��W1z�Gd!�WEl���}Uj��-����a�d�������	�t�|TJy��܀���	'�{ל�s���9�H��k�nt��#A$��T�l �N��%�h8  �(��?Ћ�;�������k�b<=.�G{===�D�׾�5,^�X�¯~�+����_�"�;�8��������_$��+V�����[���Ѓ�n݊Gz��vJ�d�����?a������FT�i���(9aVx�x�MR%�x��â��^2��p�qo�]�;�a����^�K����u�����.����`֤���+7�A �
O8��"�{�Tp�-Kq�mK��T+d����bՆH�3�`�<b����� �=W"��r�פ�ڥ�ւ��|���L&EU�!���"?���k�����l��@�r��	Dc!,^r)l�P�x�o޺|�q���*�������Kv����d �s� �hT�^��]���Lܫdo��H�xc��
��*���h�<��68=Ke��'ஹ�Y��6zZxi�V��А�Q��C���[j��y������NJ�k��V�娿����\����s�~��}�W����n��3/��+�����i��\)'%�/�2�Q�F!/0�4�u�ȍ����D�\x��Xv��8��)Bw:9�������ۋ��*i+�X} yW3�Q6���wU�����+@` Uh�R%�GF���V���SM@j�-I9�l/�&��d��c��v�QYm�UL��d\ܔ��r3��]Ӻ�: ��`�������A��,IP�4)�QPj4��!3�J�RY�k��
�5o�f/�9��@���:2���ɷ+Q,<x=�w�<6���=���P@��S��K��-�𡀠�I�M�T��8����8g�G1R)�o|�^r�`��κ��__���m���ޘ�Ӂ/��)`U���j��'P�CY�͋v:H%ʪpX�E� L�O]c�+U�(\(5(�3�))熋�Z|r-��R=J�}}I��W�%��AޤZ�n�|�Fŀ���N��+��t���fإ��5Vp�*Qz�KY�J������P���<�:x���d��b��|X�h+ A��E���{t0Ը6 ��{p��[�Ff�O�� :��k�)c|�M��'�@&�{�;1�n]��c/@��l��<4�k�wx��
��@_o]������i�_��J���� X���."=�d�mFc��?���'��_'��z�B˞ښ��c-9_+��xu�������ӨR��(J��5�H7^�5�����\v@ '��3�iY%:N�ǩqm �v5�կ���l�u}��n9������y�<$�U*�P>A�w��Ê'����]�������\��+�-�;R�aҧ�jW,�������.����8�ϟ!��|�5�7�'?�� �b����sp��c�W�unڴ[�o@��@�P�����p$���(�(16���^�4�qߧ����\�t>�g�}<���k ��o|Cz	,<� �����z*~�_`�Ν��cWJ���^��M��6�1"p��Ǯ��o���}N�H��L�6�����K.z�xzw��009A>��X&���Pe'�o�y�ۭ�G�~S�>[`ˁ^��Ѕ������ħ�#�A�Z���NÏ�~/BL`:�(V��[����=�������U��������.�Zb�3I�Y��?�4v���{7�i��T�������z=�I�ȿ�
���TH��d���ߺ����W�8�:�����p	��N,��r�t�M�:m� ���y�������|�U���R���%�g|}6���Y��Ĭ�QOȩ`E12h�V�(�!��j\����55���"�/�wL  ���O�F��U�Y��V	����"�XƤ\��ZH�3eP�jI�҅�0s	c����nX���|避؞�W���'ox��Q��)�U��Q,唙�u�~	:�.?���,�.��ƙ�,��o�����Ͼ��z��fܴ�:�y�	E����6f"D����@?���> �߁`�$x|�*��LTG���1е0��j
^3@t�k����Yge�1��h�i��q��R��8���	�l�l���t(�-�|���RK�D���
��Ck�.9�+e�d����b�%�*�j�%����"�d3�� Ȭ���{/jUf�0��'M��-��S�E��(��2�57<Uj�
�{п��p?PʢZai������}@ͷFFU�<�B`s��f�PY8nf��&�}٥bL6\�c_o�,`v��cQ�dY�2��iJ����jʑ��j-�a��4�lxSp�r+5�b(S�x8,Q�(��"b���]�|��;8͍BaQ�S6�{��E�M�C0���(Lѱ�(1F7MQȨ2��+Y��)��x�񘌍Ȳr<,�7�f���
f%��Z��J�˪ZsG^��1+��փ�������4��h�����B ��j�Q�xk�}퍀ٚ?�JX�9z�����U��D����������=�����q(5��9�Ϩ?���֞��_O�c�ԃ�z���~]-��'ip��Ms��[�Z8'8���l5��e�Ys����كi;�Ҵ<i@�9>�"V����6`��]�ܒ�U�~��9$�y��A+��ԥ��`X�[{@>�����?D']W��ϊ��%GZ�~��2&�S��� E��,�:���fz���ԥRQ����R>g'3fb�}��v!��'��i�$���?��
E��Ѓ���QB4���g?��fu�E�
8�z��: `r��s2���j\t�G�Eq��A᷏���μ2�T�C�nʚ�rH%ƑI'1�Ak<��}������eĘ���;<xPѿ�n|��O�ꫯ�[��!�a��?�y�~�i��~����ᮻ���)���/HǊ4����J���.|��JɀS1��	���q�E���`|�z��@��)��e�N���w�z������_��C(:C�NcKW/��;�!�����#���(�#g�����/��>Nd��f~��3�`c�Tl|�y�A|l��Rˮ�_��.�3�ٹ��>���%�񩠟 ����cLDi0�ְ�����/ �� g�%.�J��I�]Ȓ~�X�\yv�K���4*Il�Fc`tlC���5Eq�����n�/���_X��>:N�vQ)��U�7��䭗�¦)�A#�DJ��D�uR�]K¨vT�v�ܤ��u������� i?<�)s��Q3�(�0R��}2&��uIs��,��, Q2c��A�!�RY��Ҝ�-+n����|w�G��>���?�� A�Vs�����7V��g'y|�CQ�����Xn_�P\$/K���*:[��?��]��ډ�^�=���E^�s�>nO�	�jSE�7ǃ\�����6�5�@t�m�u��7\+�[H�k�k�۵0��d�vS�F����[<v+X��͍�j��MqCU�j0��Bu�ˡ#\�n�$�޿��ZN�܀ٻ,w��O����>,�e^*�=>�k&}�45^���X}��ұd�9�ep�PU�
U63��Pv"�6�^�ϸ =c)�$�֜����?��{Q� A� �, i���I�����{4�Ҋ;XEa�������«c��a�Cp[Mu,9K���"�@��	7$]W�؍C��oVah�N Ţ@0��~U5{K#�ڨ�Z�`M�(Z���a%�h�F� ��}�V9UKd�t9��P(�I�Df    IDAT�����z�Nd3���!�~�wO�� �5R�y�(�k�7�W:�E"�B�U�	ʫRM��V1kX���X��=8�gz�j��[�q�s�r����1�;���W|�H ���{@�N��uP��5���A�$�@U��s#���^{�� ��@�׫	{ n_�����?ĩX���'�����/���0�wZo���+-|U�8X���qB���fl+)R�UUm�	�|2�Vf����*�!���@�}��sU�_�q�ԁ�'�C�-j�l綀_z���P��*����x��ړ�E�.K.���]>'=a�>d(�&��#� �ڣ��5��@ɾ���\�CQ
u5�TF���h��*A�Z�@4�G��,��0�������2p�3}.="J4'̞��p�x����"
J&�F	꺻ੰ��D���γ�|��7]>}�-؟��٪6�{��6o�-�Y4ބ��='�r2::'I¤����I�����8.�!`��b>�B.���~�~|�_�m�nA&��O<����[��*���=��ƫ������{���`������?��N<E ��W����ҥK�5^ye�z�-�����M�$���?�1.8�\8k�ݍm���,a��$S�H����� )"f�N��"��/ol�%'�ŪM]�O�P�z����fQ�&�����ӿ�Z�!E�\���l�o|�v@ �5NRZ=H�F�p�W�s��/�8�s֬|�w�s�*��ʦ4�O��9�󌒡�՛f-�^�Y%�a�����)�����x<���ף̹�$IfQ�t���( ̴S��R-a��.��������;k�n��o�޾ax�ax=a��&�$J�ʭ�C�ٌT���|m&Ԍ2���E��JY�+��ǂ"[����O(��ˇb�	�/'�_�PLOG��(R�#��M4�(��L���h��y�,*m��/J��Q����ӘN͉���������+�]�7^ٷ���G޼��U�E:N<nfN�@G<��#G�f�&���C0ގ`s̪R_�|���h��pڱs���+����ޝ�E�w��yp{x�J�qp3��4sD�:0^p��]xm�TB�j� >��(Ù����qd�@qHz�Ϊ��۠��;����!�(M�ϭ,�ެE\h
00BR�R�ꐘPn�9�*	o�����i%��fXI��5�������O�TFu���C,��\d�6�*�#t�-W�(�0�"��+Nۦ��EK0���e��I�_�B��1����^���
=*��eH�ҢB|8 �@�?f�(C�6s�������A�� j��fa��Z�@��2հ�SYt�=X��x����Q�KƝz�4na���q)�9q���HT�g�^5�|�f�Q���9:��k�ӓ�X.#�ɠd$����)�*7BQ�`��ʬNΨ�����21�d����L���`t,�\� 1��73 ��'�,k�'˔���@'�����������u�&A��a�����gR��T��%��ց��\�k�_
,��2���	���; п�kک$�5[7�kd�u���uMg����RY6@Ŀ�4�~�r��P���������_g����@L�^��4�H:8�����o�@�xJ��
���\�ʺ�Z�F�%f
?����B�]7�|nT*��eF�� k�6�,t
H����jݙ2���S�M��phpD�#~�:�1�kTӃ���ާ�X����O���3K9A+���j씲����J�ݿ��fS�\��;�{��y6�UʤY�~.'{�hԙK!�sbfG3zvm�;/��R:���	�)�i�����V� ��f ��H�\ɦ{p��%H����^�f� 6�kio�9瞋�O;U�ž�~��Cɴd���cB��B>�Z��������� B~7���/��;nE�P@��?>(�|f�ٰJE!��Ħb��g>��s�Y��O�m[�J/�H�='0����q���Ϗ>���$DBQ���1Q���~�s�:S��=;v�������~�%ǐȤ���2�]vB!�97ʦ4��H/Gk�O���,}��8C�NGP,��2Xr�����,���L�xk=����iW�M�t�Da���иo��j�{��?���~ ���QI�Q��lio�`�
JvY�I�&	0H&SG�x�5%=/����Z���I��V%��%+��t�kX<Xݲ(�����SV�Y�Y��s�4$SY�B2����W*=J�z�+fQf�i"��6�������rtKvx���Au�LN������<�n7|��V���n?��fF���F�v���$�N��l��"�&�r�Y�
�8]�`�Y�I��@`%�+%T�bg���;�^���q�A�������*o���ɧ�}o���O�:e�ҫ.�9�����#��x��W��K�a$k"��	_�N���t��ᦏ]��O>A���n�X��υH$$��	����i�T��(^z��W�E��O�^�M��P��al{o9l~W��U3�Q��^�ֿ���dL,@�!J<�T�]p�C����`�����2C�HE%C��{��'�������$�l�ڈ�"���鑅��H,�q��ʬ52y�uZ�D�-�e^��U�N&\0��iL�r��s�iM�+��	w�g,Z��g���\	�C	Y1�v�U���ې:r ������O�)�����k?`��Ԇ&R�8���@���RC��ٸ��+p�%��pz�^�ʎi� �iK6��u��i� ��l�ͤq��"҂X�Q41f�yؕ�m]���u"���Sc@�I��r82�GWSf%x����"�OQzJ�7*������P��@�IFܡ�M[Ϋ9�U�J�T����8� @�	��	I�t##cU�bYmX�>0б4�	
���%Z7�����_C�@rBSl=Pѽ2��A�~}�l:(�5��ve|� K��`\*D��^Y|إV�"��NS+��E=X�SI{f]��6@�_S�7);���ؒ�����v�Q}p��������0����-�Dm�:;��]�� {Q�^ �F��Q�T�t2�}S��
�
x�I��9 {�~���[��AA}|m=/���ڡXUt�c��V�'�Ru�c��T��Y}V^�)IP��$`j�����؛�uŉAw}��rҶ�����7���+@ ���\˸[�
\'�[��&]!_,�k�����
���R9�������s��6D��صqV��U�@K[��f��,+e@�b>�a��� G16����8|�7c�����y97n؎��a��D�b�ٸ�+p'bd|Lh>�Cê����O�+��hXV��J�A:���� �c�s�(�=��3Bb�����Y�믿^�~��Ș}�K_��\( a��}���K����}� ��;＃-[�Icm&��ף��	'�����I'/g��[��Ï`����Lb\��Ц�f��O�4Ebf�墘��q4w�Ĕi��:�ؓ/��U��|g$*��ύ��_��v��J���������G�����ʣ�L)O#�֖ ��Z,Y|���`ӆ�8rp?��	�Vz��?�뢚�CZ��129�Ƿ�G�=�	IVx�-� ������r�հ���auB*%5�L�[�:>�R��|IL�(��~��Q�Q�	%�Ru��c�
��Y��ǃc������>�T���Wr�"�C��~&}�(���]1ӈD�h��.�d�be����H<Uf`ON���IB:��=�t^�,F�*=�T���fe��.6���誰�{h&Y�����m�_����rɡ�������翽�`��ϼ��u��|f����Z�g/섗m�`��#x���x��5�𶰑�}���_�#���S��ߝ>N�7c#9$F�Q!�M@���d��)�%"��mƋo��+�u��i�/��ׅ�p�t�-�c��+p`�{�����*c25�U�r+N+7V�|��v�ߑ)^w�e������o�f4�N(�����UF�jF4+2ai�!lf 5��jb�����L��+��L�>5��C@�� �ڞA��:$xh�,]~�x8I}p{"˚���p�Gc�	�b�TA�H�q��cGz�g�z����:�Q���/��L�9ĭ�hq�~>^�ਚ��sJ%�3�oX�c/8�G1�O�Iy��H2u6@ wͪ��hP��M��ۉB>�1N�ba��Q���ϋ&�4�QA����:puÔ� lim�8M����L+J�HX��,�$�A�BU`��h��l�"1�п�eNQ{����/�	|.��.:C��=����a<��Y
7U�3�l��:`T�dQ)�/��Fy�e��IO�ζ���ؿ�2��^C*�Q҇�����C���xu0�0�A���u��R�d�G+��}M�D�T��mu���C]�=��t[����?�y���~,����d?|�ﭯ��]�1���"�kBe^Z@Z��x�J7dn��^�p�5�y��Yb�C`4 ���r̭_UŬy��cC=o��n͟��C} ��n.�Y�w��w���Pn�j���-I�?�e─�k��P�!���%趚�� �~�4���bq�sR��b�I�QsX�U:A��b¡PR���r���U>�T�t�@�a�>��T�h���`צ�X����pҸ�aɘ���V /+�Lʹ�jʹ�����7.��_��s�
e�{�ͻ����ﾷZ�=�Y�P��d��Kf<�h��J�⪋n��~J��Q*d�}���тo~�����[�
��/��_�R����s?s�g����_��ג����{�t�� F�G0}�4�ٻWn�L��o�Q��h�@���;�m�����:?��O�p�B�6oX��<� vlۂh8�`$��i _*� 	��i�%�TvT���BЍpS+:&�@g�10�n<��r���:�er�����޻o§��Șe������g�޺]p�C2ߙ�b���]ÔIq�p��wL'܉m�ס��!�p������$1F0���<aҋ�#�y�*괽z,�y<�ċՁ���Jn�sK�N�1�C'�����v��B9G��ߏl�pxι�aQ�48�I]*�P)1{��q��8����IY������Y�Q�{���#�(�N����p�[Q���c7���/�k�?�r�t/�kR.���s���cf �ǻo������R#�"�I2I(�"=���T�#���L'�g�?}�͋��ͫ.8��9?>��
���G��?~}���?餓&}�֥8n�4��GJ���=C������]B-��QǸZF�WFGS �[#8���p�E�%BϐڨPE �c����P���A��E^<�����TB���uH��z����k��{��8��} ӯ�Ni�W%��,��Z�Q�����+����,lцt����X\up2�X��1�:_NX6�����a]l&�ld��\�L2�&Q<�j��4��c
��4�t#}EQx��"�E��a+�]�d ��uP�߇@�	Y�	_Kλ�*�Ι�d���q.�b��pa�o��|�ܡ����D�ʋ���?+A#0PJHbe�Z�?�@��y��0/�<{6���F�p�Y�=x�R�sK���&Hj�x��r�HM������(_+��
�
\�T�v�L���>tv�#�Ju �UyQ����O�����ٜ4R�Q*�����8F��DLwLVg����H&�+d�lnmJ�E�.(�l*��`PʋMC���� Z�!�7�X�����*/ Q����ټ��M�p�/�\�2���|e�@WQ��ݟ6�B��VO��u&��_F�̬����������ZʖA�q���� �*�%�81h�5J���j�r� ����:e�[��4`�r~s�Y���v0���b\(n�<dT��末D��۳=P�`V(� 3�{�Ħ��:3��ف�=p�vB�+��"����5�~�a�,�}ph5�r���F�7UD��}:�mץ �RR��zgl��-M閷�����P��	r�j26�*���%_k��=�A�
���ʒ6#�f/�Mq�I7\�L��w��2�5/���#U���h�Q=�u�w" ��%Vy�{<��u�=e����5,>���r��T�.c;�+Wv����3�a鱂Y@{S�7��lĚ��B!�<n��@R!��v�^6�^ǆ��p��W��eWa�V	�X9ٺe7��?��W����9s�aѢE8��p��A���!��	��X2��e��l�cE�	&�JH'�̩�����m�n`������glݾ]UYP����.�{v��K/�$Ypҁ��n���U��ob�ʕx�wd��OA$��0:<�U�Vᙧ�@��z�g�'?�	N:�$��|�������P7���e<H��2�pϘ:M�T.rF���D[:Q��1:X��o�ƁC}�DH�,#�M`ʤ|�s���[���m��pa<_��o����}�v+sS�M!�W賊��(.��"����o�6l۴���ړ�M�4V�MQL�2Y��6�2��h�ƵL@ �SK�G�ΐ��j�[�J(���b��E�X�*��$˔��H{�z���*�s�J"��{P��T,��Dt�dT���+���罠x}jd��L�7��5,��b�"4~�l"\��xg�&<��cش��
��5�ri�
c�����/��>'�\��=���Y�5��|�K� �ES؋�o���l2y<���b�F��J@��x�%�I)j��H#9����~�*j�Lv������oc��D����" �����-������={f�e矅k/�Ӣ^���\e�7m�����AlܸcT�-��!q#�ᄉc���������Y��1�0�����Ǡ��B�@���ӯ��K�m��k�?�*��s �
ý8�s=ƺw �>��WL�(r�<Y\'*���S&���T�|d���/:�	Dn���I	�F ��!?���E.9LQ�	�AO36	2�N-z6��#��	���h�A�2/|tC��&�����G���������Ç�#T "G�A&V@(��׃`�+�,G�H��xq4O��ؔiwLA��Gɬ��v�Q͗л��{� �{ ����@@�t9l:���kT�le���SYMa��1�cٔ)�J��L��Spŝ7��Aw�$i�}*�^�I�l�)<�Z���G������!&�0�py�k&���!����"�<u
�Ѩ�:�BI� _��R�P�dJ>B㠜�2+  Hԥ^��2��\R%b�����}��i�����rFYއ �j{s��C�M�(p��cQi����S��G%>7_�K�����>�"\�LT.a�@�@�G**8�B�E	�SΖ�:խ� X+0IK�=���FQ�ӲiVvH{R�]%+N�t��������dS'���
+ ew��)�T/J�Y�ESat����t6!�{��=��a�r��-�L��$�N�:3S�����u�1����| ��)�O����y�d�P���A������� �hjV�e|�A���s�LY�?Ng�c��ov�%����:�ASU&��y	֩OoZ�գd���
٠�	-����x*K���̲��c�iM��2��OUV��RU��c�� 5���DSo�s�@�+��d�**�Ȋ�{�
�)���4�s�a���h��� �G�r>��-4 � J��TG/�*5�O��i@���h�[�M�����T���~�̬��g��XUD[u[^ס��u�SVBK?>���O h	���b��Uز~��4�T���Gw]1y����uLz{���%G�Ĩ�wވ�^�Y3;P6iz	t�9�o����2�ך�`>ο�"�I�Sғ��g�x*��є4}R�M� ��YܫG�N�a��)��׾�믻J����xC*]���՗��gs.���� FGǥ�{��c�,��?R8    IDAT�d
��Gp��>I ����Ta*T�IIա��e��y���_�+wܱr�����~���A	�3�������mm�2��p�\Z�^sG'�&�B2]���7bժ-�+���;2:���Zq�7�s��>WY��C�4{j|�%t���A���`�, ��i�/Fq�֮Dz|D�P�$���,	�|6#�8h��0� �i�h�J+ܬ>ə/g�j\f�KW�<T�s*+=�8��t"-��b|�
�����˓j�
!�X�I�!Ǚd�"Y.x��*�kJ�`V\F�d��5��x]�I'���K.���^�����d2a�7���݇���/b�Ɲu��B>����� #@ܿK��?�1|A�{h/��6^[�c9� J�fjUMA��e��ꏜG���{ϯxEx���\0.ʗ�DR���c^��C�q�1�>7��3��2���|���>�_��ܾ���J��W�Ҷ���z��n��鎶����8�/�;̛�	#�G�d ��a�}��]��7lŶ��H�5x�A��B(�y�B~�}�	�����`�L	��팄|�9g�Y1��b8��M��ċ��Φ��6M�7�*�-l�:�{7�F���H�'��|6�r�D9� g�/A$߁D*�Zh!kM\f;t6(�ǂ�HX�`\x�Y6�
��?J���M�Ur�<homF8LC ����B��D*�#��K���A�+(kNx��ʀQ�`�������S����`�����l��e�O�7�D���^��5�c�bF��; ��1�̠���C�D%�q�C����� �\<�7���X��hu�s�<��_�J�I���Í�I��W�%�0�C��ȍ��U�Ŕ��A�	� 
yVR ���U,�H͔9@���0i��l���5��hT�.�,�@G�I����
E�ۨ`����Ȱ4�
@c����}<\yH0���t�=�0�wQ7�5��S]e�U"�9�l`��HY�AVJ8GZ��:��-͒�Q���Q�"���àU�r&<�vdK����oh��|n8�
璃@WU�$ش���Kc��-Ҍ�z&��8:*z(�[6D˚fh� f��M�0�̡�*��	5�O�>�&7� �@2A*h�3�" �T {�V�:�b���%;�T��h�V�v�&LD�6@��'J�U�
��<�̸ζs>�y��&ݖt�r��(~l�&{�(T���Fs��q&�8'��M����С��G�_�~��[�g�嵺�l 4�Wu!Z���_a�M"Г�](��K��WX�6�"�W���`g@ =>N��֐���r.�G�,��~Z*%s(FGl�'��`��E���G��@ $f��Z.�ټ2c0�c%��t��N�)n����э�Z*Hϖ�5�f�Жs��O�y���>얊�	h�9�[�(2}�X�����M#�sP5K*o,��^�ω��^����G���^��hP�t�����L��Z�׍��Fiz&��E�YC�߅�[�c��u($Bq������T��)���2EU)��ZEzlM!�g�І�Om�(����[���[wx��y��q�1�e��9�-�� �I����bT&��l�d?�����6�����ŗ�Bѳ�?��_|c��r�/��Ĺ�Ԙ�BU���7��*s�!

�<16�b6�ϏX�>����grg���c�ꚫ0k�ll۶���a={�A���{JR��`9bʤQ��Z�v�x3��Y�@�o���>��\Q A�QC��Cs$�O|�&|峷��)�{ ��CO��|��FU��k�J�ժ���8�Dg׎-B���#?��ah�&�sR�L4�JonRB&^U�֪WL���d�%�H���R{���(煇I&H&�]Nr)IeE�����@���^�}E�n7L�zz�HU$�y�၃��e�M��f儙Ϣ���������߰��"[�b݆-X�v���H�
Ҕ�$A.�@����k�����O%��f��}x��7����0�Ax|MR���;�ُ�o�7/:բ��V��'_zc����6w�� 92"qלAIx�r�ʥ�k��@�D13�_0���;���;�Xz��N��=������]��s�����ⶥW��y�н6mێ�6�z��h�x�+�����k��s/bϑÈNj�ɯ���%Kp�i���)W�D,PZ�LDs�xQr��Փ�CϬņ=ÈN] w�YJ<:;\H��o�6TJ	̝Վ��?F��=G��uHʌ�XӦMA{{����z180,��֖v�����U�RGGN8q>�%�ɗ������=`��Nʓ��/����Tu.�f���-tV�RyZ�S�V�u�
�"kGQ���L�ç��8Q���g�w�\�_d.+
�x�U_�C�bf#
���Ș�dS�?��7<���Ad��s2;�Gs�A�#���g�6���i�CP�|( ���
��m֔��|JXV�u��-�pf��_�@hRθ�b\r�Ȗr��h�mwW���Яh�]u�Y��k�#@��`�R-	��ZGK�ڛ��-B$�Rp&W���|�9<(U*��@>�� �ĝ�� <�@��2��8f�ع���M�����l�w��b�TJ���A9 ����V�^UWl��V �9���Y*
�i����$������)�V�` �M���s��7B �MH����GG�L�EQ���( ��@����H�_]*W�Ge�"jR)�&���T���(eR8v�\̝9>���y������s�A�^��M���Q!)�K*�B���:��j޶g.e��������!Ki����Q���с���3h �Fϑ!�z����������U�;B����I���/��9�`ZsK=�1��R%�5���Ё~��c�Y��h��r�x��6��upi��`?'�VYq��ȰA���2xƩ�aHRE�)ܒ=�������g�ܩ������2��I��G���h8�p���U	u�_�����{R�����qH��Ũ�_��P-���U�dg1L�*?�
2�ŵ���(�|I}֪���a��*	��A>�JB(�.V���^����c�e���cI���������ڿׁ�}=�^�S�)�т������+ȭ�|�Y��UA��ܸ��mB��G�RQ��)��Y��\N��>x����YC:1�X��O�{��r&O���H�)����?b���ȗJ�T|�e8��D��k�.tuu�Jl�t�z{�eO���j�lp�`<1,����׾�E\z�Eb<��_�۶퐽�|}q����J�󜷸쬈*�,�����228$��'���C�&FG�Q�����ԩ�q�u���%�1::�z/��\^���E�(9^�`D�\.� m(��1�N�ǝz&Zۧṧ_���(̊Mmm�SծT@<��=w݌��w'���3�L�Ǘ������Ҥ픀�r�wV��ڄ�J�P�^��]5$�b�%U�{L�X�l�N�v-�����Y�0�6��B:Q>]�}��)�E㴢���^��!�HL��:ax*9�֦8T���9��+�e�9X�0�1���1�) ���0�� ��I�
"� ���;��1/~��o���?���0�<���8xh7I��}{�l��^�p�b����� �S��������/aWW?��XK�a��8��*ܾ�BT�V���,#�
z�Sp�È4����e?#�Ҁ�����>��5T�<������-O�v��������~�@�_^~�;k7|���t��`.�Yv#N�?�֮��>-h�K��.D{P1N��X�n=Vnڊ-{�c[ݗ�D��f�,��%X0}
��,�!?*EEGa�U� <��y���Uشo�����!���qM7�����&?,���s���ְy���׋H�E�,��0�шL��	�(�G�/1����|.#�Ķ�	�X���o�;�~����0C��**I�0|��8��X�����'�[��y�jE�јEc&�	&\x�%/d�L�������f�l�I7G^/�3o�Xp�OJI�����\�}^W �p�`X�p3%Yf�ܼ��7�� |l(����{0�{��0@�Q+؞X!�� ��:�WŪ��Nv�Hy����W�D��'_z�Tr��\X�!`ҁ��QVL�f	����P���L]�!j
�XΚ>3:ڥI�%���C=6yU04<���Q�,�pL��l���k����	U��Ě�̱J���J9@e�j�LOdL�JTV�(	(��dd,�< �$����sf;�
�3A):�Z1s�T�#aQ8��3g]�4���������T�"���Ho?zz��&h�Qq˫lӅE�#��R�� 5��
x��dl*��id�%G�������!t1�,��pρ�\���#�;_(*
؊��/�2�/��ɸY��:���k�q��	 �/�jR�L�jq�R%I(��)z�|�V�Ipf��
��z�ϪQ]e{EfN���s�L�dS��Twx�%�縋���~yH:+j?Pcbʚ�w�ĥ�g�4#�':��A�4���@I�@pV	E�cfV<]H#b���!�s�O5����'N�4w"�H���MSb��ժHp ��h�3� �R�j�[�4��ɓd���S F��|��4o@�H����jU]9�\�"��yU��,\{U�w|�rGz��X�._%Ry@[$�~�����l=��١ֵ�׊e�%������:]�2k�Y�lpBe�� ��:����go^��i�bd���a�Q�)���ǉimM9+x����k�z�{���
FU:GůGK�z&Ŏ��
�M%����Vܾ�JLj�k-�Ux��5���	��t#�70u�t,��b\{��Rڷw?���Fbd\�����'p�p�q�Џ�I���0�RsgM�7��5|l�b<��c�?p��[�k5ŭs�\7��l2Y��GV��d��6%��9���R6�G�4M&��r.2�L��ٳg�䓎�g�.�C���_{o��򹢼?�������� �bq�SH�Yxʩ�x"x���x\�XK+2���/ѐ�����L���+��C�bϞ>�L\�p�2�r�����$�xt�_\�k<ê��t��KPLO�m(�Erlx��|jr�k��U��``xhɱ�|~��T����I4EG[�P#y~3��4�c�è�I><����@*�5��Ba ��x#�d���Qz.U/��@q�Ma7��|�]��l
/��{�E�I�H�&�O�A[fSèXz�"���	p�Q���#��d�ު�x���S�2z��0sJ>y�Rܺ�"��«o��"S���HZd�]���(Վ� ��07<�(#�@�U1���p~Zg��;�_�?\vEO�\�˾���<��`���^����|��t�/�1��v+�8~.6m܄��ߢxg�s>�,Y����C,�_���C})���<�Գ���-���#�y�5X8w:�霔��V	^��>/����<�v!�1�7��LJ��!)Mze���`ΜɈ7��ylڲ#E,\x�l\�0��xXp���Bd���E�pѥ�	X(��G}زl��ln�67N4�����Z�c��n��-��p�P�-_ï��IGI��#����/��*&�QH����T��L˹�����,�H���
t�5	�yˠ>��(t��Ȧ$:�9D_e!=F�
R�#�� ��>T�Cҋ�` � �g�P�2d�Q�����/ p�T������s�"�u�E˲)6!�i��ȟE�C2�U��2��"��(�q�bzg&w4!B�B&-MI����!�A��U���p��_2��`�Q|Gr5�q��ԼH���
O<�8W����^�p�l�۫6?>_���ҙ�
0���Z#�K��)���K�K���R0�&VJ�y��Jp�JJ6�D$L��rK���R�`7��
��� ��J�is��Rf֜Ҩ%@���Ѻ�gX���4iG�Q-��q�98㤅�����B���̙�:؇M��Io���'V�fR-μP�t������:��gHu��ϩ]�>;�BT��>�9&r�	��"�;f�����˫,(ב
j-��h�3���-�xMǐ�p��Z��j VA��YT��R�:.S�G5�k�Ή�H�`#�9�T������5E0��M�); Pn2��]g��it��gd�s�0sJ;:�Z��ڄ�x��?&P�KB�=f\1`�@�,}��J�ť�#[(H�� L�6��Ύ6�����0)��@"�C"�C�H��$9
Eu?T�s�̸�HfϚ�yӧ ̽�,J?�({P<.$	�"�Z���+���{M�3���2d�
�� �,-�
ع�z���_+.i@�糞����>W5�G�/=�������#I�����E2G�>o#jc�D	�qׯ]0����h�E�`�dj&^y�Ily�=ᤇ�*;.���g.V�B4J0ƾ�\	��(�A�Tn��*�����g՚u�l�u@=�;'�y�p�g��)���Q �upP�ٯ�}HX�e�-�&�BZ������>�%�_��_<� z����^~n:���D��&�䇵�V(]��9V.	L��D"�L��S��7�GKKN=�DLg�&5!҆���#g�І|�6DV@�I�XX��fϞ��'�i�f�opO>�^|�UdrExA9S�VB>7>��[����+F��蓯�?��{��L�9�����*')�~Ҫه���@�f�y�g0�SC��Yp�yĹ+��:ø�]��>�c\�t1��>�������<�~���f����>�LS %��x��@4~SU�� �q6�N�N�3E�Je&�h��q�^#J�g���A[g���o��k����K/����_���,rE�_V%6s�L�� ����k/ǯ~�O��0��?��E�H�����Wb�� ��a��N�w筸��O=��<�

� 2e��D*"��֫Sh�NwU�L�I�e�Z١�ܔ��3�a���M����羸n����nw���ܵ�&�w�|lٴ���o�ko���g�y&�:�t?.��x���lH�
X�n#V�]���a�O���ŋ1w���
�����;dfn�n�xz�N��5g|*
�`$����Y����{C��
�{�4L�9#�$�n�B2YƩ��%�.��H#��@P酊܈�0��%�T����j�%}QaRV�~���C�&0Ţ����"k�[~�"y���S��Y?�Tr�� �<�Z˶����C�
7n�tƭ�J�f�Hg�0���j��Dx�S���Q,����]��~	�8�I��%�Z!���%��,K����h��z�@�6~UM)�HO��*k*���i@@!-��oE�ڳB@���B�"w���b�93�w�^��/<=��1�J���>(�lf6�7)EJ�&��˼U�6����ތ�������������d���b4�s6n ��ll*��R�,N�:�ESf�3�C�t���d9��Ё�q�~�1<�u����=c�a�u{<+;Z&}ǥL)�3P5U�@��J
�Ae!��,'ηP0����������}н�ZA6�G�d`,���h�DE��9�r�E���X���FD� �|��9T�)�]8n�4\xƉh	{ġ��w�-�#9��b��J o:�B�I�ZK[���u�u�!��ah�%�������M�} h�9�k* ��;lj���<]ACϚ�E���
�l��� ˣ��[ �`p��@�|\E�Q�/@��D-_L�@��(K㹮赠�G��h� 
R����YU�T*5*�j ���?�	|�
Dk�̯2��w�����Pɉ��i'�Ǽ���' b�/q���x�^/{~�B��� O���bQ-�Of\I�b�2+�����i)<TK��{�74��D�-�=�C2�.��q�8v�T����������)��I�r{ѵ��mގ��$�� <~�q�-����Q�C*P�+�i�X�ש��������O%y'����v@,�DK�@?F?G*Τ�J gɂZ�|�ƽV�9��j��$F*I��Ô��5�x�׭b�A�<�(��'�� �]�>������گ"    IDAT�G{K���2,[v%ZZ"���Z�v~����}�}������M�&Q�����T*�l�flH%2˪"G�䟣Vƥ��SO9	���êU+�u�r�$b`J�)gK����A�n���NU�cr��M.�}}����
�Զ�dM7_���H�J24�֩7��RFkk+�3���Ǵ3��q����ؾm�$���&�'+� �}w�����1<��
<��gp�w\xd�p(��9�JpddhH*�D������&̙5>�;�m�>/�E�`��P�N&�X1)[�&e|���G�1�L����E��RI<�^Rn��F8H��Z�L��	7��@.�D*���1��D�&���؅ޑ�&`P.����j�J��zǤ���#72�i�:�o|K��T���g��#O<�#}8ܤ��~��\�$n�a	����"_H�o�n���S �#����g�����{�3gM��?q��}�e���_�o��r� LwH�A�]�G�LV� ��4�)t@�F0S1���Mo�p۵��S���{Z��s�c�������xG,�;n��>[�t�x �wlCk�$��̚�������1ӧ�=�b�������9ԍ#���6�'OE����.T�q���J �Å���k��a� j�N�kn$Kx~DB!il�E�R������ǡ#�ضu7����@&3';UDڊ4�i%Eቒ��I6��`6$�-{=��g��Z��)j.6�����br;�Ò�'݈Y�!"F}�'�oa���1k��K����tbf�T�&��WndS����8MV.
RN��fP���:�J#4%�Z�j`tԀ&Ϗ�#u��b����2F�/{��l�.אG���H����àS1ui& �Vv��]��T�� ��Y4]! ���7]��?G{�B�����t	�+x��#@�'��PE$p��9�)�[����(����>�	t���t"�fi9�����2�adՀo	2�xhaZR)��(���,w(WP��<9�yr0���EM�A�
,=s�`Hh:�����5��5��\��eeKIߊPI��p���c!D54�C�%{P�eC��ՉD����dF3E���x�x��d�T���[9.�VG��8j�$�O��E矁���E���d��P�y~����Z}�Y�f08���T|O+*MX}���u]�
t5MHg��R�{A�l���r,J]4uE@�*0�@�G;)?��ld�2�:��*�4�IӨv�m���w�A� �j:���ܱ٘Mw|S�)]�ݠ����/Ҡ��|��̼W��+Ry�YM�"�jֳ�eU���$#Q^b�@jc7���0�s���لsN9���DɃ���ZIhM�B�*��"���(���
Z�Έ!���z��J�{2�L��|�Hq{�'е�G�FD�}�L�ufϘ��N���-��悋"g%��Q9�UY~>u��!7X���k6as�A$�8�Q�%����z�N��8�J����A�� �>5�Kg������h�״ =��\��!z��1�b��GQ:�uso�&i|.e����ă�ۥ�C!���U1�UMl\�>���"����D�ң�z���֖	���?2ЇΎ8��f�r��hmJe�������O~���!D�;
F�3�(���˜3|Mm�D�nV��p��=REktj.�X*�����5�d���_�ʒ.q.
����Ī/Ar&��,��=�t�� �.+��Y%3��aYdk���ğ�y�|�wM��!/$8�1�]��jFL�x��"_��402�m�wa�.����r.�b���޻o�W�Sz������X.������s	H���,�7ED��`�>���s/{�����,U9�U]����n�o	-��a�����Ѝ�����+�3f̔
_� ����	%���2�F>��x�N|�S�JZ-���ρa
�Vڝ^��ֱg�_����r-RF�@�����/s�eYy��>'�X9vW�[MNJX�B���Ì5c�,-{<W�������m��e � %�D4Bdh:wWN�N����<���%���K�?Tk�j��:g���������i4��i���:ʮɛ⏾�{��C���<���y���p��p�}Bg��U�!Ы������b�N��B���-�2�S����w��{x�����$>x�T|Ƿ����ͻ�k�5!h�<R0��'�yX2Ă��!^��k��k^��'����/�ÿ���~y8�=xr�o���?;:��D"9�p�G~W^�o��?����_BrdD!�Hid��q��x��12�~��X̬!�/!�7�h �N���P"_M�sk�Ï2��(*=7����*m����U�$��	�M>~+�iFї�? �!o2<t��"�ѐ4�Irb��/�^ (l*�۔�j��"I�{=��J�,6��/Gv-�S'�#��B.�VW��#n"���ك��A]o(�P$�T��@��E�Næ*ȖZ�$�;�4gBl�D$^;O�<u��u���tx�l�X�/䰃�Ӕ�� MK��=t���*���@a~hV�d�D=��ڐ��ҟ���l����9����@�]D'Fq���ù��j�
�;�o��ӡCw@z=42�	<زi�c�
,� n�d%�`�@O%�vׁl����euR�H����g���r�����P�ǌ�z
b~�1\b'S�gK��p�ף�c�m:���Zz9v/�-v��Pz�4��ՉV"K���JZ�0.ȼVI�����up���$�S��]����&Ć�bQP�R�|_Pf)�����h;|���̌����$?s�rsv��p��p��طm�^y�����-�Ud2�㎪�iP�B��]��S�ȕ�px86�C��σ�8S��y�,�&dژ{[��$�fraag�3�3�����=x�|�	[��3\��B(i]N��t{�>Ν�-��i״���.x-̛ރ�OA6�Jd���-r���*��!���[_O�y ���		?�}����[�G�c&6G�N�I�9�;�ض�� ��<Lg��\]�]==l��E瞅��0�lp�Ȭ��c�������溒b�H�g&26���H������>�GD�%-=A)�5��e+x��i��^����|�LN��9�v���&1u"t��¤]�D�K�^�ˤ����
y��^z�V�d�F���S��Aȟ�0�
ef��3��ƀ-�>�ٲ�}��0g��.7� ��?�$����~~���9��A�~�/�ؙ���A1
=s�K�G���HO�Y�^1v������T���a�	:?��%�>�d�Z�bq����^]��P�}�#��ǯ��H��U�<������L�,��e�٧�=�${��M#H��8AF/Hb�}�+�߃J��	�G�RB��F��|&i��2g3�V�.�Nce��s�Y���J�9���N�n�h���8%��X�~������<{�Ss�_������%j�� �ϛ	���zU�ձ��"����ib�܁�KU�>s�-����� C\�K�i|��G��;Bz��{�؈ 4�\��ଳv`n�4y.���	��E��Ԛ�,p��kbA�u�i)�\�z6֔4�NEx�{���^�{J셢�4s#W�4�v��XZ�G:��_�'\|���x���*p�1�ς<+w��l_����ڷ��Z�|�*M���T�ԁg�K�C�V1���O�����M�H�C?|�>�C,, wP�[��u:U��5|�#����Hg��������~c�q�����`?�3e|�oᙗ�C0���?�!|�}�"������ _���kN��<O��cJ�B��ĉ�'�'V�J��ժ�U�����߿�����_}��� x��顿��]��C�?���L�����} �]�Ǐ/�|�+x��P��x4�ljY��{�l�G�~?���r�DCN���BjE�{��p����h�����pa)ς��~�z�!����k�k�����p�� V�y,.���\�!0pR��~v6��#iT�*^8%ɉ� hkT���$٘M���ϡ]�� �P���B%�A����U�bi~�l^H��ba��m*p��A�`Ӗ����1��Q��E����**��z-;�#̅��Ö������Bj,��뫃e8"�::"fRzKp7/c��z���ώe�!S�x ���7�Day�ZI�v����2��k�Iov��vVG]�-����Uq���
�"e�Z��#� ��8�+qޕ�"[) [�[�W^��g�pڵj]�^��	l��pB�H��ˉd<��H��n?2�=��t�PX��u��Iu�Y 8tp��&o8�h��0����kD�4	O�YS�Оp�Ç	���������#$I*4gbgX�.[��(��@�
��3�Tʘ��C|c�@�Ϊ�N��J���2�� �brj�$q��)���d�U,7���b~��;��L���3S���̉5%������ٵ��>���0|h��h�����"�R���	V��]��j+�
��Z�֤3&'`=��y׍�4��L˔hX�LM)�d�LL��݆Y��	�*Hmؖd-��-I�v�%�UBH�d���mqL�ɭd��da��y<�h1Av�8���m̵��F´�SVW��S�KSr�"��x+q��ۿ�b��ې�����$^pҏ,�����X�����j�eMAl��o6ǈ�Nh���D��D��ÎM8��pK:�#2%DJ����3!���*%�J�~��!����,�DRe�҃L�(����p�I��_�S3�8rds+�Z�J�����8g� F�{D���Nq�@ilWa�o�^d���o�᥷�c��A���h�D�
$��p�z�p�Kj
�R���e\-?	��,ޏ�зwj��{�������01����6�݂}Nk�����]$0��{I9ɜU�Zwxa�t�o����c���x�����sϡV,��gM>� i�S2u�]NĢ%Ҕ����>��?y�JHY�'�|����
o�}J�P�zoP�B^7��_�abc���j�<�4�����Z9�v%�6	�jN8�����L
\0�X��<p��)F��:��gC�8�c�Гi��-8�5���`O���%l�gby�Q���gǜ�$�/đ[f��En nO���@4�X�� C�y�-����W,m�YX]��<����8�h���n~�gϣ�[����`~nO?�GgR�cA`�m?:⹆BgxF,^x�RA9�4)���yR�4�~�i��=1�;v��p2�fM�X�.��B��zC{��vbuy	�\��u'�굢��ս��@(�;��L_���y�C�[Ρ������l9_�QU,%���Y��� ��}7|����� �Ɲ�aa)�?*~����.R������ߺ����K�#O�P&u��W]s.��2�0�?�{�?VV��n�MW\�Ë�~�$����x��i�D��ϒ{��"z�t\^�u���('��n�b�21z�k/���}��<��_8=�߾s�_�yb�W{.Ox(���I\|�.���a|��;0���p�O�"2�(�h�0����ql��瞍�.9M'%��Z˨x�&/�t�/�<�����౧V���_EÝ@d`M��e��&����|h�+R�`'��W�<�L��f�j�Lg&��s^Ȥ�>�P��*e�t�j��*V�x��@�C&A��
fO���l�xx]/�A�p'Ǝ�`تc�x�K�!�7C�o�#شe�d�.��At�n�,汔ZC�
� �#Z�����Tpb�m@J��Qv>�H�	��7���Ǯ
9�Y�=����6������h��ͪ��88�h[����0N�2XxX�R5I��Y�7:N��LA�
�u�b�a��"8>�׾��})��,�4���	&���0.�$V�%+	�ߛ苅ߢ�*���a �l�4�ɕ�(D�%@{n�F݆$ȸHgʺ���l����7.���V0hm L���d�g�l\k�w�s`�Z��;|6L4����gI#;u���&;�:m8����k��;�F�x�ֵ�y�f�B%ݨ�Nx��ؐ84�t;�Ƒ��B���r:�t��t��1�"�u,�q��i��i�Ь��f��َ����~�=�0)lIC�X(H��K�6V38:���l	�BM��&!>����䎞T�����P;�5S�3Z�Vyg���7�p0�v�08v�ׂ�P�|�Z��r�+k&x��ҟ��yLWP*e���0�]��	1d�/���fvA �}��F����?c��F�R	�E8�{n����mw����8Xo�7.�y�R��u����<˚��i�2��Wm��k�q��ٻ&���-��o�	 #�` Q�PZ�햁wt��~��J�:���e>3�Z���o:�'OM	8=At]n�/q��N��G�TU�Iu������;5���}/�!��ŧ�<5��Y�K�C�u�7�.�_?��
Z4���k�Ju��99�#d�Rb6ɫ��%|s��?��LA`?�w�gְI�b�^��>�����ޯvqH�q�l�#�1�qR!
Z���޲бU��: �ĉ�ߋm��@��g���"�xnZ��d�<7��'�[��ݠ�L���[���?��n|/"a�|��ƳϾ�����ĉ�rq�:�q�a�[{}�Iҥ_)�9��(�Ѧ���X��f��H�Ϡ�&��>U](�'_��pN����&>)�5YD.D�W?�5E��2c9��4�,U�yk�l�A�ꬓ��=͸OYp��*l,�A�CDe�<!M��yv�M���H*n�X�iB��߾���?�����S�����?��9{�ܛ5`�����S�%��
��0/��$�ڮ��_������к( ���Q!�^�:ŧ#���_���"FFF044b�7>�r�%��ʆc��Ć$c_f-���n����o�&&&FP�t<#�U*Մ�hv8x�8�y�x�Q�/��.�ڒ�!�<s�\$�g��4:�/���q�u�A���܏;�u/�VJG��Dj�"r��
z�on�4��������O?�?�f�Sߌ[n�$�;�k��x�Q,,������]���㟽�{Ͻr�Z�P���1�/�|�)(t`x�r�(�ΗvL�?��.�q�M�v\�E��S��CC_���<���8\�`��ƍ�]��/� G�Ʒ����ȈL���$Kk�hS~�O�'v�ރ��?O��R!���l���ق�g:�r[��w{���x��+x�g�Qw&�@&H~C�dG ����l!�7� �hL��T#��

��xR��xr:3�q\X�T	�Df	�;hԊH��P/籶��J1�f�"+i�g����O���`����U�-��)-_3�m[Zӄ�h�́'�G}Ɩ���"C����ض�l�oى\���4f�WP%��f&r���w)�H�Ŀ��A�/u���a��MW�0��+�=nL4K�@�����N:�Vf	�S����*�d`F��c�9�&*a%`|~�9�}�Q��E酼H�b�%41��{�
�T>�T����g���>l���c�F���!�eV�З�iĤ��
�rzfG���H.10(��O�Y�䪺��Oԁ�r)�!�F� ��K5�[&�-�P�@/�F]�������;�C��*��@0h��� �������M7���D�Ru0�=�E#z�B����%�d���F+���HHd�Xȇ-婒�r!�/`�P9���j�H�Uu,��钿�,��Ψ��]Ă^�߽��َ���r�6�)�>7����x(��tczq��W��v�����.�Pm����5�%A!l쵓�d�ڴ��vw�.�dx#��H;Q�����Y��Q���m�s6�Cr�L��-M�䙰ҵ��n\w����^k���I��!���<�τ�k�����"y!��n���H]~~u�:̙��\���;�����B���p
,���򕁨(�� q)qbRƉ���U�̾�    IDAT����..9w��=���)���	~@�)�
*g��ȱ�Ν q^�}�2>�y�)�\vى7ŵ=�3���.��y0��cf>������BJ�?B"��[�ؿ{�}aM��$[�o��X�	&T�"������Lϼ�6ϤQ���J�*���-ʞ�zq���G C�ؾ�v#�N�m�����i������Wٯ�� ���b�1Ʋ�KC���"��ÔjmY~��Uw��m�G
NZ��6��6< ��:�6�vb�`?���}�Q�8tA�W]]q<��,���E7�.��V��l�>���w��믻� l#�;sz�<�J��j��r�n�?���=gM�%���y�1��F> %3%� &@ٿ�yEU�����j�
傰�:5�M1H/�F�#��B�((�'��������2/G�z�;u5�(�۪��RLn�4�����7�qϕ��h1��^��Orp/�H�Ӵ��`C�����4��ND��6�O�3�~
���C"���^ZƗ�~z�	�.���D�mx����`�WV�q��!���l�:�H�`�k�]@"G02�^��8�eH�l��l� �.�?�������'t�C\��!>c)5$���ra~V<������>��<�˭!�+"����GÝ�y'�����Po3V�D�Eu?����E$X�Z���@��Ͽ��o���<�G�{������p{�t�P̢V�` ������/܊R��ǟy?y����q��=|���-��QD#N�}+3J�a���]A<�ӟᡟ<��`1W�+< o *R8��fA�f�A^M��:t��\�����6z�'n��?}�#����� ��o|�^;>�����P"���m[��^��x ���P �y���@"�g�zG�~��QRJ<2`�c�G#��uW㼳v�C3'���Zp<:n/�nB�z���gq�xm� *]rt��008��4�"J�JV��pD���d++)Ʉ�{!���x�>-T��� GK�r�j�Z��%T�)8:e8�uuz=N���p�X-���hx�!���8���F>��ԤȒ1��a	�ȍ
���Ф-YrL��~��0�}7������=H�"],ci-�B��eYizeA��d��(�,!4�pJ�P�	�C��Ȑ�H�ɗ8���ZH8��Z�sKX]N��M�]͡�_3��m�auԕ K�rN�"vJ��8s:�:;2d���Mc8z�s�����	A���R�_NX4���F�ZU�||x ��`,�쵔�0�g�a�լ;����������>����h��ĵCD��{�="��I�L�y�� aN-\�-C�d�^$�Rr�ZRҾm��_S+�
~vg�A�����R�$)�´\'[2�T?)"��ČIy �pHE߇� ����V$�� ��@c�Z���љ������h Na��èXk!W�`.��4(] }~��:�譗e@6`��6�`�P?F#�Q+�R���g��S����/�e�-TIʖ�8:����"��¨T�14I;���evW�N������.6< ��X�^�M���0%� 0	H[WB�$)��aA���Y^!Llm��P�:Mn(ԤraI0*��ޱ��l!&�Xk)�j�r�d'{v�hC��@5���*�,z��-2�]iT�N�����ɀ]d�Z���}���Aŵ���p6q�{q��qD���e �u�ϥ�bȳ<��[s2��h&��L=�CC���X�Vh�%�E�������Xmcy5�7���󨷺���Lؽm �vm���8�m}���K��P)FM)�>l��fO�^<x��=��l=��PDv�	RAE����ݬ=Q���`v����(y�`c�����bcA Ȋ5��߆�B�t�ӭ��5��qz,6K��([X��k)lY�ʢ�G�Q�2A�Z���¦�$�����8}�-��4�s��Z]y�� ���Ʃ*�e��9l�:��}�pݵ�"f���B�56���x#*D	�Y�WX�T.��'�]���,��P'*�4�5�I�ku�,�
"��,�TȻ�x��W�G�P%��9�⟌/�m�<~B6i:M\y�����kd
Y�f�p�8�:����."~���Xa�Gg�����$2���H�Ơ�g>ak���Z�O�Ƈ����.�yg� �sL��Rk����-<������3�r��:q�?>1��<��,���g��U@��i4�u):�y�d����A\���h��5M$�A@Wi��ɱq�B�Ԏ�ŵz��CȤ��j��_�"���#��Q��Xt0^C1	�|���Y����P,���{�i���=G[���E�W�%����a9��w��{�G(ל(V�*FixجW�&n|��?�/��o �m���œ/��#3�(V����c�����閐YY���Ŗ�	��=<��Oq�#?ơS�H�:h:�p���Fc�-A���q�0İ�gAPM-���2z�-7_�?�����`��ǿ؄�����O���?{�O�ON�c��(���=���y�x��!lپ]t	.������o�W":8�@8�\��b.��x瞵�r��p�]R%�X]gG�p8Ps9��{�����h{��`yv��|Oj�8�B�Ie ����� ��e���X�C���vb�o�n̜�`n�8V�Qέ��*��VA/'F�ֹ���3��[�J�_�_X�t�Z����"k�����8TOq�`Cl\ ՠ�.�M���	��®��Ǿ�.���$�?�sE,����
�Ocl&)|O[q��L�չ$Q�ݸ|A� �7C���G常���7^;��Z��:�E��Цe.�<���N��=/�u�7m�!h����lɊyt ��r���ͪL�$�ʎ���tȗh712Џ��6���Y-"H�;���O�B���R*� �͗��O���E,3<���-��]�Mbl�YbG��+zC 6Deʭ2p���QTL��t���U�M����T(b =z�N��\(�Y� ̳��*
dCI��dX"Y�"Ѱ������`�.''A*��ٵ���:�I�\�k�JC>�?�����B��L̺Xʗ1���J��J���:�*�嬦E;��p遽�<<��x� ����Xw���u�N��x	�p:Eচ���Z��cs�8|r�J�Gp&|v���Vo��������V�ygQ�	��l*)�8J���6	���a�����.)~�;��.޷�#a_U�좀���~��[-#*��Eh��t�x�Ů�QAJ����~r�_ϗ	N�2!��s��_z-r^,9��QB���p+�܁�4�`��}B��:<�6�v�˄�N"ɻ"���^�G��};7���0���U)� �"z-6h��Y���N�rE�=�<�nD,J턗�ȏ��4%l �+>G�_<�Q?|9]�[Ǧ���iT]��QP���i��=[p`�6$��:��l�)8�߽�ї��� r5���*���M/j����"��N�o2[�eZ-�܍S۾�����=��Ov矟�N��Z6�;�������}��a���t��R��zd�KSkZH8�&�l�����Ss���E2���n�_��̓}�V�x���q��C�<*ȯ �F��L���H����2v�،������ ɘ_g���m�L�8���x����T�6� M�&�O�_�ki�S��.��Nr����s�D�Yv�x�7p���O=+�;_ ��'yks���B��ɪ-�~�-���Ʀ�a�Ir�CاဘB�R����4���?���4u�8U�����l��H�fU�=M09���1�L"��������W�����1JE>Ө�s!A��8<<�͛&P���0��������t �"�XS����|�<˸֦��0>>�I4�G�>ƿӧO#�Ja��͘��4��l�p��ƫ�-�R���P,�qť�`j�b��
N��uB�&d�|��q�7��J�$�E��B�NQ6�<�$��=ૅ6��K��p�u�A����|_�z��UN��x���iD��뿊���Z��{�C����1���J��l�� ��󿉑h��*��=��Z:����'�փ�G��F���j���ۇ` j�UPf�������g�;�li�d�ݷ~����߳����/V<��|��q��p�����xb�?��;��+.��� ����/��R��1I�4��{��?B��$���mINE���g��MW]�}۷	�I�Q�1��`Pq Mg/�����?�R;O�u����x�Q/��l"v��0�v\dnb���s�/�D2C��Z�x� �KY�8���N�i�RSh���:����_F��yM�X�QU��R��chu\� � %b˝�Z���m�p�8�da�'�XꆒQ��[�Ax�Il޾{Ͽ�ѭ��d+-d�U���c;!��9�f���lN�<ة�؍�M�+u�}�j����"� �cm5��_|E�d���`��wk�H�]0�4_f��Ȳ �����}� ���ykB�s�������2�}��(7*(7j*ԡiw�&o�x|�016��Sqժ!@�!�򳅔��/�`v~E8�>�PXxv<BA/��1)L��T��āh4.}z&[<@	=��	sL����W���5G�L�F�����$���}&�$�^���K�d��/R�h)�Ù'\+����4�2�r2�X�9S�C�/����&D�ZC�PB6W��jF�5	j��Ӕ/�sc���H�}�{D���Z3+,�_���B�YG�����.:{.=��?�>����C�F4z*W��4��;�^&n4�|�lI��KY>5��\�	�4�1�̊:�͚��x;�ߘ�ڂ�v�n��	�~�Zv�,l��ڶ<�=	�b�:y�V~��6t6쉀:���[r��&���^�K%t�daG�I�=��Bv�8��y�(X�G�!;��eK5�h����,F��$x&1�t_����e%Gv������!�򺙘�[Cx^��G����p��;6�&\ݦn96s�f96K-��c���4;L@{��K�`��F|!�Ԓ�@JB�Dne��B��M�a��$Ws5��[��sH+��'a�J9���7��K.��PϜ��]��K*ȑ��)+�� �`9��s����çe�F5��Ã��A	�� �^��ɒеȕ�ɯ�$���~h;Y��V�iI��	>�/6d���^���.�8D��>�߆o�
6����F��2�EzB:M1`��Q�!Qb���KDQY[ų���ǎ"�P�ʪ�	l�e�˟R�:ȦB����v�݆/|����k��/&�nrY(.B��&
nN;������D�@��>�a�N B��O	c����p��	W1vBF
Y�@$N��#�.�{����;��������.�E]K	ʚ2RƲ�k��h���]���O`d�DW�Eio�<.!��0��$������E���#J�q5���'m�&�)�y���+V>/�v��S����}=*'z��,2*�1oI$�06>�\��Ϩ�wt[h6*��Ţ�Kϗ�V+F��
���
�s��c�A�����̌�G7mڄ�۷[�3��ţ����QA�{ahpP1/�͊��N� �a���*h��&���	A�y�I<�G%���Q�u�l"�}f&f�c,��%�R��=��_�#��}�"�K���>�;�q��.ܾ�ԉؐk5���GB��-�_���#�o�;�<��_|�up#��������oo�{/؃�׉&���T����퇾gdŶGfVQo��'�׺T�#���G�pHk�0v� �U�m�}w�r�_��߿���~���+�z;��C���?��p�?�srvo�u���GP"NDB
����	|�;╓+��IHO�!�/W���Ӊ���ƫ���Јa[3������s:m4�)�F��i<��)�U�pc���pQ��x�-�sH������c0��@�8�A�&��k�V�rN��x�簶� 8D�A]gKw_̋ZfK�'Q\Y~�h�R.y���f����C�6����JΙҼ���$L �׭�q�JB�ny%C�;p�ڼ����۲K���J�fӘ���V��t?Y��c\��3�{r��^���$o��XZX��'P��st�Z�G�������I�� j�V�f�ϟ�P��c8:'7Ȏ�B��zl�$��q�5�ƻ.��R�@�x-�V��v�&'é�aL�Hn��4�5���9N��[���
��>���Q7r�~���	�$	2Y�^���	ǌ�!���5�ă�C)�,,.c���N[��M��زy�T��)��!Y�$�T=`�Rl28;@�`�Akj5�T:�r�&a����aL�� �:��H^���e'�����A8[b�i|���\��T&�͏�'N�¢���*UM����6#��DGdf��R��i�^\U��%���V�������dOa�� b~���R[Q'�J	]��s����ۥ���,����V׉\���tY�Ǆ.[�[��.C �,�������̬Cg,����K��V�hC8d�g%r\��S�z7�"!���1Q�ђ~t9�p�{���V2\�.S�>���2�ki�([+�Ɇ��J�-)[�GΨ1�\��B������wE	��`"���i��2dlө6ɨe<�5)��mQ� �q46��V1&�^��y$��#g����@{��a�Y����ER=U�����S5�t��d	y7�����r�:f��d�-�Xׁd�}	$�~��E	y�m��K��|Nĳ�j���)<>����*��$��+�#`A05֧��G�I��Є�G1�2�U�+=<��WWQM�2y��ĵ^d���nْf!�� �z� �ɾ�^�g����!��	���ɑb�b��^������x8L�YXҘ��j]ym�z��QK�Hs�Рr��t��"A�3kx�'?���|*EP&����_��̧"[�q�����O7��^D࣬ ��e�Ra�F	��l�0[�!䇞9��`&��flI�z��8�!ω��0�&�T��}OV�J��r������/�/��-��5��T�Qj�$\Wl5����������P\���o4���ę������P�e��S���Ԥ�"/s�1G�)�Mq&$f�1p,5 �$ľK�9����pziw��}�y��H�e��yo
F­�R��K�P��Tp���'e�rAf���I�[u!��UB|H 6S6�Q�����#��kl����YN��F�a�DaieU1���[N���L����)�<u\ӌ��1�#K����8:>�`$���XYˢPi�����p��-�~��nL|�!�=��/ܿ���_v �v���x���cf.�B���I�(W2��������o����u����������r�!��� ;7\��~�ո�}��^�������~�����n�Z��׏�"_j �������`*RɲQLwO}��^��T����]?���{��O���tջq����6:ddń0�M��7��_��}�t�#pGcp�����w�1�a��8���.�ܼ]��¢�F�G�=���n�����'�;����� 1r2d�_����V0>֏=gM!A-t�� �&yTJ�zp��	,LϚ]�������DP9#� �ת�S/bm�8��54����U��!U�TB�x�($.V=d�9`'�r_��5
f'�����\n�p��Í�b�O!���|�&�6n4��[w��w_���Jm O�F�!�>%�L	8�cd���m%~@i��8t'���`&aT�;r�tNZ�RBm��!�@wR����c���0��ˆ	�!?+eGd�(�(�[7��T���o��E�g_z!��)��פ=-R%�9�61�L`����c���c��`#ф8#o>�16�B���:���GG��irL�b�)���4���W�A
L���g�|�KKH�
r�dL��XT�"!8��y]�&��Hp��I����`�b�}���[X���'%e:9�	S�&ї��p�$~Fve簖��    IDATN�ް��nM��+˩X�4JV���'N
�ȃ����տ���C,2]m��\8������I9èy:�	pٹga�н�t��à�TW�z���ujϭ�V{�+f,��P�
1�i0�r8QhtdV6��aa%�b�aГ2��!Ɓ����"%^
�����n�U��� 8�x�硱��$UNd����mR3sg��_l��q���:P+R��"�[G����֖TP�4�� �% :SZŃ����T'��?$�?^wWe���3W��:��<$H�0��a��D���:�5�P'�·[\��\{�ᤫ�D�A�����^�P��lՐ�15ڇ�ݍ�c�����$a׍?J��"L�h�������������YzRT4��U)��E"�TA�}�(6Oc�?J�\8:�D���)ȇ�B��A��������C&_�\4��#}1\y�~��mɦ��MaF1N=�99=��χr��L��S�%�|�(N���A�Ѱ�,��$��Lf����n[�'�3*Y�����҄�eȾ�3^vqa�+a|uk�d�3S�s3��޵aEvajs(騉c���)kY~5���0M9�~�HI�F�f��\�
^~�i�>x�n[>�;�5���Mڷ�L�wu�m���o�l�u�\������Z�&,9;��;6Z��<q�L�L�C�5�N����C�H�g��s��H���Hؤ�V#�1جw���M���c�q�������Ln_N�W>@�����X@6�ZV���7	2491�zW���D�%�/�y�˰�n��H��b�qL���	�Y)����R���+��� ���{�h�,g
����qǝ�bzvE(	[�����-yѐ�luv�{-q�&ƇQ';������`2o��L��sB��~�TY�Ĳ��ӧgԼbG��!+�]��H������U����W^yy}�&���V�T1#O �!��ˏ����L�2'܋9��\Z-L�����p��{p٥099�`Љ�t/��&^|�~��A,.��X��6�%8�e|��_�_��籜i��'��#/qBЃX��:VgN P���\�����8o�4�@6���ދ�|�[��r���Gg�&�rDrj]���T�3�VuHƹ�Y-��:��_�������4���_lB�L�������|�>��_v�>��� ���=��)��?|/��&���yѮ�Ь�0����_�����"�'|��N.�������4��ޣgA�YÓ/�ZэH��Tb�6ҹ��y��$!���+�aח�YbT�}�ſ�ӗ1?=O��dЯ侜YA���`2����ԅ�O��I�Yʓy���m�C��׋-[�h"@M��`2�]� R��-�T"�!�\��IXl�e6e��M d��BȪ�hE	ǆF��[0�u&��w,��BQ�L �<���C�b+�5�R8��@� QrO�IV�ȡc�k�x#��(-�D��L��a.Vv����V�eT,25�"U�����r��d����X�;�J��o�.��l��.����y��{���j�U�`jr��٩�4�j�]0��Ǐ�B�م��Sp�{��FU���Q,��c�!!دB�Tj��#1��i'M�� g�wi�477���j��rrdE��PJ�+�.�+h2���r��U௔� ��Ѝ��E�r����!L�����֌y4v�]X��Ҋ����pTk�I�@��"%�J�2V��p��G�z���`C#I��T�6=�DU��^�St�[E��A���E���������A������L5:dwGD>vlVBv�F��q��]Ҁ�&���i9,���8$y��SR�i�XL�U��E�v�u�[��3��R��zւ�
U78�z������#l�1�z�N��Q�&��yx��>Ƅ�P�B�(O	��[/O�����fv�+USk� �0ԁȢ��"V�2�i$�BW]�7�0	��j(�}� ���!��c��c{�F%��[?�a��@,�m�a�&��M����n�bQ��VA"Bdf6���5���<�4ڏ-�Cr-�!�g"Ԃ�����vWI�׸\%�(���xGO���4]�ˈD�	�Ѭ5$�@���[6	81����U9���I(%�]���XhJ0=�مU�,�B>�n��vMat8�(9L�(�H�{��"øD�P�6Pn'�s8��šC'�Q��� �_q^�/!����NXR&6� wҮT�ΞxY��S/GWE�q:>�b�n��;�51�gT�X4
��uH�Q��J2M���ф��)[V�� �PY�.��O]ɱ[&|ƣ��lN6�ig�ˉP�ɜ��O?��o��^��F�Q$�۪Sp@u�9�04��b���}|�un$�)�p�X���0vi�����9���%e)�pX�"����.�,OM�|4�
c|xHg+aH�v.S��	_G����b'O����
�
�tz���E�L��f#�͙6�.Ɵar�(�}�e��s�&	7��$4��dV��i�̵L�)7\/N�wZýJ[8�1��?2~F<��;$��aH/�GI/�h\~�hp9p��|�λ��%j�x�p3VX���3'��*��H���c2�� �K#���^��I��8�|}�3�+P*Y�$[+d(�R9dÌ��?�gP3Sw�c>g���pD���"��ge2�'�T;M�q�d�*b56�V،u ��JX�L�6�yghrid��څ�������aDj(���{����w,��P�wQ�2U~g7�W���y���}O>��^{'�id��\^tȟ[]�z����>v�� �Nd�{��R:x������J�FK��=N�|~x}!�!�k�wM�;T3K�s����}ꆿ���H�������o��/:�O���&v��H�����Rx���ջ��g_~=o������p5�v���ބ��=���_N���(c�}9^o����q �p���^z{�J�"��ڬ�֪��k��� cx$��d�	.��%�"���2����'�x괔�:�,�H9e(������N�:��Z
n�kF��z��I�R�:Kč��t4��*T����ꓚ�z�׼.:ҩ�V�ݪ(����\�ǰv�γ4&i7{�V�����o��QL�}�cSh�|"i�[�!þ֖̪�rґ��-3�w�[���7�M��t��:6�J���ë� 7{�|�Lhr@_�2j� S�`��1�m���L�k0�H���8�a����п}3��е�z�^���pX���f:��Y[�ԡ�~r_�Қ�����3;��F¡Qr�m�l� ���~���h�@�C!].k�Lc�"�A8�� �j���N��j �Z�u<_k��ID�w��y5	��J/���ԍx(1���$�y1�i�H�@��v�mp��Z.�X�x�A~Ƕ�j�sH�s�f�p��ך8
L��x�E��\W� B������B���a�Ƥ�Āۤf�/���<fWH�Π�ȣ�_�x?�s����V���Sc��$D,�8P麂He*x��I�8���l��8p��ضiD�0&����^�VSң��q��<r9�.ٸw�F��`�i����Q�zgA`:���>5���-2�!c�DɆ�,�*	�<��A/7d#WHI;xz]Bk5�\����0�i@��]���\���gL��1C8U�$��4��xKՊ���<+S��Ũ�{���y}9�#Q��(���PT�Hb�0�69x�m�!�=��ZJM*�7p�c�"C��j7���;X���h
��+��x�:=��������\>�^ZƉ�e�Y��J^�@\1�\vc��崽ur�� ��)�S������*c-�1���ť4*5I`����sv�=[�~�l^�:��,�Y'�sR��n�NŦo�Ǔϼ���B�axLb���B�K�'��2�({�<��O���!�����DɾR��Z�lb�u��!�T�� �"	�R@��Ʒ�6֡���Ǳ
�@.�@�&�>�	�^NBioEWtv��J�8!h7JH�<�Є韟����|V ڄ�PA�r�T�!_�q�"�iٖ�P��&Z��<�������$�%����Ntju� �5�-�F�һ�̿�b\�CA��5���J��k��<ë�|��#�i�C����Q�	J S�lP��(���_O�G�S�Uh�����D.�yD(*8��K����|��{����d�d\�]{Z�#6\�z���|LuyV8��Y��g�Uʈ�?|�0N�,"F���j�h�"�ÿ�6%P���pt��\�|�w�`מ\�7�/���4�YE'�,�lNxx�

6u�ߚgmO���@_��)�mPy�t�/�H,�uO�(��4+�E�g����������h˫��f�BQƢ�� >x�5��Gn��][��p{<��!����+(V��7q��C[6��7܈^Џ�U�ʤ����Ϯ>�K�;�Rgm݌�}�j\�k/N�:����<�9pz��khtz�R�>��E��]�d�b���-�P8{��?����������/MA�������������n�W��������G��˯�C�=��<���$���-/��CH�:�59�߻�V����XY&63,<58g�R���A��E�L�Zxk:���*ܡ�T h@VmT�����8�H`|b��R���.��?��'�dfmq����o�IY'�C�#p�,�8w44)�XɐcI�$����I��L�HX���^7;��b)�h8~ukY�͎%-mp��VS�h��cϘ<��׭�����&���'�r�Z�M8���/�Y�_�Zϧ�n�C,85�=�r�2��خ���h�����t_ؽ���pa��<
�<����(/�@��6ŀ�����Ј�$cg&g
#�0j�[���]����l��4�{|�L�٩���j"�HhĘM��7�`bx�F�=��%�J��r�D�
f�5�&��]ܠј�qDc!��9�g�Ǣ�^oK�he9����7v_�NEGN)���j����o���P�'ל��ouսx���h��b� $��atxcc#�Y#mv\�0�!q��YKM(1�)K3�Ti`zf�LQ�>A�=N�LA`�x��Q�����A�W0)�K�İk�݆�=\�,�aa����j�4B^��,\�/&�C@��%���O��f�P'O���^�r��l���ؽe
��wF��.������r��8���8rt�3�|t\n�E���{��di���b=ѷ�+��A���3X;��cc�y9M,�>8	��B�����k3��VJȮ�Q��Q.�(�.��*�RR�A��B�� ��C�ZG6���Ґ��2�ǎa.W��gA�1 ��>\�0|����(��	��h����u\5_�ŨMb�I�6�JŎ�d�sf����̖��'/AMv�Y�6j(���훰oפ
��g�&(��KU"k*�����l��(��XX+���"N�,˃��R	�׆�K��h��6�ɑ>��m��qjK�|���.3Ki�
M�d���O!�/!"$����={���+�G�׆��iu��-�'��׭���6�D�Bx��i<���XZ-"ѷ	�@��1v�t���h�E�Dx�(�*e�(�Qc�/Y�X�"��4'�$^�C��b�!���۱ԙ�l�W2֞0Dz�����Қ�D�]��'�<$��}�iZ�8��N���p G�?�N��:����
^G�P��U0�l1N������������5�?\n5H3)�Y��d�m�Yn!*t9�ܨ���F�G��m��~�S�X�~f"�6	�\�[RDb�E$!�)6M�����l��E�YM�`�c�bm�&�v�v�����0Me<#�)��lT�e	R�S~aA��Ӯ��W3 #��n�.�u�$::t^(�y���4��
��4�:$��q�ё��56�b�0\>69��O�|9�I����Ԭ&���S��5i��W3S��iҙi%L�9a7^|��'\8�agf!���x���@����9!qE��R��8��d�'�)�j%L��⒋`��ޅ��>��_'O��G�?��՜x�$-�Li�j��H4��@?\�It"!)�l˷�SF
)��4
9����;%�==?g��.7��
�
�2k�+/�ӿ;�:�H��^�D���jf!ζѯ�����_����Ǟ�����Ϳ�;�W_v�徫�{%�nǫ/��~�
^x�f�3�b&����8��W_��wmC���+�}�(��66o�"3&��2��ܖ��r��bׇTՋC'���U�PΓ��b9���*)nD�b�C�������wF�CO �Z�F�T
���2���{����6h�2(�R(�����N��t�h_X�p�Lz��Z�j�x^�/��Y$ͱ~Ќ���k)�r!��H�)�yq3���kb�S�-�	_*��G�\�I� ��v`�������\�5v�}�_�����j�4�����8j/��AX��+Ȯf��Z��<EB�(��r�%�[CD�@���,�)n�L��?7!�
/;i�&�<���]�n�$�,�9!�Y	ݤ�68���@	v1(�֪�UA�=,�d�x�a'�HĂ��!"�$:<:]��e��%��lA�";f��:\���ԫe�4	�bj�8�<����X��g���0��f>�2��4t���>�k�#4J<$�0�m-s���{Ȯ;�|	��(W
�.�'��	#�i�ۂ�3�3X|����v411�ĶM��y����jˉ��˘]Jcyu�V{wnŕ��-cIx�jW�#'�K#nJW���B8t�4�� J�ʀM7�Zu�&���}rL{��&���W�K*���t�|��#H�*pQ���n�!ȓ(�1q:#�h�Nl��ܚ��Rܱd?�} ���v6�{�"0�L�,�0X�`�&��"2˫H--�Ʊ�mt%D��6�y}��'F�'^��T�i�K� �R��Z'��k&�*��7"���Abx�xL�a,�@83dw�n�\!�R����Wb~&���g�l�Iv����'��,�	�T�j�QΧ��l���{�aj,7����Q��nBi�E�K��Pd�����E>v
K�Yt�4SJm�	�Xp��:���>Mp��
���	�<�˂�Eh��F�XÉ�,.�
B�W.�1<ŵW]&ߌa��|l��!7�C��6���͞GO.�g_�j��x�$-�t��脝o���M�XU�G�3��MI� kơؘ�� ���5�Ƃ�E}�>!�bP�M��F0B0#)Y���M5�#��m���c��[L���p�p�:��zx�D
Ut�g]�k�H2�P����~3�D�\Q�(���2��zfB`e�s[��ru��U&��
M����7n��C��H0��QecM�4���4)ƅB����w&�$��9���xI�\�g�&72S3��	��$N4Fq! �<���s�󔿊ϧ�.��œ=�/�F�o�i'���r��4΢[��-���T���6�=G:����9ْbԵ�}��̻<.xk�D^�i-@S@^�8{����}��BQ6Ձ���^�s���Y�^_ιs���%�$$H2�L*��s�����Vmm��Z�\��1�	#�H"�(����FI�C�t�_9ǭ�z�wf|��?�*��L���y�羯�
U�*ZkTAb��4L��k ��꺷&SdM�X[[�ԑ�ݤ�͋h]^�>�믿�R���c�qEg�P����oWt�V]�_lڸ{U+NW��[4�V��?��]ݸ[z.N�i���^F��9L�oqy�jU2e�	g�ZMt$���"<<�2)��~��#��)X����&�����=���b�TjuTic&��O@�>��P�����'�j�:u�2K�}SC}�����~�(C�������/_Ng�w:t �D�{����x
5�p���͠Y��S�P"��o�����"E��j��t��t#C�8������>�    IDAT����]<�����^lT�ߝ�ᵳ�h:�Fc�W��oJ��#K8y=Z�~�;б��1�]����zn��4�;w��E8�e�rk���Ѩl�^�K�ʃ����lv�SP�U��b�X��9�y�R�1�����l��i��Η�Xp^�pďd"��(&��~�;�M�կ��?��ǸtnF�`�MD�r�����Y��+܃���p���@09�����hs|�����M�%^n�1�����ʗW��tc-���]i�Ө��9/�IZ�Y�7D���KCS0���� 3�	۔!�ؔ!~�o;�7~�^�G�����a=5G��Jtujjؘ�%����
.�.!���Gd��wW��=� $@ۿ(z������g��U@ԽRmaiuS>��Ey9ei	�b�j�L�E<B*��0�M��L�Pgspya��G�l7��Q ���'��}�.(Њ�w:vԉ�x%ТO�ym~U����Ng�j;��0�AE�5 �Tt �~���*�H���R$�]� �q�M������VWcS6Dk� n<���N�'L�W�f��m�AuQx#q�gN��A�Յ?A�� �bA?�ڎ��>�3��H}���*�jM'~���pn�kt��8����+{C(�Ud�6�#��C�ᙃ�jCp���>��^�.^GN��!lm�Dg����u[aq3�Z��F��R.�J��=�3�A��}�᥆���;��u��h�K�%�d�&xݸ�(8�B>�E��ޯaп2=�r��xɁ>5,���;���U|*�Xz�ȩ��j�M�����+����S��e�j9����i�d=;:ǡ=۰k�a?�jV�%�Kt�4�e�H���MN�����u����YB�z��П�u(�}+���_ "'�\����Bg/��r� 
�����b�����cj}� ��6�L|f#���$�I�h�L]�7�ұSXZe RJ@��*�,:S���'�UJ�����j�:R`�����֘����Ÿ�v��.�nil�6�=���@��t��]mTXs��cY#[{�fO��0:eQȅ���M
�\\��B�8Q*P*��su0ڗ��QǱ���ʹ��Q{e�Bl�Rd�ز৻���,Xy�-Tj�H�a��}�M��wtQ��s���>�;�׶��}H�_k���dcP�z��Ϣ����<Õ��!�K�_O*�5�t
�9ɣ��5��p�V�$Æ��3�㤛�5r�Rq٢H�b������f�|���"[�!k�a�gM�]�^���Hi��~Z3�.�E��;�?Y�iF��E$	�o1��L*,p*�	T���*�.�8�ڳk'R=	�8�&2�M+;���Ȅg�9��e4���[��rEZ ���צaW̱�a����ѣ8z�z�^xAzi�D34�:
~1���X�ҝ(%a.�{B��W[{�hVdܑ�E��m�N�D5�R�H�K�q����Ґ��n@�"A�?�TBÃ��Ƚ�f��*��i8^Ts�(.���0�;���z�4,�(0̜��ܥ��Ia��s��QC����75���?��߯�����0�_���W�,o�I� �J!_�I�é[8�'�R���q�iIX/�!������߉�}a,/����<�S��ƽ��G�\we���P(V�!��:��=.\^~{bW����$�ڸ:�B�5��kr���[H$��S@F�z6���"6�f�]^��]C�ZP3Pή�QɢU͛�1�N�cn\n4�3�>L)�P�J�;�.РC���Ƀ�� iBSSS��������/�V-�С}�G.��fzG���C���,..ṧ��3O?�'ϠP�H�9?������&��1�>|�ߌR݅�l	]
�N�%��!�)*o��(4�NW��:Dr;�e�H��Q͗��a�[A���� �#z��7W���7����lVr�Prn�S�GW�����~?���tyV�.�&z��U��ѡt�Et9��F�I Xq��63e��Efؘ�X^��"j`;�
�Q�{������D��RNo.E�D��d�fMv�"G��@o����)�4�@�99�ha-�G����5~�mZP����+�Elȹv��!��ȾV��nDJ��q�f�*��(�=�����U�e�Ce��lF�-�ɥ�7D<�4�6�J����u�q�
Ͻ;�px�L�� ���(t}Jĩ���.r�Ƭ��9�I2#�އ���qL�bd��	�ܘ����/#�;����8{aǏ��Z��\�8����1A[�.���e�fTg���u%�kü�	�*Ux�Y�领vš �
��Nt�R�aaf����U�E4+����v2���Q���A���O-���٧ج�U��@�0�Fԝv�>�D��O�S�6�̃3��"[��q(8��:����#��n�ݠ��!��Z���j�X[���������T�EKaC���8�`���l��W!W~W^r�8�>�j^�sǩ	P�̮lH��)�銍�]`�ȡ 5����q<4i񵊬���]J��5�źl�)P�T��)#�[EOO7�x {wmE��D��@��}����%a�֤�_��mV3%�8y��Q��	�����yV�&��J��I�'���\�`7!�xXz+̬Z��C��x���8�b�g;m�g-��@C����`�����;ż�k�Y6f*��³	`6���,��i���ZF������P*�N!�W�y
���<^�j5�����q-��$8��Qa�@p�*S
C��ǣ��R�
xS¶��f����	���bE�/ݟ-s/K��#��K�G�"R�9! ~#�o�iB�:�"��nD�,�Z��:��@��Ԩj���Z�_g�ҍ	k4��3�m�a�`�4�E� �R��&h��t[��������v��k������kh�v3@�� ��i|�|<5V,�%8�|��m��vuj�M���NA/��.���A�>�m�&q��	\�|����μIƓz�l
�6ۺ�y�רյg����v�v"ƿ#����Oׁ>���א�~�\Ƥq�LR���4Dv�18�E�@&_�C�m���|�c�G����d"�:m1�\s�֕M<S_��AFϕz��@?�##p�"����t�IʲO�ג���QC#�C�XhAJ����N� >��.��g�3�E)ߤV�%���?=��O����������/�����.�o��/��%�zŹ�w���rЖψ���"z�^Loŭ������9|�_Av#��~�<��l�Ws?0h3ܪ.֫m�rz��Y@�F05 8$n|M�|F�U��;6򭅶���PM��ӈ8����S'�p�Z��!��Q�o�VJ+���,�>�����-�21���6�*�Խ׵����P�,��A5���H�l`����am�.������s��?E>����_'����	�Umc��"����'���o��d��oL��/�4<�Y]G�e����{=6�U��w���I�eC�'�D��V.c��0A1_���6�@�wq����A�! ����9�M����8	���әD"l��`tvC@Q���n'&������a���ЊPms�*?l
�Iu�(/��\ʙQ���;�W_=#��X|@(+�uD�>�lڍ�>[:)�\����eC7htJ�	y`����%�����N�)Gν�$�R�krQ)f���ΐ&ڋ�AY�T$�嘵V+#�M�T������^9a�q���BX��IP����$���A����"r����?r���U85:�����,�I��VA�Ot�n����%F*B"��hE�\���e�y��F�7�߅��荻�B[�Ѣ����D�]�'Ϯ���0��A�EA&��{��̍�#�J1�n��m�.������CB����\�[B���Ój��\�,�b��}@�IsS	����BJm$�
s���]���v�%�6���Ni5�K3R����B.�x�6WV�~٪�6,=}���>�-�S��g3�RD�qC��f��¦	��2�BemZ�b=���4�<T5]�b����sB�\?z��k:$�I��kj��Ĥ�a����S+A�v��t@E&-��� ��kD����t���r�ڳ}�����ߢ���4�]�?�7dф�>�BE���P��ߥ�b���mB�B~�l��8���c��0M�b�r������,�\E��k�&����M7�C��E��@�`�ǱD�b�H`(Wץ)u���KK8{q�kET[N9���DMe�Ll~���D�8�
K=��M	�%����uަ1���7D٬/�V�17V�! [xC+7�׸�slD屨:L���M��<L3��U��df�h)���4�c,v��{P�X��g�Am}1�_A�\��f���� -��@Bb+<��N��"�7���vC���ǩ�����+-�.r�	���ִ�ʴb�ĽOV������UI�q3A���U����{�Ӵ��O%E�U*9��8���Z�� �� \�y�����Qj�E��笽Hoa�P#��Zt�i�!���f�
/tW��f�d>'M���
��c��1�����0��Ts��~�P��j���B�D�Z��e�ģ�퍊�Ө�D��f����vE����.xf�2ן� �1��`)���P����#���@�
�S�h`fjFǾ�����¼��I�N��F�HCC[�-VQ(���4T�{����YS'f���n��[�A����>�}�4�&x�k՗J!::�V�TV:M�5! H���Y]:PU+�M ̄�6P,�~�@@S���}�p{ec����I�n��[��1�?���?���vg�l
��?��,9�E��zv�_}���]X+�#�;l<��� 6�=��%`:;�1(�eCbڤǉ��w����'�ۿS���>�}�����)�5-vk\M�F���@�z�4^���p�©!r�My󹹹�f�R�/���,70�׃j.�מ{
3'� �E$H�Y]@�\@���L|�Jd�q�zq�-o�G��6�߼�N�8��"�D��=�����-�܂�{�kDix���	�<��ڒJQ�l�7��J9�����?$י���=�wv��`{v��Ėm��x��q|�[��w��O@ǋdr ng͎]g�B��	���w#��ٹe��Ia�+	Q�0�7���A��Z��8�r���kX_�@n5g�d��,PT�qd��e����!�e�)�ݲU���!`iǆ�7c�G�����0�&�0���b�*�6d6n�*z"A�F��0�+e�����d}{�Č<����.��Rq:F�0ЗB������dJ���*
Ŋ���,+Y&�k�Ǣ
t3aHSQ��6��X4��T�X}=18X�UK�0��{�
Z�,�5������6Q
����"a+t���C���z��Q�Ě�Xo��c3���Z�F�T��^��zUkqaK��6�LzS�ni���=;�0:�+�7G&0�g2������e9tvn�`*�¯Uˣ^������>ml/�����o�-�d[�t�F��-�!ҵ�t	ý1���[�/�t����Zi������bu#��t�fqiam�v&�qB1�!��n��Z��Km�
��?��dA���TtV!�f��Q�Z���s2 ��h��:B<�s9��ϡ����hd�lߵ�8��F�J "[, W�&��av�
�T�ψ��D�
Qb�.-���y���u�����-//ayn�h��!	ȩ%�IA�$��6��~�Oi��s�T����K �����\��(R�?��VJ� U�j�}1�?�]��q|R/"@2b�,�~��'��iG�D�dY�p��� _�)Ř�:��F�,/v��!XD���l��5$3��`��X�PQa��pҴ�^B�XE�Q�����@�{��O��8c��m&'-:���)��
Q�403��S��q~n���p���uU�Fp���돨���
��P|N�,�H��
]יG�h���ۥ�iN<׬u6��7�,a�VC����ոџ�%}�M#g�}�8��/Z��և5�j���	q�x�� ŏ�N��9���g�XO#D\�a
Z7S٣�vdp��i����cf�<{�v��Z;l��r�sO�>����S�Cֺ�F�ƞ2Jי���:��˽��=3��u%A�t~�ea��W�K��ψ��'ɞ>x!��Z�
m��c�xf��DA.�e}V�� �J&�s���55�HM�)��V�܋�1Eo��ub�}5�l����g�z�Y{?o�c�N��׎|y�{|}�t8�B��$��a����o�4�7�q��qM�wLOJ&�I���?#c�z�nY.�� P�DE)�s1�����ҙ��5@��iӖv��	h�f{�b5|����@�iP�� b��~~s3#m�����~���ȕj��r�6;:e�aٝ]��o��o��6�Qo�F�~��ؚ0�af�G7A�ق�f�^�>�H4��)�V*q�無�i�{�Q���Q���WE���'j�p�h�!8�{�o?�����nٗ����ҿYC���<?�_��Wg7�$�e�M���9��<�ޕ��@��>^�j�V,���0=���X[����;��c#��*���_V�7�HK����;7Wd_�H���nur�حʞ�+w/9�.���2�!/j�4N��6f/"�i��h"����ʂ
?(l�c.�J�زu����y��������`}3�W����`pp�M��G��F��.,b��� �Ã�MB5�ř�x��_�_�LBݽ�v�mo}��x:�K5�|1�ص['���Ep��,��7_�?<�u������!lsFp���1�� �%���0�3^Ӥ&���!���sM�#�U���p��������@�hS��xR��1�P�k����X]��n%G�߭�@�Y2�ĵmb`�6����`xzs��(��"���c��02k���&b@K�vۅՍ�&�f�^B0�F��!�(>��;ɛxyuU	��rM�4�J.z���Co�nC=Z��M�8�mq�����0Z��P(��:i�ϘNy⺮Ԫ*��YP�AR��A
	7W"�����ur�̃�p�$��T��R�S[B6�r#�������D�V�'O ��F4����3	a�����B�(n�0���gN#O���sl ��6Z5�n�
�İ��ca��_>��T;nxBa�*�;�v��b1Ԯ�Ь������c��-�5��m��2m3���fh�z~v��VQf���-j�,xixe�u
�.�7_��UHQ�%��Q{Re�ė&���Ht7��|D�q8t]s�^�*�*Q�Lce~^闉�al۹��Q�A��植��B[IS��5boŕ�$E��t�S�Yi'm"�U<h�����M�H\��&f3��l������G��m�B؇�A��<r$��f�,��TO�69��d�hc͘��C���k���q�Q5��}�0n8�G� K=�+p�j�+���n�(w�� ũ�edK��x���gS�Ϙ{h��G�T���Դ�v���J5���v�	�`e=�7N�`m�4�Vng^_7�x�I����)��g���}���[@�����5�~j��8}&̨ط���!�l7:J�DjG4�3��+o�F�9h��0�l�,Ꜩ-����u̐G>�lJ͔��i��c9qI�f5�f�ZX3Q�T�1x���x��O�٪ʚ���}c�_�*˫��15Dn�h�lp���v���FD�!��Ǝ�lo7�{wO��'�B�͔]Y�Z��Vn��᜛b�ȯ�~:0�5�s��T�gis����ip�7�Cم6���ܛg�p��E,��kB��x�6���E�-#j���&����&zRq��J�:2:�ϖf!n�[I����5,�����@{P66�^�`�%���^ �i����<`m���bE�
[S6K�p��p��S�y��{���=�܁������a��عc�&q��./.��s    IDAT*_)i������&��>�C�`t|܇lʐ��]3!�����B�eu�i�E���j�l+R��8��{���V�x�mL_�O������!P�~��pS�o&��KN`�,��V��5�f{�,�9�� N��a�Z	bp�a��˥�. 5'պ�Yj6����:���2)J�R2!��7��K��Ԕ0���F9��yp���~�����O<���i���^���׾�������q�ӛB�xS�M��{��`^�oUt�&ǔ�{��yq㾰���v�Mx��a�֭��R�N��[��!����;�҉E�>��P�4�^�TJ;@�8���S�p�T7��nM	ѝ]^����+��3��Kh��(�� �^E�l
�V�HWYB��{��]w݁����Tr����������LLLj�)�M  �3.h!�^��)v�V�@{�D���i|��c/J�C��[n�A��ܴHF����a���Xo�q_�[x�;?D��F49�HlՎ�����;�6n���C�'-��F�����Qt����F$��{��,\�E'����F��)tG�U��]��)�Z����y4)�kg��{��v�!����<J�n눂Æ���ɱ!Ye2,�bF�Q�<�kD\�B�%���M�x��QP�`o
I&n*q��l!+�[&����U��3�6�p'��BE�c���:�ZV�@�I�hժ*��m�5��
C6f�i��Dr�h��hamm�/����bێI��2��4<9.71��A�n��5��AJċ��@'f. W�	�VfC$���>�(ڪ��5��k]�\ǩ�g�}��}8z�D�Hۮ����@.,�w<XM����y�yv�R�`\���DM���LK;Y��K��3����w���i��>	���h#�/ W�b%]��f	���L��RG@Έ��v�JW �뫙��5�j{�7��H�M��_��W� &ǁ�fIt�-xju46��-,aci�f�&�섏:�`Rt
ч�S�0@�!kjF����p�%#$�x�^�^K��k��I�Ԥ<��z	esK�QD��ss�e�2�����|�
��5������Ƴ�5֪OacJa�N�j��3�bSXq"�'�%&�zj�vnCiY�!� 0?���ƶ�|&�4�_�Æ�VG�|���q�yJ[�v6BјV�)�U��:�w�No���\���V�NӞ��,�\ؿ��	�%�
;Em%�R�H�G�*��Z��F������x��e��f�w�%qa����p7��2	 �b���P�Q�If�H���~��p"���ڲ��Z�����,��1���7)0A�gZ�J�`>ZF�k�n�8[h�:ZKR���l&��Bg�[�i�uw�(�.��/���7�ݑ��%�N���� ��\��j[A�۷M����m�"�I�Άў�j��^-��}���h��aq�&����G��j���-��%w%���w=����~�}���܋/ɨ!OJ3�sT����k��W�D�!��3���a�i�9��f��2�Ӧ��qP�����yf�
C~<�R�3K"]��g�TT�Ub>�����I��Ҕ��NKK+8u�����p�i�Apå��S�#��G>���!����!��@*��� �(r�fff��e�<|/��)���>�Mg͉'U��K �E�����l*$W�?Z�R�`�r��х��4�S���	Q�����p�����v;^x�U|�?Ź�9t�L�%_�dvH�+����&
��A���n��&��V��R���q�q���F�6���k=%m��&�ȻR��%k@�oK`���ʪ2�t�Оפ}s�s_Pc��"�rys���~�����+��_=�Ķ/<���E���v��[\������*������	yä�4k5����[�
����ҥE�]>5#�	�t� �q�͘�܂Q|�tnn�u�kz���x����Ө��g+G���P,B�D(~�Iђ�	E���rǞ�g���T[z(�Wp��c�XY�&խ�vn�[�q�߃O}�c���� o��t9��Dbp	�X4���H����4<�)�Z\\�ɤ144��;�%X���}gϞ����=8r�\n�&�1l�gUhLLLa��n���ěg�<���<�:�:�V7+�Dzq�{>�m����F	�ٲ����,��5���aO≔�T.�>���%t��(�a�*C�,��6�Y�57Z^�!�i�p��\�jq�C@��E'�C#���?��lф�\��F���&kT06؋=�[%Xq&�n	� �~=���@�N�@s�������!�Mđ��_Z����e�y�
�-W�H��&g��
N	 v����dum�k�j����ăe��F�./�Yt�8�Ř�BX0RLZ
�b�3U�H�-4inqK�+HD��1�D2�һ�F��Qn�^&Rp��Q��HՕk�=�R��
��D�@�c�z=Ȧ7���,�RG����,��89��ޠ����^�}�Tj]\Z���i�)�?�8�D�s�W9�ff�n]Q���4{�ػ}��BO<,�D´b�Ց˗Plg��87�����C �1��wo�iEK!�lβ��AdL
$
����D��� ��!���ɩE�R�\��u��y��qD�/���!�e�NU��P�~'�N}F�~�4 �>Q��U��;���&�}ΙK��V�yO1�����xuXszIԱY�"�al��z��s�
e$�]�SL���0_�E���hL'����V׈�y����z�]%u�fr�i]ؗL��091
?�:�ذv5ᠠQE"�Q0|j��l7�i�"V`���J�p�v�р���S�Fڊ,<i��\kc#W��r�έcy%��n�K��&'�u4�m�H����	x �����#�Q.glj=^\\������jN&�ӊ�a��Ԙ�Db�I:u\�D�=�i�R-�3$ji�?�
�^����r�+U�Lс[�o>]SX*A�U�vڴ3�56�5�vT�˚Z��=!��d�)Qظ�:j�������7�nр��9���/�x��"u�!#Q�Ȑb1C�*��1��լi���[o�g>�1\d�\�:n^��x�rЙ�5�-$5(�)0���eѬ��**���۲E�"��{��WWã��$6��[`a�������wq��Y��a��������msj��9	fݧ?�q��waj[���%m�ױ�&����^��ѴFv��!���.�H69��=�)&�yZ`����f�Xǽ��CXYY�SO�
?���87��?��'��BF��7=�O~�\�a����ӿ���g����䍔���u�+:8���Ԁ���Ȩ��k��f�_�f�I�_�Sԛ�����럛�\�\i"h��a��m��;w�_����al�v��ǿ�7��]�8=���x�u�1nY�<1�B�<Bw�?k��ɱ�O��k��B�E�J8d5A�4���v�&��׎g?�èTѥ-��	r�$i6�ҟRW�=՘Y$U惡J3�s��6�޻m������|�37����!��?=�7_��&�y��>���Z?���̙3R�c	4:]	&4��0>>����h�z�1�9y�uu�ƃ8|p�~����Y���Rn'���|�"�z�4'������P��r�D|[�=���0h�\E�퇣V������&����PZ_����a��)�|N�v�@�'���t�����u;Jłľ�Xuh��\T)r	+�.���'���о������+#�B�����f��d��ʱ���^��؈��;�ՙ�#W<�c�
p��%,�n`xh���~����x����X\�`3߀˗�F����8t{��8�
U�J%�n�3G��m,��t�xc���6��r:�z&���"����\2Hj[Aj��S})�ǲi�p]�[?b��pV�`2��X��#A����O��k��F9��߃����2�Mnm������7�g�%�b����^Ƶ��H%��I�~��+G�&<��$��I�h������$��g	ʛM�o��g�E���1�
���J���Z��͸Y����fDhĞ֡V�����%5��q��|J�dc!����&s-�  �Uɝrn2����76����l��$jN��z{1<�/�5���U��ƌE�����.��ݎ��~����U�=�YW����'����*^;uAH~�w��d�,bR�8)`�%�r�Q�|nD��">$��łHF��E�ㆩ4�r-��gW��+o`v~�hbѤ	��d�4+L늓������(�7n���9(`4S���>�q�wk�M3Y�����js���D�^E�VF� i�N�a����=�9��O���x��8��#��鹵^H��ƁM���	x��Ѵ�:�E���)�犈����ST+�ʠ�f]v�L�`qށ��O6}�xq
U��ӂ�O��O�a��nK댯��C.��ɟ;|� vl��h��Td�ָf8�,�dY邋���L�)[RWD1d����C� Î�eQM �gf�`�}&-����ׄ��aK+y,/�0���isk8La|4�];Fџp#�n�k3����G���S\��a9]���q��2*-'�
��o���V,?w
�IC�$�'��\.-�8�,�y?T�u4��Ɩ��;g8}}=��������a�{����-PG��W��u��X���g�gR�Lcl7��L�ŏ��Y�["O6�j8]��2ԇ��<~���7x6^�RN���i��,ǵvCNc�r��_ӁO}�#�O��J�!,Y<���I���Q@�y�6?�v^34R���@T7c�ˉݨ����CQ]���]�Xɔ��E���O>���m���px��F8�w�0D)�z5�T��Z5�ٟ}���'0<���6ܤ���TrD��T���hjI������h��W�f5�W��)�7�>��18�Q�Xp���4�x���Շ���^<(�ƹѨ"_؄��҄����(����P����Ə~����+Zσ���I��+6�g(.fC�ό�'O�縦m�֝eMl�O����u�t�c�5���!H&E����O�Ї�����?�(N�����2!�Z�k�ə�S�purl�>$��F�^u�\&>5�8�Cj���0g�j/�.���1��c�t���T��`l����H[�=Lj2� '����;���O>v��&_���ۿ��oyh����g�p����Gy+k�${����������u�͢�|�����3sJ�3A������s�{b(fr:��Q5����	��p�翹�_��M�mك@j@´]oܠ9��[�����<�0�)S�����y��D0rc��i,]8����X]���#�д���wݎ?��}�E�Y��	��0���:�x�˝���+���/|�o���g�	�yX�g���|�@��C��ff]��SS��>=�(o�V4�&U�Q�%[33����Ho�q�[n�mo'��<��o��kobu�����CxZ�'��}�Q��V�:��3dB,=��:`!-m"_�T��V��V����,*�3@5+$�A>��$z�n�ܚm�
=���l��1�5>dC d��P�������0�c��+��
&ɏ��nj�<��"�Ƒ�;�*��ː�^<��,.�c3W���>��'zRI��+I�
S���\�$��	�q�ˆ��UO@�r:��z:����4p���1���yV��5�'�>Ģ��5���^����~RFܘ�<�K�.k���9 �����1>ù�/�7�|DN�6�Y���2^��b�nSEe��ǖ�Q��/p"7�.r�99`��.+cx8�Z�QԘ���
��+	7��&�7������s˘�[B������{%���#��pz�px���T.#	ax�WB�N������>��J����~��1�:sQ_0����u�L5�'���썝h�ȓ�SWh���l�\:���7�k\�հ��@�"��4s%�Mس7�t�.`��C�!�<�y��!W����]
g�.���hW��uoX։:ܩy�M���`ь:&)�_<5ffWo��9!���\��D^�pQ I���xT�A�VʩtJ�4E�lG[,���s�Po[�c+�!l��>C�I57.iVҙ,VWױ��"�����n��@Q��ӌ��ȭ��J!�f���/� �-�l
���)��>R8Nd�֎�����X���3;�%r,�����F�C;�6��XZ,ay%��L+�u]�d*���8��a�xJS� ���.4��>#\�	n��Tj`n5�3������E�X̦�֜�*��N$��̨V�(������	m%x�����eM�9]$�-�V �����#~��'q��,B�B�Q��<Y�G��,
�튣"�Z�vC`'�H�
/5D�M#&��B9Y4�rl�wNmAms?��c�.���}�Vw���ӓ9�#EU�c^	q��:r�5�����?� �{�(��������aSGʅ�K8�Ϲ�َ4j��M�3J��P���}5�-��sM��D5��Ťpx�TikF��U#��c?��}�|ESy�?$!3^
�	�l�/�\,��m���ޅ�>p��F8DK���i��\�;M��U� }.V�ߗ����3N=�Z=�ߍ���e�x�wR��@;݆��ϯ���/����<���sp]������}����S��[E^]^���S<��w$ 6�X Cãz�ex������^���ӧO������\4[��1�#)Df�q�>d7:Ϯ�����8�J%�[�y8<2����߰��a5�<�#��7��7G�M���BGG*�,i�v������|]�\��W&�&�����K�/��8;�2��r�ʖ�R��JU.C���j}�ω�!�$�q���irIH��Ԋ������V.�������{��ɷ�i����۾��w������������;��PƗ��E�򩧕�5��;t�ؽ{
��6�~������u�Q�%S��w������AO�\U�assО�o0��ۋ|ˇ���=~��ić���D
��h���Q'T��.D8R\+(�������(m��+�a��I2����${�����ě޵{&���}" ��R5>��ݡ���(�,$/]��������zFH+Ӂy���
�����'�\�gЮc~�D'��q���	���7j-,�/aeq�3󘻼�#Gn�;�y�F�?�y{�2��h�
7>�� F�����w��V�BQ�:6��9���i�S*�Q��ht��ב�����y���!6��S�i& �xYH&т�͞��}��aű˹���A��pS��9�o'n���cd��W��_l���ҦޭV�(d0�e��|N�4VL��8z��wxQ(\W��/��iCn�
���߫086e� �<���B�:3%x�T��u��٘��������z�u�U�%9��G"�M��g�� O��p��Ff$lW��!&�	A�L�]O�4y{t�*KCȢe9����AT<HX��ц�5z�s�a�Ɛ�����NqzS��^�˃"�K�l�7�Mo`p0�����T�M~�~��-P�����{�/�"[,����E]�B�s��uHcAp�L�����I�����N���BC��5��PؚˋLۉ���������iX@��+�%�/��nt�[���6vp�w���`&"SVc�5ˍ��{Rq2�k(�3@��X0����;v�@��C����&D����֘~��T��Q�k�����j<�\gt�����-�[h��f�ڬG5˾�?O��E���".�=�b��f�z�p�4[���n]�P�X�ɭ��B�%t�����&�bl���t]�h����@�ƉT���L�5pmNnG*dޯ��h,�H؇r!�j���?�T8��\<s]&OFZ2�#�w���F��B��3N2�c��m�Cyz�S[Ӣ���`T���j�/g�d2e�ll��O���Ė�´*j    IDAT�CS�Y�VM�@��
ٰ�.�|V6�u�y�2��
ES�Ky�e����F�06:�h$ �h��<Ξ9'�����1>��
�l��x�hz����gj��v�";�;v
�?�4�e��/Ӵ�kV��v29�(������^�6G��mL�uOX�i��'�Z)(�rj|�r���g�!p�ڨ��Ɖ�M��DUm*��{���׉z%�����s>�G���>���3.�駞E�\7)�.f�0��%��lԩ�26��6z�dҸ������X|U*%Q_���4����T�#m��p�D�Z��\�o_~/�|'Ϟ���G<٣���V[�X7j��>�[�z��Lo�@�^���E4LS��NH�&�,����m�X 4@˿�nR�Ʒ44����7���[�2��h�36��)�ǡ��_�jU�'���c�͋'P.S�@J�5���ކ�����=��S4"���Ǐ����_|M
��a��m:o�_�y
�BS;@���/�ƌ���8�K�}FH߲,g:+cS��׶W�]����Gv8ġ���}���!���ׄ���e�}%Ӛ�ź��i�! ���\A�,ꐱA��ٲ�}ޛ�7]�ܩ:� ������Є�����k�d6uЪ�	�Me�+�qш�w����M�S�gW��zx��������~��`�����\���w1���~�Aw0r�7����;1<��˿{���#x����ˇ��x|A��[������@������%�����F��V|����`*�r�lP�C�(�i�Ɏ���b���<{��mG��6�,v�)�'O�Ⱥx��|n� ��)XL�yk3��_:���E�6� :א��mbh�(��ȇp�}���H�:�b>�qΣ���Y&}�i�Y�^���g���D<�j	�G����(G]!x-$��(��h%.lf�P(䥅�U��>��|��_^\�����W��,b��V|�bpx���w�������
�&J�6j%
���">���)8Ca�u�����V��?��=���\/VP�WP���e4�.�Æ�虜8�M�#����v@�E62�M!g�r11���!���t��S����C{q���E�Ը��|N�����FI�Sv^���uJ.mɑ��h?��D����Zg簑�=sP(�f��W���`ЇP�$r2ԅ7k8A(�����|1���F��9n�q�<l(����@�,y�}��޹�h�������)_�#_丙�1�Չ�� ��Y�u����6��� RL;�dqנ��*���0���ۀ�Z�o4��~�ʴ����fVt=���]�&0���f	�V~ҏ��6e��L���2~���`u3�p*��v��W>�qs�!�#���A8�П����L�bOκ��X<7��C�t7�����v�t��.�p��y�={	�2�7N�YD^3! }Ğ���kt,�ݚ��)S�`B\G<�E[_G~3� �F�����~�ޡ�ט�!;��R�(rl�LH�i�,J����Z>9������R6J��h:���lz-�x�uz|�}pO��I�G��/]B�I��0�&�"�H޲�5�󛇼��n:m��k�e�I-��@ۦ��pJD�\''
,�,��/��M\Y������F�$���hPS6�DX7)(C�p/j���2s|N��ˡ�BJG��E��A� 	A�o6�6�T⡫��-ݻ��8��書<���r�Ed
%�|'�c^���q`�{��j�Q��7�������tQk�Qi���)㵓piqNwP^��3���὘�:(n<��g�����3���?��^��t哟�gqi�2fg/�Y߳k���tO���q��@������8���5��B���׊�	LPO  �5����D�bu�1t}Y	�l�iM	J��ڏ��>SQ?:�,N��C"]��7M �n�ۦ�`�ǩ� "��Ѹ#r�޻o��>rF���>��&���s����/�x~�s>fėlT9b�CWCy�L��I)!�QӢh���U�A4^<{�,����ajj}��W&�L�޲e������B���x���;���h�b*4Z&00T3BMM�T���"���+F���`�GڅD$,
�Xvфö���i��~���+���g4S�I�Sށ��&0�ͤް�<��A�О���_~�a<��+�U;Ңx<N��WJ��2���?��w�P.uv�����W����Z,�����+e�K����5s�
���>����VG$�B�A{`7v�+��%��sp�-��ߧ�ZOOGo����g�e�ʵ&������3��p����%.�������mj�U��� �v0_\QWnY�k
�|�d޾$:�0�td�[E�V
�ǥ{7N�&k�Z5��Z��Z�e�9A����<��W:朤���
h�ӫo9<�~�����o�]�WuWb;�����/��W�<7NOo���p��7����co��?}?}�I4�.����?��n9��ῧ#N�p/J�'�w���m7a0G1�3?�V$)���Á�ۉ�+95K�.������[N���`�S����F���7B5��u̝~��_�UJ#φ�K;1��X�`��m�̧���~'≰B�<ݖ�N�&=��_L^$�j ^��+�Σ���`7m�8�Q'���G~g#@Ȃ߹X������ؓ�:��n�r�lk�k(fJ�Ɲw܍���aaq�~�wx��XI簞+�Tn�\$�����r��FvDbh-��yC�s��f������Ppoہ�F��KH_��6�rF��p��J4�E�Eϰ|�U���ӡB�@� �Z�b�i�1jB`	�<��.�ȳ���p��"9>�| ��ڐ���Dg^��2�؃�-J�&�M�k2�#�s�P�|_���W*�]�)�d�D�P�h�I�!�Rt3���JQ0�S����K�Ɖ-���BUN'D�kB�>>"��P硞���t)D��62��Y�����R.�����_�	���[Z�+\SK�"n���#J�J��47_6\S�[F�X��F/�VKt6�y��{رm� P/��*�C�V�HӁz�%���8��^|n�;w���#��LF�d"��.�Ue���j�;H�jiã=��<J%�<��)x&�J�3��a�ٔsp��<^~��lI���X�JZ��\_�gs�D��6ȿ����"������ΐӌ��U��1���F��سCCC(�Ş�x��rö)@�im�ψ�}ͦ
��6~D�E�*j�N�DꢬyMP��'Ytq��nh�bk#x+Ź����<���bx|�����Y6�M;Aנ�lޘ`N$�^+ �a׎ql���P~�~D>I˴�N�lҰ��q![�b��".��au-�k�i]ۺ�6���W�iU0x���'�a�����pRi�]�h�؆B/kҪ5Q�c��p!	I������π��K�̮aee�R�+���E"�'�g�IVvtʨWr�F�m3p��r�ZF�>� :��(C�N����e���䙳!l�06:(����,!�x���XZ^�p� <�x��Z@&[�������6�];�!c��[H&ӏ�.:��Q� 'N/��Nca9�;�h"%Q�ֲ�M0ދ\ZsnKx���ʂ�nC�����ٍN�kM�(�MN�C^x�uחp�cj8���� R�8�!����p5���ݬ�I���^������?��{�n�E{��c�?����N3ׅH$�R��b�����r:�]��j_Y�	�i��n��&$B"ޫƈ������#��w�n�|��֭��ڶc(����O~�=��\��y��=|����^��g�	�����v�܆��=�DBx���X�����3�BBʭ�$)A�A��I���Ɣ�]�P�pP�H"�&�i�nx}&�altw�~;�^D�G��	�!���SO�N�+���&���NMm����O��w�.G�b>��_�-z�!K(\A�����-���[u�WVW����N뺳��ԚS�f�	�=��ƍ�[�h 3�����GNh�b�%�y�8w84}  �YK��#��#�`��]����9xֲ|���Մ���:<���Ǵ�u{h����چ�j����x�ɳWu�Q�k�ѱ&�T��^ty���L�/�:!��>7��1��hh4�/䮸g�1�%64a�����j~����]Cuen������?x��rǑ�����7����>���_|����}���{��Q|�wcߎmp�O��?<�~����R�1�k'��N����%TJ]��FP����������;�%�앃����7Kx��2������J�I�	�ހ-84�*��s�M�Сgw:��f��E\~�V/#�:��U�7��ti ,�	D�M��=���}عm�v�|N<�H,����6�/�����XKo`׮]�6�]y���A�I8dUXd��4N��~�������4����PC��b����'уÇ�`���**.�.b����6D��0��յ<f���5l�pG���������-W�A�;0�٬Pk���Ku��������l��2��&3!�bT�-.'z	h��5T�*]�6�M��9)����4%N��mzW���<��=�Ć�1;�($�1Q&w�"1���-C����.T���W��b�4;�7��Q�ѥ�E��/�`7�z�h�wj�����I��z����/��j�ShM��Q�6:K� "�Dxɣ�m ���PX�]�4Ʒ�xwr]���L�̰/#�fKʏmG�Ɂ�\����!kH,����>C�D�h�ki����4����B!+��'�������7�(�b�n0�`�r�h0�����щ�����C�B�.�&D���r��uN�7Qz^;:��J��p:,���I�5�S]i����
�܈=~�{���+���_��J�^8�~tQR�09��t�����1��>���n�bn�������Bv3�	A>�����x�Ԕ
�^�\0u��Z����/�-�٢ؓ!E҈���,q!_�Xjj�I�J!��(��e�&���2�g���y�gϞF�RP�50����5q�b�B�]\䴒�Т+V�S����q"@>4Qb�vZ�6'4LE�a����{�(���L�99�:U�rΝsR�Z�-��,�adƀ=���3��26\�}=�Mh	� D�D0`�BK�j��9VWUW�u��Ͻ��������j�^�N��g��{�7<��D2��s��\A,Z�(��
�� ��d&�R9�ρ����c� Z�.X�E�(�)S#MɊ��j@�ZC�f@�\��R8�d:�׃��f��@_-
GF��$;�Bn�W��ci5���%���J�Z��e�u�a��]�A89i�&`�P��"�wrd��nv���j,�KcS�1��T�"���2���}�.�ڶn��ZI� �/����;��u�F4��ڊ������x�R�����^Q��t���TfgN<Mpz̘Y(�g/Ǎ�8=X�4B"�Y���US�I�ͦ5b��ȡ�����i&A�G�/s�G_U9�j&�Z��XF�ۊ|,���_CnuI����{�b��nSb�K\�5QX��x�46L��z�]x�����/�B���#S����O�6%Ґ�DF��%���/S�:�a�c̤K�˭�v�~�p6���~����ʪ�IBO8�^�G4m}N
�+D��R8��%����w�y�Le�]�.�Z�#�ohmE ��}���|��`��U���1LNL �H�5Ѹ�g�N�K���A��^��T�F�<ig�T���`�Y`gV�w��"e��ho	����'{���Vp��y|��?į���y�8���2�����������A�P9#��'��ѣ8{��.����$��bfn�PH����p��!x�~Q�!o�ω��aQ�}�?<�x��}l2�5<'�z�E���L�4���ꁄ�q�#���?��?c���X�$�����;��b	�]�DB�"FnQ�IAԌ��ٕ�k�۽>!P��@:�e�6X(|l���A�lF^��jBM����N���U3 ���P�x����M���d�	;$���&���r��J��жM��ч�|�O���!�o�~u�_��3U�eock���Ň����ك���N͸z�"~��_�ĩ��=ٱ{x���ꗿ�ɉX�sU1�yǑCؽc#���Ԟ��%|�zdy�y=XJ�q~$��7VQ�4��G&�C��.`!�>�͌��V4x�(�R"�R"���f.����%TSk(e��xPE�lV��T2h�@ؼm��O>��턭\���	P]Zi�D�q|��Poz{�d�`�<>>!�OKs+�u��g�ٔ�G���2�#�d�ɚ`��qD�1�#	I����㮻މ�@��r&��p}tB��%�f�pcrc�XY��8�J&?Z��c���p�7�d�!��KB�`Í(��X��`���B-[���I�^�Ģ0VӨ�b0�R0閚Sc42�pM�#��#�v�9����1�"w�\�`d�"];M5�ڊ;y?���R�A�ٛ$~r�iv�~?6��nC.IY�<Hk dD]x�~eVb�`)���4�<u�X,(\��s�G�$[�BD�����}�16q�UjJ����v�	���{�0R�U�@��,r:�p�<����Ȫ�+�4MyB�Z�a�o�s�4�p�*��Ƥ�'�J�Gb�9��3�����L(���
��Q�k,B��h"@�{�,�=����V2 ���ի��󶭛�y�:I�j��\�1�k�C�9�h�V�u�#0�~����w�	1qb@.vŽ��;;�V�Z�ɖ0>1�h<#/��&�#��(��ɎX]Qϝ||<�覭+Nkk��T/�,t®~@�$�T2!X�x4"ϟdY�b���M���Q�E����#G�|�|����t^K���wbu�*���B�M�\o!���q�kſAS��b�b���s9�</<���^q1���..�&�V���S��.ކ"�l�؃��&��Z�(��R	��&&&�����ٍu���W���d	�K�vu�}:v�s�$�"m(�`�^l��P��n�,fجYF&�F�jFd�U�k@�X��"I���nooC���x�6i�3���;��-���gs$�W2NxD�TZ���b��~��\c=B�7W�.�~۝>�54 ����[p�ڄ��c�Id>�®�p��n4���RHg�|}��>��� �ػC�m���_+c|f�G�I�u��]�oC)�AduED%��������q`v��c�����,`"\) �FLxU�B}�
���BA�$�&�%Wܒٛ1+26�jTTc�|LdT��Z�����M���W�Z���.�ղ8��)�͟�)$'V�q	/�RN�j.���߉G?��V�
1m�ri_��?���Q����T%豃^%6��f�d0���Q��v����g��"�sr1�5e����������$��&�+�T6N�z�!���q�����@SS�4Z8��¼XU�"���t�l^��{w˔��������_L���l�-.gxx����>}�s��/Hל�����BH�OOmQu5
<1_�I3������ȇ�k�X5"�,��ً���?�����G��)� (���߉���'�@�D7�*^y�e|��'1::*
�F�E��,hҩ��_��PX���E�H9mX�S�ދ�=4�D����d�aA�����M0���G)���9�^�ի��q��w�/��/008�\����~�x�X�dEL �ɔ��Z�c���HT���H;����)�{�g��ʹ��ȃ����r򍍀�+2�i�|UU%{���T�+�a/U��y�����M!�K����]��we�K�=�*��E�B;6v}���w� ������W�~�4�4��2b�p�ߏmף;`D�\�|ǎÅ6��އ��N�?7&瀚M�}��[ZZ�l����t�պ��Bt-Q�l��L
'�O`9Z�3����ˊ�����ϔ��n���U-�Z]Etqˣ�⌴    IDATW���th�\L�kL̄j4��u��L�ރ�>� ���{���$�i��+M=�D&�+׮�[�='�d�m��H>�NI�����=}�4"���:�-���G7C��%�V�R�D'�Ue�>��BXYɄ����Cp����.�(�u-Ǎ�)$�Y�L6��6:���U)��K��o��w�`� Q� S� ��
�Y�/Nv���m���!_��`nd�XV�`��Q��	��y)OgDv�X.�A��|��$9a4�nC(���U5��B�cqRU�G> o[#f�9!�� `BBK�RQ�:�,u6��Xj�8I4$��r��wd
���n���f���g�3���3���������D��v� @��^+���jMLFUa��@�N	!5�� 7o��l$!#��)m��jH:)VOY�K�B��_���=�
���������N.ﴸ"�`H����zq~F�7���p�L���7����!(t^�R[��ǋd��ɩE�$��Ĩo��=����Z�)�&­��Q�r�t?5����+�i��_e5e��MyP4�Y����$(3�n;�n�L��<
�Pŉ�M֬�PQ�Q�wV=5�RJX�K'��8j�_�w�CNG>/{���Ʉ ���chh���'D��r��S�Ј�Ⓨ��uID5�VI&ד�F��I�-J"\���B���s�H#��ߕ�Z����N�*���n��R�J�J��)�H�!�,Zy،e�t7HA���F���tZ��V191�kWG�ɕD1g`�]=Dp��`s3�8a��D�($p�@U1�;9���ٱ~��z��@	sn3���#Y�X1� �@�J�''q���ilܸ^��8����T
2���9ȖL���;�U>0kQ�7T�D�����ᒂ�X+�鰈0��;�V����Hf�S���XKea�:D]*^���^��]w����|*�l����'q��9t5p��;�n(�t�Y�`rn�^���}�0��C9���Y���`5��m�oCs[ 7�
x��U�N, �����(���"JB�dLyI���&�7j�vs��)��Ĩ֓A�^��v��rv+���rq�X$�x��_!9?���)����2�P(��>6*��S�È<�� >��`��A��,Μ������KW�e�0f1Y�椓됰9~�X�d��mҽ6�H2�)w,Acɼ"ܳ p����	>�7�8�s��I�^�jiD��W�D����N��%5��u`�!P���K�
i��yr
�
��p:��>���ؽ{�\��Ąp)2��?(Ϳ����+W���D$���(��ɳ]�+�9�K�+�����>���`�d@*S�o��w~�#��W�$�3���|�s)���O���x����PTR�/��|�K_�	p�\6��a���^��SA!Js��J<l�h�9��I�&����gB�cc����}�u+l��zA�{��0Ꮿ��Qd���������He�x�?y��դ4��U2	饱 v��A����ӏLN� �R��hD�X/�yC���]� gs3�~�ٚ�uQ�
�T���	79'��r�����g�K1KIx60(�B�'�{���k+;7�|�C���?�]R��s�X��_~�aW{o7`*��`]O��؂#{w �UNo�p��|[��o;�ͭ-B
���0l��-��]�PRf-�2SϘ�e&�*��Ud�L,��ʩ��D��5����z?jƒ@�,��K�w��d$���
⫋�O����Jr��yT�Q�~ld.�����pz���3Ё���8�k
�4�>�t]��B�+�Ï~�c��`۶m�Ŧ��;.p���q$�j\��Gss#��:0�nP�諡�B+R��ˢ�_�-.,`iq�h\
 v'��v;�l����x:�Y���E{{~)�s�KA0zc�T��Uk =�a��È��X�AU�Jg�ҭL���nĝ��6_�����Q^[�ݐ���D�F�C��B�����<��VA�;��4����%$?J���
;:N2�n��iLƅӳk�Ȏ�;�%�,7����''�*�[,h����As��Ax�UuM�E�Y��%*Qհ���̼���H���I��.�H�q�j��@R�XD%Z�i@~�t�D6�A9f
$��vv<	�bW_�
�K��?�κ�4"�t�dڢƋ��J�S����I%��ت("��$iF1*qtwt
ƛ�NvIJ��h��`�X.D��S�9�5}^<n�n����G��m�0��&�#���s`gkݺa�_�M� �8Q���L�x��ͤ>��J�?�� j�ӌ������_3_���Ѯ�&�2��YK�G���y�V����C���Vo������`�@(�����0�Z�a�F�\[T��^�8'�U"!�J�W/�Y(e�5�XI�$LM�O�ߧ_���)n��i��>n����SI�z��`|�Բ���M-���K
�{��\1�VΊw��PZ�vb��t� Sޙ�eq�����{���%P���.]��b�S"�&J�*el�x\f��m�pw<�
|��V�xe�A=�eFg�Fق� �M��7N�f�c��h
`,g��q(o?��*��p�J�J��$�'��Y�b�����&x=N���8!�P6SI����$�&���Kk	\�ō���3�>�v���މ�N�L���N����W�����}X7�֒�Y�O���So�����0��	���T,,I���8�<6nہ��^���^����&�IP��k�p�v�zJ,=��t%����Hɶv��c�4�#�W�6�8��@Uȧ��
��|��ȭ���CO� �ȓ�$�'�͂��Dĕ���(�b,�{`��a��r%�|���FF'��v8���l�������eZKN�����Ę�T�w�܉��6i�,��bt�:f�e@�WG/�Z��s����"��e]5��U� %Mʘ+�P�bg32���o(a��
ZjFC0 �^8�"�B����4�ŷ��<��;v��@߀ȉf2Y)���payyY�t��I9��%��<�U�BnWr�"b�8������᱇އrA�x� ;~G��N�<+Sv�f���N��/c�uR���C�Lǂ����?��P)���DrZ��$��ϋ+;;���ݒ�K}Z�����[�L�'æ����8m�՟t�4�'����06�;��@�>�臥 �3���x����ɧ�������bZN?M�1��7B`}�:����]��o6��	�;��ǇlbSO -��}�75����d3�D(_N�)�%�\�Db(�R2Q�Ϧ&'��A��/pY����&�q$���7�8u#7*����}}��}ב���{�7���?��q����Ó�}#Z6���.x��8]��ہC{�c��A4)SFqAePeuOMiJ�1b�vUL�XHE�J�у�%{��V�[�`�9�LW�0����
�V��p��z��A�-Mhlv�q)�afl#�#������ER\&�Lx�|R�ұ���mN'��*�zP��}{w�=��[֯�j���0��'ß��ghk����%x����&geˇ^�H@�flij������bm�.����fO��
��La~~��>�%�\�~�!��$sy��c��Εqmt'ߺ��˘�ZD�l��ŇΡ��}�;/T��!�) �)�=�b��Ǫ\�Xe)��^�!���E>��ra(&��M�|��Z��*���C5�\��A�H��pz`�AD�5���b2�o�1&�7IA�MC�&��+�?v\�ɤX�����؀vŭfص��j���S��L�H���ǿ�X
˫a�I�H�&e�h�c��ÂO��2ac�\3�b׋�����	�WϏ��$���h�$ҥ��S�ȓ�;�u�4�l�k�"D���/Ө���hp7��f"�͍��F1Oc" n���%�T�ł��c�RN��p;,�nmB_g�$c�J:L��gJ�3vk6'.�����02:!ʺ�M2*�����/�dԣWP�b��UQb�,�Ѥtg9Z>G��I�Y���S�Yk�j��,�Q(gau:WL���N�4Sړ	�U%�#�^��Hp���-AT��u>w=i�JQ�$�"�����]�F9���}�A�*�XJRhr�zA����%�=��1�� ��8�I�TfүQ?4�C�w�œ���*��C'k�V�-?���U�����M��/�p�uV(˛��l\׉��6�����D��jq#+b||sdrLX,����K��,�v��'R	�j�k��D�	%pO:&4�9��D[��X�p�aVWdXaqm`r_�O���ձI���)�ؿW$>�\&�0���1�)�f��MA�r��06	�ޤ���22��t�U�=	�c�0����}&_�P�)6_ʰctz	g.�`~E�x�o����#�c��	B!C��^������wo����au +��\�����eIV��=ر�_5
J�S6�$�P,�l�:�v��Fk8�1h��&*/�}�LQ��6�@�s�΍�.��"I
�W���pg���+�(�4U3ِM�D:�m3�����^�!���a�F^"��i��x�Ĉ�%Z������{�;��>����`xNo�� �8���	��W��G?�|�G�q�����������9��$Dy~&�A�(�╋XX���x�AI����Ec��v�	�ㄅk��	&�4\�=��o���H�`�T�8����'|ʑ�ٗP���2«�Or�}�b󦍈FC8�F����u�����%�ޞ~uͫ�hll~���H�hL�O�A����f0r�J#���L�Y��+��g��c����C9[��(��_{_��7p���f��A"5'���nç>��8x��{�U<�կ��ٳȦ�0[,h��(��3e���ø��z}b�7!nNg<T�S�,��|&M���J�q�f).n��i�I�,$�LOM`qq��_��_"P߄p$�o?��L��4���o�M��`^O���B�1��5�@�uȧ�M��"��P�5������
��s  ��*����꽴��k>M�Mżx��h���K�O��Jk�XGQ�\N}c~��W��-/�X��7������R����/����E��`o�Y#�]N�Nt�{�#�c�P3�f��i�~��#M�Iv:R� �)ae!"�*������9Oť��/��JY1���J�p�Ri$Rq�+9�7�aÖ>��86����q��65��\���$R˓0Ը�I�R�D6�S�)���.%����$R�{��}�#hooG����2=3#݄���e``��꤂f��BO&R�0�DɅ��Dss3::�D堩9��Nk!��	I��/c��$OT]R��!6=������!��K1�N`zn�ύ`lb^������R<#�4t�c��}(��OQȗoUD�X�V��6�	�(W1?:���`I'�4��B&� �C@%-�Cf3;�twUP en��.��h�dC��;qv��8d2P�����~5�b	Ԉ�5[0��*�!���B����
!W�S��ps��u���M�dsk1*�j�YTةgQ��v�LQ�H���)��)Yo�͓��ʝ�A����3A�"n��#�#2)�4��X�f>�THF�6�aM���������LHHٚA9,�XUY�#|3<n;~p9l"�⇄�|� ]�W#Q,�C���ɧ
���@WZ>���)��Y�d�h�B� ,x��u���1>�Ϗ�>lڴYK����&xYMa,&V�b�8N��.*S?���0�S"���*�L
1�Rqم�L��8	4����r(�ePٝ��������]qv���DH�ZH/��I�$R�@Wҡ7<�x��T�D
�|�MMqd���Ϗ�]��!|(��9��i:?A��L��G����[��25���CU���&�R\F$���*1���ˇ`�Id�+1+�4RK��2uRRlXׁu�:���/
���b�ӌ�����	��xvy�(U3�W�9,H��Hgk�;d���Eh6���n�$����4���4kk��~��Har��H�
(,��+8sqo��$r}�wl�ƀfC^��UY���N�A�2'�����|�ӭ�JB�&��J��u#z!�:��u�a;BbU�"�E�Ë��(�^����Y����qx �nGO�G�L|�]ÅKQg�a߮����B8���c��%k���܍���@�[�Q�O��Fo���Lϭ"Y�!���h��_�
��)��?B�y��ę���B$:)~PS2��0�*���S֍�"���\�BV`�TB!�>��b6��g�����J���e4�YXb�c�@�(}U���nkQ��*P��i����XRX��sWp��ψ���,�[Z�W������RB�t�*r�em��x����t8}�mqۍģ�箻������l�������я~$��=���$���$�I�f�)?j�{�`sX�07���l��o��fl|x��8(x/#�čݻw����O���.S1~}��ߕ�G��	Ŕ���ʵtw����]�l�Rxr��[g�g_��k��X���f
y�E�00Ё'{�>���F������s�.�I2+�ӕ��"�߉O|�q�߿SH�4Z�կ��}��v�k�$�G�gVIf�:��^/�˚���a�ҍ̈́(��9��K��O@�Z��kE��7!�V��c���``�G�Ŷ�۱��ɧ� ���p��4��&�k�F^k�R�R5���S"����ޝAq�����f>`����@�a�	�}���ҡy��)��)�B$L�/�+�zY/2)�{"&s�����D���N���rBOc�Jfmn�@��x��������!��^��O���ӡ�aw���Zf�r4Dk�j[;��#��s��tU�y�Qcg���7p��<��>'|�4[���!V��:9��ٴ�M��6�&�k�iL.�I�F��LR\\;�����!$�+�.cfb�Deh
	�w5��K��hne&#��xت�tCs��.x�#\�~�w�y�o? ҍ����я(c5�Ǚ䳂��}Z�����<��ч���$���[�lBOW�@�l�XX:B�Ț!:��&���N����8���XV�*�Vĕwdl
�/�#_��O��"�_�"U���І���x��͏L(�ɱW�x�M�=�Rd�bj�.���Z�$�"�,*Q����V23	NS����KB1�;5Jw�I&>�n��@Ȑ���w
����M��ۂ`vn^:U�ZY�!;�$#�.(Jr��+t��z�h	֣��>�C�޲��t��i���S�]K��;@D�+�XE�Ȍ��2r$1�*	��3a��T�@I�fg�U>Iv��xX�$	SC��k+�n��c7[��eEs%9��Ś�$��$5Ĩ��&Iz~�����Ex�4��]�\�T�dR�T�lV:ۚ����^'�,|N�V�����2)����0�W�8-��V�C�S} (�E��M�=ݦ6Ԇ�9���
A�d4�b$�<��J���_'�]�b&��fZ��
���8幭�����Ĥ�xQ>G���ia�HWS�1�	��ߪ/��.5����/ѓ�=vC�U��V�[ʱ���-�3��	W�$W�|e r�T��,�7IM0���]��p׭�wJ���߄	�Uu��F���E]I��\N�)m"�)e!���j�6���Z*Sa%+� Z�4�91�߂��&�fdk�Ob�֡\�`j"����XY�(7M�e�2�L�g�JS}Ë����J7%dRqx�fl[?�ގ&��@�i��Jq4��ڧ*����f3bi�G�1�ǹ�ゟg���݁��Vt���p�d�=�@"Y@���V(��LF%��ǫ��ب�b��O�M"�;v���UVi8��X�~��Ҹt}\x[$s�l�0�������,��$�før�
�=�c�V4)�XF,[���Wp��b�6bǖ����ˢV�Y֜TS	EҘ\�ڍy$�8�]BM    IDAT�0Z)�L�#-y�r�I9
��*����ݪ l����,��7S���`"�4�t.%M�5��шH��P����+/!��
�6i��r�6���Pn����40�R�!�x[M���#x��?�m[ש"�?������3��g��ć>�>��G��R/�%����Cb�c�zrb�7p��[�|�"ҹ>�����O�:Z��Z�V���/��^@,��{��&L���8	��LS���d���I�Y�3a���$����(��g>�)<��G�v�P*���˿�׾��$�w��R�S��۫�x)gY�	oCrX ���K_|
'��2���E�x����x��G���?��_,�����'��O~������OAh�H���Gp��^|��Gp睻�Hdp�̛x���091.����Q  )@ֿ��cr��?���c!����Vdn���K:DS5'T���d���F���{	$�f�R13K�*��������y�c0���/}�z�D�i���K!tJ�����zgS��	�-�K�y�o!�,bՙ!�F��Y|1܍
.D���VL�/SU��x���ffIG�PNFa����3P�g�1�$��1�&�E^��}R � �B��:���{>����;T�����ߏ>��J���� i*�TJ��-R�Y��c���.�}�\�x	�j{v��Jh_y�)�;Q~�T�����;cxp
i�����X�N+L�6kf2e��5������,2e�C�z������&�>u�r��0������`�T���G1����gQL��\��d�*�;�N&W<̫顙F����÷�Ё}(�3p9�����ի���3O�&!�^�AZ��6����(��j��B�����@�t��Q��`m������GTA���/��%��T��aq�(xaq�3�\ހ��G�Q��[��2��$��&��mD]k7���&�ǒ)��Y��|0Q�����5,^Gfv����"��a4s_P�J���P� ��@MѡYMY���bRV-R���#�Q���#��ӽ{�<� ��XX\{s#Db�U��;V4�'�y��8'A��b�]�A��aag�p-_��4�%��C�hD<�)J(����������t蕻����ٱr�35�.��92V�Lu�u��l����tb����N$�n��+:۪�t+F�	&1�"Qk���I��C2�����$�|�(���j�Tu�'�.��ь��4xB$ʟR��ԍ��$���5Xqq|Y:��BQT��E��3�6��r*Մ��L�����$k�\�v��;1�ó�cg��v$�xv��I�%!R����R��$Q�8i>����ȸL�o%Q��ўUST�F�On�GhE�~ 	wA3y�� �%����4����	8}n)�0@>���H�c��⇒�c�QM*t�J�0�R�
iPS�R��oeQ��a\�L+7Er�d 	�s)�b�����Z�	z� �LJ��[~@8L6��"M�x:� 0Vjp�-���@w3Z��i@&F�UМ�$k��
a~6�|��σ�&�@``-���{����0��WV�8��I�=v�ݶ�*���L!�2�R+���B��U�	�R�B�+�Z��j�X
>����a��"y�$Le3�*ɲ4o�	f�kN�jf��&��:g�A��ɁQ��!
O��_�V�&����_��Ĝ@ٲ��n؀#� 賋�%u�/�-�¥�k��;����ʖ�8w�N����Zv��� n۵�=m���
���b���,�8w������5
���1˒��!*)��X�]Y�U�`�O�x��5l8XlF$S1$3q��ɕM�,Khh{K�Jo����'a$�����J38%#IL���j@�{�FZ�Sµ�C���ģ8�o�d�L���p���p}�4��h�����L�DK��W2�M"��\�g;�@��%�����H�{�{/�˟��:�d]%�i�8~_y�@��Z���Wj��T���X4�HL(%'KN)���b��t����Jgd����9�ݻW&��R'O���'����Il߾]x�����E����P<�섳111��}�Y���)��Q5Y
OG�P������c���=#b�<^>~/��g�pq�f���B�E�wܾ{�Ql�0�����_���2����|a~�{9z�Rr���I��)��:z�87���	x�>y^z��'�z�;�K����,�dƶ�4���f&'�c�n���/زu7^�����~�H$#�sy��J ȧj�*gu6'!$��V�
�ќ4�U#�?�f� �{�+8<~x��a���h�k��>�,�J��j����W���J#Y��>�H�L�lV�/h��?�[�i�7�[M�K�4J���Pw��>x���N��c[����I��]��(�kȗ��X��f��fF:���˂�� ���n�$����ۿ��(�p��d���C��w�%� c�R�N�F� �{&R�XF(U��\c�i,�ʈ��9�v�f� _�b-r�`� r�8�]��ř	��!4�,@:���K0��2!��h.pX��%��j������܉-��1;5���i�w�������҈����{���tTĠ��.Gmbl$�N�9Ew�*1%�R�(���[����$����䏋���<ߗ���L&"���M�|���P�.����q�r$�91�A"���,��Xe�M=�a�>��E3HĳHf����5`����8४N2���iD�gQX^B-A-�TÀ)-ң,�b��7���UH(��	F�Qk�`팊U�8�z� pl0���m߄w|�!�|.��	���9�fAŮnUU��pJ2$um�q�$�Cr�͂&�5��Q��c$݈��3��	Cz�����%�`��Z*��Y:3�Dn�$$�o�T �]�l���y�D�\�:H�s-����ʁ̓KW�aA�u�D�K��$!2�Xt��=�{}�`�n&��Y4�.���'YD#|�Y��q�$�T]��8�g;��(f8���廬���0��^�'R�⺴��]�ʊG��g�C��6x^7'1�mUj,�TrR&ԫZFP��*�4�E�U��f1�q0����3r�W�@T|�	3`�����
._��J�\	�� ��D.�k��%�*t�֭��>!��f��w��u~L����ؘ$�A����F�E������XF�5!?	���aГ0�c&Zͳ��$M?,�^Vk"� ��̥&Jc^�\za�s��p�V����n��	��l�Oe� +#'�=�}�"�uv����WP�|Zby�d@"������V����׃M[��UdKE*%,�$qedc�+�:<����f���я�[�a�#k��jLU�Y�k�Fv�Ua�j,&���ˡF�q���� ����������I�$J���-Nl!r�b>�N%��%#,E��o*�M����`|�l8�	A�i)HN4�D�3U0����D5��%�عu+�q�>)�f5m{��^z�%��1���Ac�W�<B��}	���(���QY5����"����h��	�p �+��K7�!_�?�f�Dk;������%e�:���V�ʤ�e$ɂ�j��jn��bq���YX�5x����#�"�Jh"9�`A >���b�Â�J����%�}�A��;���H6W���������Hz66��Ԁ��.�^'k<���4�>(��	���r��H�dO������������X��/���B��_�?��'���.qTȱ.���<s�7���%RP�����$r��(���/p-楓Rtuw�����7r:쒛HAp����{��|�::��#����Bdry)fX��wv�qh������q��P�nQ�aA��݂?|�1|�#@�P�"2�*��'������W&P(�Y�,�\���A|���Q�����c\�r��:��e�ຽz�\'?���?jڠ����yJ�x^r!�g�p��>_+�q��S�Wb��i��FĘ+��<���D���M����p�{Dh-��_9��(l.��%�Pr��3^R	R��y��'<����M�, p���oE���� �yzXQ���v��0 6��\L'Q)$Q.)�+*c^�K�걛��N�l�kh���@�R@%�6����o}`�O?}���S��������_O²��Ԅ�YL&��~���L,���l6���{�/^���|T0��Y4��}�>ܶs;|8I4dG����i�A��	�\L`t6��ł��>Z�`5H''�M���[6uS��]��Kg_�BS�	K6���8��E��7�`�T��#��@P ɡa7a���رu3V��E���С�ص{����|W6�ء�7�d���~>���2�g��>'tG�4�I!��t=��W�(}��ZX�gu9$h׎ݢ�R�"���c'p���0�=0����#��A�lB2W�b$�ƮA�o���E8�N!��ưP]��v3�n;�6
��'f�� �V�| ��F�A#�b��M̂�Xm�������vjf�W��@
��d���q�R����]�:�t�s�tIEI�0��D�&���4����C��`��uU\�]�smfS�G P'�ⴡg�Y���(�t�I4I��lN �BF,W�S���aI�v�]�v� �q�`0<T�#\)���L"1�L�x(���_��Xt��n�HP�O.��"Q)�8�11ɏ#�%�,ȃ`w���Y��ES��,v�J������؄Z~��M����E��.<3�v���d09�/ٰ��e @�2�b���F�3U�t8�t�4wT�C�j�M��X����	7W��O��TOqK�!�hqu�t�!܁b�[N
~��	D�Yx}A�NK�"�Q�	!�P��֤[����ū��H��>���q��~��v���g��U�^`)��t�nr��4�8d~�I�ӻQ�$A�\�E�t�Y s���,�J����?�E�/��)�+��D�k���I�E:�2ANg�PŧS&4�BNK]m�6���C� FY�l	�3��A$G��Q�?���j*J,�D��\g�\��|
�:̄������{�m�@�O�.Hϥ��F���OL�=�3��Xe����kYL΅D4��a&�=�ص�M�����-SńqIA/v>�Ћ~�
�χ\$��>{Q�8�>�	9G\�*?�Z�lH��*��n`jn�B	[7o���[�s��zʕ*���i!iڻ�n���*�-���z�$^?y-m]h��9g��B������@w;���t�X�"������Q�4�G�L[�x�3�:�\q�Sc����Ҫ}��9�=NPѫZ�Љ��&x�lk� kkaL�c>���%�&��aw��8GwUY�
'DL��me>@j����n��~�|�?<���Q� �?��/�W���C�`�{���ߏ��V9Wɩc�X)�(hJ"<�LJ�I���G�m!��}����?Cog�@C�>s����o��8�e�V����|&�.]���֭���"x"8{�N�<��Z;v���M��at��y,.�cÆ���R��+e�:uO=�N�:��"������4x��(	Gcr��t�a��M�Y>����wp��(�%�L�yru�����x�>t
����������!.\�&'�|�)����m�.ix�u��ˈ�W��l�s�M:��˧ϠopH�<�������E�n5���Ƥ�ω������o'581VE�ݽ���mS�w���آ���j�i�p+N����oC��p՚�tFd�)��u�lZ�A�!�ߌ�5�ݘ��o���M���&b�����:�5�#K`ee&��� \M�8](��Ȗ+�B6��&&��'���Hi�y8m�wC���^��8#�����Z^;����lN�.���
��Ԗ�ݟ}�{~�ٻ�d�.����wS��wN��篿�L�j��l�'���I�X��b��hڐL��m{p��Gp��9}�i����u�M�loŝ�nGO[\v3�4qXa�*WE'�H����lW'c�K#5�dpIA@�aq�#~��~������+W1r��Ut7z`�&�<q	��)Ԩ�c�Tr�Z׌֦V����dri3��;�o��X��ĸ$�w��Nq"��ȏ�C��kmkFWg����"�i����v�qR�����i���XL��(b MV�@ilB�
��vm߅]�v���M
�_�t\��*��V��C�bez8�۾�v`)�A*gD4U@.S��<�&-6�U�k��1D痑^ZDum(D�R(� ��	9Qg�8X�j$��:�]�����q;�YgA@Q`*vX��,�jD;�J����;����G�Ey�ȟA�;�l��ž4�A,�I�0��L��CbJ��}"[�d�N�7���UU��Ē&�����
���+Ja��Q��/	";�<��ꋺ����d4�/Ovcu7G�#��R`�����.3�%Jk���@�F�@��H\=���N�T��Mf��0�#	gs�b\������nd�K�1��9�$��*{W��r�R)r�jE&CGV-���m@b���U9���81�5O�����p(.u�Y����nB:�(���+��e�D��ؔRa�[4�& ��Vp��Y��py�ů������&���֮���$>;~>v��?�������F���nJ�Z�vy�GT�DTV�DDi��(� �����~
��_�$q����ݚ���k�n�^���:��V��^��A<E"�{wg:�Z�2�{�n���p2Wʣ�O"�b�`{�`5�d���I�Ǳ�1�298شe3�&�44��01���ό!� �ƀ�!����ni��MC�mi��Z���"�뀜��481)�J��If�(�������arn�Qd�8,tb�^4x,�
��:d�A�J��!���m�
�Z%���
�;)σ�����XD(ia:�R�\H/Z�L��*2E~6�*nL-����^�lZ�����r;��p��eї߻ewܶS|R��ȕL��{WF��c���Dts������z�]����ND35�X�����1�����b��@k��Zԓ.�J�<:4T�Lo�֘��P��:�7k�67�pS�~���L޸�lZ C��y�e��,\Y((Y�2���]���h��{�a|�Æ��g[_x����~A�\�=�h�lXMoϠ���e��T�;���}�)�(ɥS"Б��ݎw����C_W��}��I)�Z`�:04����~���yG1
���7������k�n��V�?���7���] x���{E��d����J'�+_��l�BgTKe���x�O�T���X���.EC{�2:�c�Y\^�u��ٻo�pΞ����~c�pz`��NƑ��14ԅ?|�q|���%�4����_9&PB�ss����y6q��q��mۄٹI\�rN��Y��y#Jj��wzb����/=N���
J����<xPރ~To�qR��5���).����M�CP��H���E#IF d�fS�C4�@!_E[{/��zē9��/E�ٶ�����Ć�u��=oF�]N(���k��_����9X<�0��}���8|��������b�F8M(�(��"�J����]w@2��\���x4������hn
�I!���	��#��4��f�����#��2:���
O�Q�ҹxlz����>q������T$�������o����/}��o�Kƍ��z�̪+��A�:.�\
�M�X?<(���	����������'1Ms�G��[6��ÇD�i6�=X�z��}=�8��fE�FW��^[ƕ�(R,��`'#���蓴aur�R�ьx4���9��O�i*���S:��k�[G��T�����Jx]~Y�\�R��-��jÎ���a~vZ�-��.�*8u����I	@�䲛��"'%���hkMbnn Ը�uB����+���߹)[�� Z]Z���,B�Q_ZB��uuX�~#vl�%Z�WGn�d�!�7at|��O#����D����<    IDAT�ܴ�k��a�!iW��55%��F��G%�G>�Dry��
��y���!�*qR�a2��H7ْ��@kK2���&d&l�$��CUMjb�n,��m�َw<� �u,���c'#m�N�e(Juꄛe��H�	��("��)�aU;�,��1����]pk�;�4����#$���?t]��nu��ɩ�|�K&�Kͪ\O�T⯺�1Ѻ$z2�]=qf�eW�E&��k�ȣ�M��&vQ�e�seKT�����>��Y���y�R���Z!AOafy�ʕ�\R�3U�l�յ(����SEp�3����,.���pJ7��{�'��-IK��Eau�t�h>���=Q	*� Tn��� ����*P�h�]��tlI{|�ʮ^ܞU�MDi�j�]�c�B��E��B.��>��g1�<�(DF}�t�Xq��].)8bVE��ܳC-
lhhR���ov�4���n��?kdh�P�z�u�/ Gl�2�ѧS�f�N_��� �$��f':ۻ���$Ϛ
N$��J<+��^�����uaˆ~����ͷ�8�d����`�$����05��k��ǫH8͍�`, ౢ=�ǆ�Nt5��m��e1�KgYq���Jԕj���,X�ep���O�a1s&&���mط}:�0����P̪�,8}�T]k�x��eW),{Oa�E٥�T�xn	�S�@��JG&�B�)O3�����5��ӗr�y����؍��)���J"+q��)���6�Z�T�����2���u�$ߕb�Ks�v�
R�U�{h����z�7R8u�:�V�R$��l�PQJq��"!��9.���N�6��&�Z���G�D)��K�}#aU&3(���4+��~��Jg�8��ܼ�>��oN)���[���N�<+N���6W8rh��3����I�}�?�7��.V��u2����@��L<	C�$��V����T��P������H��k�������>��;�h�p���������ŋ�8r�J#1&�w:(��k��*S�|P<��I濳	Z^���E��M�S���s�}�1>�g�}��:)�a��~;,f��o^~�e<��S�Lfy�|_N	�:;TN��$F��ǜ� 44a���9�m��Π��N��L�b����?x��>X���%�*#���y�ΏHA@�L����t��������!2֬ژ<3��W�ɸ�^3��G�ϒ�DP]M�@��䡇�&��~�3;���Zi��G/�>����dG/~��l:��&d���xͦ�Z(
����/	wR���ط/����c��}hj�A�xI�����<0:6���;.|J��K��{��'�����?����#�<l� 
7*�L9�HG��x��;�G�� �2~���ӟ��+x���§>�0Z�}s���X�ʄ��B����2�<s��<-�.J�%�iMn[��W��]?y��aus����
��={b���~�L�b�`�סfQ
�L.�S�9Lvoۄ�>�!�ש(u�ө^�ɿ�؉c���]o6���Eo{'\6���%��-(,H�Lx��x��l�nx��RX���g�ჃR�F�yqt%�+#�C�߆j,����]�����f,�Nɏ&����C�K[{Z����D�\BGg+n߿G�+.]8�K�/`uuN�CF��L��l�B1/���� ��RE�&
����4�W%�c7{ppP>5�~m5$cS�y�=Ĭ��7��=|u�B(Es�|m�ώ �*#Q 
5��Cؾ��e��Z�p�`�7��1��aV�w��=��9s�7f�M@��(V+��c�5�)�)�yM�ww���11�1�^�DT@Q@Pzg�齜^߽���$��~����s]s���|˧�ŋt>�D��-�䎦_�GZ��t��fezQ`� ӫ� H���E
�B�\op����\�jѱ��T�FQ��O��\(7����`��8��ᭈ����=���$[�
�$i�R�g��*����|a"`W��u��y/�$u �9W�G0v[���$�Х��d�ϧ	+u k1�شu�I���v�CJdv�17'h	�7�{�^�[��"<��6�.�Lz��U�:�Ҍ��.u�V��c@����֩Md`(!�7�5r��&�~d3q�5fM����R��.��\ �Kt�t

�����t���\����\Y�ѯA]C��ג/$L��J-Z:P�}�\�y���b(Jb�ۜ���Ak]�=�й�p�+��fUi�s!_�2�� q�@W� Z;��s�A�u���	��+�0�.K�Z�����݉�:�gc�7%8.ڎ5���]�s4��&��_��r��#�
?��T�%��|�"A�����
��`�bÈ��X�Fɀ�����J�D�t�x�Dh���l�!n�x�6ـ'�ƺzT�W(�Kfb"�˞�8<vo�)u�؈i'����zHKU, �0�i�%�'�<a0$�m"]��mؾ�	mm����EA�*��Tct]9�"{�tj�1�dB��'�L�~C���ۍ��4v�>�]�����5��][V��N���'��;���DN�	 �j�߼,��0l��N]@9iS��T�͹ynm�\�ةS��D4|��6�Y��$v��4	s��D]enG�x�$��F�u����?�e�Ł�G1�|�2c<�4r���9®ql�SF�@eU�L�z��΃ز� ���9���@���O�ĩ�%�T�}����C�" {��a�@r+Ut��EK�Q$�QIZV����I`˺u�;v4�Б�db�+/�D\&���S�E��&f8����ÙsN�������6�xk1�����(b܄�8�$$3Yu��4���0�����U��t�x�a?��v\s�%z��ظy}�����2�cR��p�5W��K/�����K���?��R<����oo��6x�>�����/����p�5��x�� v�G��#?�1,X E�t2�e˖�OO=��7J�K*>U����|�&r2�7Я�����Ĕi��}�װn��pKPR^�U²1�Y���7\~��O꽽�x�õx�/oc�'[���=F"5��"\�'tc��E.��~��z�1,�0�hko5\(KZ�S��1�}O�~��ș<묳0f�|��g�r�J�1��R�B�1�2�U�_�-�`�44�3�8��ᷱ �9�vQ��.�Q���{.n��Vuw�g�%[�`8(�f0��`0�ؾK�.úu�Ȼ"����+���c���Б.,|�m�ٰ��<�$t��������.�O~t���n��/���{�����ŷ�v��
�B�Yr�ƺ�|�������_`���q��N��m�'�ix���^��.3������XB��?�{γ��x2�NpV�b�倏��
Y��N�?o���<D�h=rjkQS���^�ڻ�����"b�$|� jʫ1n�8=$:.�T��������V����M��;��F��v���K	�7�iW2�q:P	���G���|��/�d�14�ڂL�!�"ʎ:h��r u��|4��NdVV��oP��|g̨��0q,F6Ԫ��*�G����[��-9�(R
��#)�P�'a�ԥNK�[�ߑ�@%
�H,fRB>_�P3HĢP;��}n:t�t��v�:o�ZП|��7lG31߱<vjA�/����8㼋�F�7��@4��aFޏZ&�!!�g��jjF����v4�(7�B������!("\�@�=!��X�lĽ2D�c���2K�u��/0Q �?C��^&�>�z-�5J�H�R�M��8)�X����dF�*�q�%N�/��U.2A�$ٵ'e$+Kը\&�"b���2q"f�<��w����ު*�����9�܈s9%w�(d6O���]:�T�M�"I�,>�Q�a�c��.`���c�MU�Fq��Q�u���@�x����9�w2YJ�L��֖"9��~�
��TT�,@�!Ǭ^N�؀j��К�(��i9<��8�30dK�YX�X]��_8NH�&T��1;�d� 3(q(�7�\,��� �1q�3ƢHgG�:rL�i�N�b.YEe@�{��R4���H�L�$��W�ΊH��y΁�(��&���A�-*uP�TJ�c'6��S�g��o����6tmQ���_E�	⡋�*a����s\�Q�	���E^��_���ء���q�v��4��Y�U�>���������GRw:��I1׶�z(�.�3q%w�s�j�y�21xYU�G�V����%$V�	�
R�"'ճ���aAN�������%��חBM�(�Y5��",חQ]����\n�CJ]�x����X2��Ã��!�>x����g�xs��2!<��=c*B�F�Ѩ���8���t�l���L���K�X+X��`�Ɲ����s��H�qʘ
z�"�v�Q�q�m�"����`޹s0a�з(���Օ]�t� �C1������f�g�'1��1�Ա2MerN9a�s$I[�&vJ��2ز���9���#����	�v�dD&/*�~�~�֍��5��}!��7�s�aw���^89:���H���ի1�|L�h"�s�"�_��NnV�UXrt���r��?�^�~�t������S/b ��/�x��)�>�ƴ7;΀��\�D
ϐ�~��)�f�=*�F���}�߄;n�I�i���ٍ�=�8�Y���p�ӧO�5W_)u��-ë�.DIq1~��7JJK�ǟ�����5N��_�[6}���G�妛�����?�0��.��\;�o�~�Y%)*�x�����ʐm��N-yJ�H��!�_%���p:X������s|�H2� �)�F���݉��_�b�2�������E��H.�]u��j�1y�D���n�X���\>�ѣ�h��r��~輸���u��y�X��F���,����w�w���E��e��9���8BQX*O���jOe� �I�!I�k�r���е�uc��x�Gp��sU�!��϶��ہ��J"a%`#Ga��PQ����;���/a�*&\wõ��k�b��jm���z�����t�^�±�^uؐ�Ó��K��_�_�탵�����`���[�ݯ�����$:{z���k�e윳h�0{IMm�޿�%�%���5��wp(��ӳg⨺���w.���)ƍ���K���,|k�_d�#F�a\{�,B�"ԕ�p��q�Eg"pc��!�?�3�����*�2Tx``�'SR�8��e%���n�\4|~�iII��z���ջ���f�ODq��u���E�U	qU������O��D?{Z�G
}M�qt�f��� B�D�>%'	?�GPY^	���r^Iq2K�>c*Ə������P	#�R�p��wD&bfzƙ�c(��"1�|�S�L|H�%�6� &�ڋ��}�Ed�	��!�D�pw:P^Vf*�4���W�ISNA�P6���k6c �CK[?>�b/�i/������Wq����s�I.����@\-e�X�*�f�{�=MMH���(7g�_vB &y:�Qe�ݖ�������Q(�&#:���9����7]}]D�$�ǉ	�OǼ[�A��ݽ=����j2��
���S����Y����[4�!U�YэU3�F2��	cF���]�8r��?��e�B^,B�-%Kx�ԂU��hr�����!gGBH!C��Tt��8h��@2���Γ�g�<�;�diΠ�����vttu6����\yZ$F,1����`D�U*=��Q�r��[h.>W6��U%a��B2u����LZ2��bȩ�{ &�&%� ��Ta�G(EA���)B�@G���I�aV�����/XQ*���k%���B�4K�N�3�y0�crH�ʌ�P$JݕJ�L�e��ބ#�*�����%y�����qs��o}$�5Sw������U�;-3��\���n�O\(*ѯ��g9�Z�Xv���d j' ��Z���$c��'�j��7�.�������=Nҹ������*kQL����	d�rHfd��rr���lg
~���2�Gף����2��f�����;���4j��574u��/v���PUW�4	��"��x	�1���U%p�#!6(yf�ǃpq~�SN��Y��ȣ�c ���F��@,�?����ȍ��:i<��	��t	\�"�,9M���wX�f�Ɓ��<&{�/(��j�̦

j�5f�)�ۇh��G;����%��J��3fOWB��*��t�D�T�@�2�<7l܎��j�t�$�1{&��ڒ�7�%�K��B��I*&\h��Jő
����c��	�3���YDbv+	�J%FVB��N(�a�.�����̲'���b/b�=X�r���p�����!�A�d@��1��k�,�PȀέS�^rz�n�<m��5�O=�2}�	i���b��q�6c:&N�,��ۿ4�X�huE��ȋ�������)�����rӵ���������;��?�o��5u|.��B�v��hQ�O?�K���]�w����������3�>��`��s��������[�!���E~�W��t����~#j��Y�Ze��!`q��q��;_@�[��*��;&�s�Y��U��=x�/˰��5����w�ܤq�q������A@�mSx\��'x�7�i�.��͈��R
#0m�I������(*��<��)��FiY���m_�Chǎ\��tW7�����)�3g��D�k���KLr��M]8��5�T�M7��Z&z,�x<:J���l65,a�99s�P�1i:�/�/8WEe�W���~� �S�ǥ�C����\�y�͗��+/���T1醛o�e�jqY<М��n�����c�B0��ʦq������X�����3O���&��=���w �b�֝X��:�޻Q��d�����q��K`����{�m{����E���xl��ɣ��ew���J���K��t����F����\\����F'����\��3�q�N���;?�W\p!F����eB�VŌx<�C[K/z{��8�(�Hz��!Q�v�1#�H����~v�v��zxH*�2A���A�Ji�GIꮀD��8z�ñ=[��k���Rz�" J������b��jkkPR�IS�b�sQW[��Q	��r�?ڋ��v��S�i��ʤY�`�g3�G�����_�v��S�NU����s�pQe�L����H8,fyYDb���G��8�/V�r9��x%c�cO3>ٸ����i��YsQ=j<��b�F�2��F(8�������2I�t*�:vm��=�(�$��S�|΢�����@g��^Ɯ,/Q{j��]�f�������)�$��4�J �� F�N���n\�p]z��?��Ŗmᒯʘ?�L��:�t3&����~�eśDV�T�Mݐ���R� ��Ϗ!�@��z�,�{C\D��{��+�
AuE��|@��nu����ݣŐ�q>c��y��S�!���=^Ub��Q֛.�Ȳ�aHX2�	C�c�`��y=���<	�߻]~x�AU��]p��x�'\$G�����j�D"�-�H �u"R�s�C�qYvz�p{���4���JN��i<I�Ӏ������Xu2�Ξn�r"%e��ciU��0at���) R+��$Lg�:��P/�5�bDukx}!���5+�nNj&Z&d�@�4n'
�E�:ɠ���|3A�1X�v��ft���܈�--7	�)y-v���i6L�p׵��U��{�^c��of+?ِ&\O���i�7UL�I�浘N��ü�%e���C�/ Ln<�Y��yMX�#�F���|��,��0fT=B�^�������#�Σ��[�Hi%2�v�ڇ�NzP�8$gp���1�b��b�6Tc��Fh��(���X�˰/ ,���w��������7��*RP�V�@�T�ǎa��\6�p�O���{ى�:�Y�(����    IDAT���Y�Yj�p��^�&�0&�^��k-qA�#�/�.t���������^t�j,�scҤ1h��R'%t"��#����D��׻�����ӏ��A�W�a��31s���=�O�P7��9���Cq�W��o<�e��c0�A��т�1Ȕc:;\��0yV�2�Ŀv��^a:bL��{��N�'�Q�&�*7%�VQ@>>������c���s`�˱Τ��y�8��&���q:��W�+.��o<x7&O#�\.�g�y���o3��bǽ��F"
���5I��\�B�����Te��I��v�C�PS����\q�$��|��#���?��wi�~���n������k/c�͒Kn�����C�Y�.|]�·�z+��C��/~�-�6㡇��;o��֭���'�섀����)%A�����5� $@ۿ'N��S�}��A� �WV��Z&�1�'aΜ�ߗ�o,���#�}��E2G��´ic�oݏ�Ν+u�|:'.ي���O>'	`vrY���"�oĈzL�:}��رs+b��]��O�v�[�~�}���^���-�� fd���K�K]c3�(�����b��dix}|缺�4�"��]k븜�<%eY�g��?�k`�܌ع.򠺺�dZ���/�?���sѢ7�b�*��ׄ���Hˋ��TS3<͹s��Ysσ���G�?���7��}�M���;n���#U$1��g;������]���������ȏ�߽�b�|�i=ւ���*�}�}kyk�j���8xL1@oO��-�w~�n\}�h[�����X���xkkˮ����ӂ�.]����7z�����X��G_Z��;������2#����btC�?o6.��L������Oa��-�j�Ÿ�����<��ŗ8�Ԅ`I��R��E�(�8b ER�$7u�0�zB���r�A�޴�B)�rd3��%g8/I�I�bR�*��Kc��,��=�q�P��.t�u�(P &ԘI1[#�EYi*+�d�#~�<mο�L�X�^��U��6�߃];�	;��Ձ��#��NGb���ɉ���a<&]v���UY]eE��ww�6{b��h��F��P0�Gf�#Ǣ�v�&;�c�E�Pɬ�����Ŗ�-(1	��R��C���P"��Z�sVL����g�2�n>������v�ri��g�LaBN�NG�"r%�)��g��R����Ħ��R�HT����j.a>�2�4�^�t�G͘���e�58�z�dBA�L��������C�CQ���S ����i��T}�@���(�Γ�7U>?.��"p�e4j��~� iY�E�l�KyPXDs�ba�ǒ�����*D�ڂ�6�^'�2���%�����g�RI�3�������H��f�I�Ɋ1I1ĉLLs�Im*1���N��X�Pe%!H*�l�{x�Ib���=��Gӱf%-��18��k� g�`�#;6|�5TuVp.��y��X�WBg��=,4ϟ.ڄ*ף���a !����<���!�"j��Qo*�v��3yB�2BGh�dt�D�3n͇i���4_�U���t)��%�nw�o%KKl5ո,��0�8���^��m�$���Q�:�Q�����ߣ�;�t�0X���(�K"U��kkQWc�'�S�X<���
"7L�����y�3!�6\F�PK%v<��(��Գ9�Ҋ��A�B����\ԍ7�BAƏGI�gL$��_�)Hb�a�~�k ���VD����W		��$�t���8PUA]m9�K#���/���f&�y�TUk}�z��ծ{��߮��C�t�СC8|���&��)+�%W(B[W7��܍M͈%h>H���G�et�e��Uե�(���-J}F��hk����G�嶹FcF�Ĕ)���Ơ��A��U�<�� rL$�|��d�5�q}4��/iU9Uҏ/�&����*iS[��v���� ߟJ��P@y�'��OV�Dǁ�J��y��:��PH��.���f������]����&���2��/.ģ���:-��74���3f���L
�2�0K�&�LG��&�^V\�y�=H�⨮(���_�[n��U�2�\�z-��o���u���U������_l�/<��G���~��I���G$�SN���s�UW)���/ŦO?÷�.n��6lٲ�?�8v�ޭB�7���q�R.����ēO>���ujx�5�5!�q ʣ&�TQ��$>���Q�8v&i'^[�6}��'hd<1�\Q�����߸��;�Tao1���X��JA�v�9"�	�W|F|>L�Ə�.�00أ���-��Q���@�,�1�F���g��X~<V'��k`��&"�Ѓ����@�z)��Nv�G��6I�!Q����"�������3$\,�q!�Ȣ,R�s[g3���Z�������o��^~�u��Ӥ=�<Er\ȓbу�4ʑ��6���#I���=E����p�MWcTC5\��zء����>���G�6Cgw�܈/��l<��;�K�d�[x��g��Ջ���*��^�l,|�,Z�>��oFt ���r)�5��1q�X<p��pɥ#�.��V|�.��Ѻ}��~�����o��o�K������t��N�ت������U[&��9瞁�7֭ߥ�����V\q��زy��mm���?P��Í�#�b�gb�8�ט`0L��&���z>�D"|��Q|��n���ȻK��+�nBS�z0��RwݕGmU5�%8��K|���p�S����k�6 5 O�!'8��L���GK�JDJ�5��%~̚=	s�9��p�#jQ!�²�����/ɸ�D��a[&
�\c��9��Ĳ�ʿ-+��fdOy͚8Ɍ���#����F_o7��f�z&"�:U
iڇS�2��hɼ͝i,|�c|�n��#���#(wL�;$�-�^�=-��s+�D�A�#�Ews��E��.U�(3J5�+�S�!���%6�[��9�h	�͆�1�}�*_.+ $�E��#��g��+n���bh;�!+�,�kHL�.�L�3�pV�Ւ�$-�J�=�%�uq�P�gt�,z�ɸ!9)He��V0A�u2�����(�Ӹh�:��"���Ua�2��
��uJ��M��j]_ow7b��8*��LAM�C1�s:�����P��Ug&gLv"\�zg�Y��	k�ګ$u�3!��\��Y�i�КV��Dc���}.���z)��E���lZ�AIq@U殞~A�5�3�ii��0��$;c�}�k���=��zU����cI��5J�	���c��I�Kx�BV�H���Lʟe���������Ҟ& ��0�L6a����G!�$]ָaJ�:8	tS���݃��V%��0!`�$ZVD���t1AR�eU���&�am�Xl�]{�9|��Ֆ�'�Ƽ�Lh��pT�5��DƓ��-�0��cѡ�CŒ)�?�F�:�uͼ��������=g`W0n�J�s�P7�fYY�J����&:�c�W�=��O�|&�H��U�S��CF݃DV���n����,#1�vj�����ćןQe��bq�~�� ?��bP�
@UUN>�d%I��=�zL�d���L����V����"(�q���Q��
�Cq����8������7�y�)y0g���(՞���wt��څx��
�}Z�,�#�
�=��Bn�ݿG\�X���PG�$�|�n�!���G��/�;`'z�'��+'������T�x��楀�Õ� /��B�vlX��H�$㲘�΄�ݪ�K=�	����g0��]�������1i�hK*��_\������� mD�H�4u���]�h:pP�T�^1�zV�@_�҈"0�#l�	AMYw�rn��F��b$�����գ�|�稩��w��)�:�k?Z���v�С�
D��w0n�x|��F��3T������7��M�y��`<��SR
x=��O�o�Q��D<��{A�#�	�����`�6����͊{�{^ZZ�{ZW݈Q��~���ؾk?ମd��&Li���W̟����B� �,[�7�y_l?�������*!�z��y���C"9 H;�,��Ք����C0"r�\9�U a����xب�}D:�oM�m
&�N���ğI�k�&���!�5��㜹g��SNA$Bkg6~��>��n$r)�[�
m��h����.��~���)6��������a뗻147�@��r��ޗM"��^>4z#�?Eyy	|�^�z�(2� �2�Ǐ�t�����>��m��K��e���}�+(d2X�x1�y�Y���ᡇ��w�"������o���}m�YϦ��t��U@���յx���q�U�!�,^�:�G??������~��UB��/_����U�wx}�).�1zD5�̜�3N��Q�%8tl�<�:�X�&&M����N=	�/��O<)�|�[��$I�4��aܨi�(����)�$�t��/{���8ؑBA�e�xY��u���q���T�	z��Eˡ={�m9��V!�ӌ���4�I�J�j6%HK"��Cj�Qnt��I�}�t�Y�@?R��M�V,|�%|��G�(-��ֈ�Z�$����=����a��\V�G�#�(��`X_>�2m�ɓP_נ
W����Ac�(̘9(
����T��^�{L`㊠�+��Wl�K7�wЏ`���LQ�''՜�$k
��EZ���09Ȧ��|=�Y	A�xB@��<rE��4ظh��U�%�_US٥BMA�L�k��y� ��>xp���p��� A'��#�$��$7.>$�2�bB��,1�����$s�_a�Il���� ������� E�-�MYMG�	aF܌X9�h�G27^�����Nt��j�3f����5��`ժO�Ŷ���WTWicf�MFB�A(���r[�T����p��i*�F�ԉL�R#�H-gS}grgP��l`P��0�<?�u8f��»��!w^7y���87q��h��(�if�͘|�Lk�1�7]�����K!��um�yH���E��7�t2W:1�9��6URE="�9%6C�
S%�3$&$�2���/�;�~�Wk��::�dJ�S$����"Q[�y�Hp�~lL������[��Ц�ꮁ�0	_��.+�sg'v'ȾO$-��'JڪAQn��eJD%�2�YY>[ӕ�.�;P�J�e�=�� %)=k |L򕔐6d�f�9r�x0�KC���y�WN�OFL�LrXU���}�01v��"�d٩"������D���r"<�%��w"�a`pHssܸ�2Xڵk�B:�V��R[
�Xq��B*_ 	�L�2?�b4��B"���<�`��ys,0GzO&M���Ic��f�{�^��H���4{�Pz9�`'2+.޿}�ʸ(����B*�p���ʽ����0irM��3ɲ�x/-�!K��N(�!N���'F�+�#�.�^�|^x�r����܄M�V#��
�׃�0	�"�q4�`I���6v���p��W�_��&�T����W�ģ��
�xe���:�7A�u��-�J�z{��	\(il�5WL��18�+U�ڪR�}������0r�X���W�VB���M���p�M������e�E����_��G�HU���/GgW�>��֭_��Þ]�q��はݯ���o��g�U ��_��\r��8ag/���{�y�up��	���:�qk�g��g�1M�f&�#�cD�8ttG�j��=|�AJp�0D�^��ķ�s?\x����=�%+>��o��O7�@����R���&�<e�8��=��5��G�9��Y��䰲�B�f� ��ڬ"ϕ�K�>#=���{����������R8cܡy����W��ܿ��q�����K�p���������������]����j�|�t|���@I[��$��/v��p)΢��s=G��tI[��:�Cͭعw���_��t�e���A���.��$V�ی�_}����Sr����o߉\2�%K��S�<�c]�x��o���oSG��eaѲ�ط�]�*��3��NG[3�#a<x�Wq�u�@��'_ŢwW�b����{����[��]%�|���^{���b�xZ\O�8�ϟ���QUN�T`��_����8�ڊY�L�m7]�UUx�Ex�7�:�t���E���N����8r)�@���H�@9)��i������bKɼ?�>%"e��N�^�S�F�Bլ쓹���훱{�:t��C>5�`�!�>U���4x
��`R.�5�e8��S1e�8�݀ƆT���������=����O;Y"����
���HS�Ƃ�U9�ܨ(Ŀ#߀;�HbCQ#��+`)-����Z�+]���cF�Gq��C9m����
1-����(FG<��MX��n|��(�~�C�Ȼ�:�Z��! yT-]a>fr��@w[ۚ��h��A� FY8�X1$՛�vli?���������I�Ԥ籵W1��*��_�ўHg]<s/:OG{ڄK-ʚj7.�G�pe
&�@^���Ǭ��~,��$+h4j0f���z�2��a;���n��v�� Hf>��L����aax	w3�usL:!bĠ�c���{Mu��	�0�����/79ڂF�R=^�7&I��2�r��&��'X�sS�8d����d��x]J�S����<}=��'�<��@P�����N�H�9�@����{����@����:W%ml�� JD\��k��/]��Xdw������ �KBdW��g�^jY�-e\�T��:L<����"x���}�\�}}=rΎ'����K��".��b���A��-`�%�A�d4����f�ډ�̉ȗ��IE.!��=f����?����]�Ф,�;�EEY)�K+��Y�G#�,7k�#�U���o�[3X�hA��|Kd�e0��(XϚ�0�-ǻ�)�卻l�Tp��$ OiV�7S)TW��;)�R����4�y�,E'�I-��4���Ld�@渞y�#��D�;�-GuN!�D�$�� 9F�{�5�C�V� �I0RI¦!X X�h¸����5��sʐ�����Tk�����ˤ���͊N}v�0q�9��At{R�"g���%��"v��H�AI���`q򶊙��Z�m%
��D�-E
�Z{�zFH��7�o�8�[�b��5�w�}$���f�RRaɆ�H@3&i�/�C��t�t�����[1a|#�T* ����P�
��b��12������Վ�^��eyHX|)� ��F:�3��.�MW�CpG��iç���<��?Z'y���;�<m�*Oj�����g֬Y�={����r�(�|�rt��˩��#GԋP��K/�^�����y瞭�Axȋ/�(���Añ���L�$�zT�WB����0y�ɨ����!�\��C�Z��'��Haڬ���7�å�%��7���!,~w^��b�~���@�K����Yg�Euu����v Į����$�G���V��b��Ƈ]� ��r�L�ŵ�~
����o:��|f/�*���q���1C� U�~���W_+N�`�ݽ꾏7	���y�	%ܐkG�b����w��pE6o݅�7lBssJJ+�!q������"e�inH�^sk>�l��\)���^���8�EGK��U��(���>��$��c�ҕH�S�㦛�n�nK���'�}��S���{��������X���l��Ö�F�ABt����?M��ݸ��K$��ۧ^Ţ���z���_:�,�������~�%O����%��_t.�}��4^����CG���g^�K�9������ �1J:-~u��MA(\���>-�6�/8cG�1�G��Q���?7B(�t*M�h�Ɲ-�r!�����F���5OC��n}N�@uI�~ڏ�����z`Z�D��%>ds����;��RR��ÅT�����8ef̜��cF
���ȑ�x�OO`Ϯ]8s�̚1S]a���ZXoCT��6�jV61#;�	ĉŖm{�!A[    IDAT{Z�5��WZR,��P�����aƌ��2���˪1K�T(.F8�G��	�C��EP'7�t��>��6��ݝp�K.�E��3!��t�Aa�`�b}�hm:���f���J��.u-�����ˀ�T��+����I��/;���(�pz�!�WD0�sp�yg"�s���K*(�_�s`m�6���ؐ!;!�[���8Ye�	�9G#�i))�!љ�VV >�{�e���'4�H~ �$�	7ɪ�����A�9�xV�sUQ�����OHF���D��!��~���[���ꑁ �m\m6�A`+�	*�>; Q�&k)~�HيֳZ���!}qʼ*X6�;�2��B��)o>��Omz$�:�g���䢛o*����n Ckf_�m�f'a�;�4�	��ۉ�/�,�O���xj�G��@�z�}�&vS��E_�q����J |�L��N ���<>�0V��d��I�-��Ĕ�����y^�v��V~y��΃]���Y���[�d��1�F� �FB�C2�c�Ȁ�8l�]�s�Ԭ��D�������vA�,�
 ;!�xuR��@�hdg��&觉��r�Tq��d`���(,��PřfvL8�Y�l�<��`%N�$�M�p���T��ϕ�>K��YQ�X�"UV��^74��q�2-v"�K�I!q���08g��*5��Ò��Kd�!�����'�``��B	L@�"���(�|�Hjb"�;\R�R5�*V�x,^:���.;M#��s\��,)��duʲy�;\B"v�-%�AJ��U���t��çkW!��eL�lN���Q�P7ў�$�g�&�"�Gq$�[n�w�q3ƍm@��^z���W�F��DuU�x(t�f'�6�1�~*Rx���,r�Գ�QaJ}O)#�T����Pp^^V)��Ν����Oc��Z���!�1%%���f%����O�?����
8σ�9�G�\ ���;�D��w���3NW5���^I�2�c���B$R��$���ړ��5z��� �.`͆���bь!��R���p�Sp�_��g��L<��@���o��.�_���?
O�š���=]=rt�NEY	�}�-�Mȥ�"�WDH�eW?�L�0ЌHȬ�3�f�ʎ_���~�y����Sa��*���L���,���R)��s��k@H#�^_?�Z;����\r)�:�Zp���Sg����8���Sغu�<Q|�AL�6���fD���+?X�����W��c�y��6a��*WkOm،��Y��.\r�����KQUQ)�h�H��q��s0z�8���؏��}	���-�߈��u32���\��^U	���ނ��{��xi�*|��6nBgW�~��q:;�XU���U\}��ړ~��+x��[/�7��񃿯����.����V���s挺��k1atJ'H���-�����hiu5ʫø��+p�������p�[h�DI�Z���O?]x6F7V����O�1��n��^��>�]�ўV�ہM{ۑ����B"�EO7mʍ��8l,�E(,Bq���H�!/�(}m����؞�qx�f���+�=ۛy%��D�je�MP�ȁ�
?N�}2�9{G֠��(֮Z��.��ڬ30��^����,-7Z:���6K���ڜܘ�i�?AxV��8��P��ߧV:c9����ǅ��ᔓO���p��:%�!�R��Qm�\
�2�t9�z�a������(.����:	���h�	�A9!Y��k���]��~p�T>V��yn0��@�}��l=o�$�7尡VŖPu
l]��OY��7��;��[	A��<[|Y#�)�/{�7�&6����;��s��{#4�G�$�#[�捖�S�L-���Ҩ`Z�F	��7Ҽ�a���j%'�`	C�rI�A���lC<L���ʀD�T%��M%VU�\vmR �s1�t��Tj'a�SpCf�$7RS6mb�i�eAC�b��hV�p �z�|�ÄD���t���$�Oȃ�D���cd��� ����v��x��N��4|����'�v
�fu���xB��2��"dƳBj@&W1jR�8]Z��AH�]�
���g�#��H�r>����e�;=3�[�cs�q�W�=ޕ�B��dW%1�"���x�����؟�@���9p�q#e0#l��%��Z�ɔ�1�U��Jؐ8N�
'HSrZ��K��Y0^�}=^���-�#��T�i�F�����P�0�,uJ�]��3�����T����s���I���[҄�r�c`:v`�HȜ�( ��H�OPVQ���"���	��5��p6-����]�-�Ǚ���o��y�r%I�M'��s�ǍT#��R�a"7�繝��p���g�C�Qc�$x�e��@T�o�����<�d_�~�b�#�g��5��\�)�`|r(���Zōl�\�A�[����e@t*HY"�&���$̲��Ɠ ��V��*�����߂������sϾ�����E8v��n���#\Z&!����_�KF.K2���t��&�����ea�Ո����&NИdg�����]��k?�r:9[6���J���bu��{��!l`#욒+AO�tR�Bp��a�������'M���T��~�m���B9�$r<9W�l1,v�X�`�j�F8`�U���+���/v����XVh�ljH*V��N�׾~�y��(�%���ko��g^\�#�]p����66�=eŜd�]۷����"�������lZ��@q@�%)���d���p������tT� �$�'����Q��~�r��y�ǃ��rA���%��X��'̞1K�)&Rq�m��O��Mx���úui����٧�?�1F����Wb�ʵ�b���~̙s:�>k���z�PWF^U����I�Y����/��矍�.�X�����0��{������Nbْ�r�w���|���X��*,Z�G;:p�M7�[wކ��$^\�Vmځ�:�14�?%�	uv���>@��� �7O������%2�-�7�����ǟX����Rq�P(�ޯ^�b�ǿ��ƫn��"��ك [����U�b���Q;j܁ ����r��t.{���e���/!��ǌi�p�50���dT���^�n�R��:�:X�ҵ_�-p��7\�h4-<&'�H-�b�� ��TJ!&���~����(��c��vx;z[�r1A�E�G�ȶ�P�p���Kr��'�k�ĕ.���碐O`Ųw�y�:D���6e
�*��g���bi�rq�2��;w�@wgH�>��99rj�qwL$Y�ۃ���c�޽���!�֍��/��s�'i,�@<E�Ј��$a��l���4�9/\�J|���.ބ%+��f��;��#��"�l�$,� ���Zސ_�:�VPj�����:t��6�p��ѵ��v�_�!L權����ϤK/K!��`N�\�#a�v�\�}Ʌp�=h�iG"K��S8S��+�I�"����p�تX�At���0XWࡊ#����ɖ|�00b���B\��KN���xצ�=@�UwvZ�A�� �L�o$F-�H�v�Df,V`W%k���3a�p�i�&�� 2'��5��Ov�e�	�)&#3&���G�d����|�����	T�.�@�ץ붓A��K
�����'�-�$)��2βǃw4�z��9���l�G�Й`�[�[����a3�B���_'�v���A=;�L�>��Y1�a>JY=�|�ENg�?0�#����]���Y�!���4�W�`��Zɑu}
���"m>��Ngg��W��� J��^�
�P5����,*�e�f��N�:M�s4!�!��ɨ���l���*I���[�)����/U�������YU�5&�ڙ�yRb9���rӵ0P-�e�G���5����dë ���Q�,_D�ܴ`t������j��d���\�)8�P��&,�;�����	�gJ�	IV�",&����mu0�{?m�Td�>����:s�)";Z��G�LA������ʿ(Z�w�8�'�l���<+Q0]�deX���g�<��*!�)���(�._���Di��e��R�!)s������_,H2���K����+p��b��FdS�3��/�g?�w��F�BUu=Ǝ��ѣ?ٶu��e�>s�R��.�$��~P=���Ғƍ�SO��g����:��ءommǚ�?��M[��b�+3w4�ƳsVP܁/&���u��@ǿ��UJ'1y���G1k�LU���I6&�xێ/M���ֹ��(u��}ɝSJӖ�KW��/�Ͼ؆�(�C)%9	��0��)x�{p�ٳ������;�W��g_zM�:��^� q�k@e�8�������!�!G!�X���|r��2�$���Z��1ޤ��_b���	c�y�,p
fSU����!x��.���{�����Ҷ�V��Ӧ��t��g�_~�̘rRTet� I��.����;����	,}�}A�2�N9}6~����x}�2��b���`�|�#Rt#��O��\��S&a0��ҕ���3ω�v��W���/FYe6o;��_x�>X���|���ŗ�G�@G[+�9(�����!z�{+�x�2t���[oƽ7݈x"������ԓ@�`B|�x�R9�{{0��_�������e�^����Gc��/ϝ{��W���(!x�Ppny�/׾�h飳��������z�;�n�Z�߰{��g ����*u���.Ăy������K���O�3�V6hp��z҄�j͜<i�HKNBC2l�S�# �R����?ޏ�[!㮄�_%�5jlJn���.��'A�6�#���绰m�G9�(�d��v���Ļ����Q��U��>~��3�1�ÙÅ���7,�)3&���0�ڇM?�`o/&������͛������knV@2}�L\��*444�[�@�
l8r��i�D_�]{vKW��s���-<:��nC��{Œv#n]q։��I��|�.<��CtF#�j��t�ÏAU�(���8�)$A�o�Q�a���ٽ�--@gK�"���߀��l�+\���J�2���L%;oȡ�� w#�ץБN� θ�<̻�8�>4��1M�m��0�ª̶���Ą�N�3�)���V:�ɉZ	A&o��(Y�4�G�9�b#�'�B�	 $	?�ު����H&d��`ᘭ���Y�[�^�&)0R}�9��|1����K%��*����{�x��_�'�����f'!�
N�d{��U��`�-�ϗ@V�U>�"I�$T��>�w� ��^���e�,�K���X�u
�qq�c�$�<X���0ؐ!�,lWD�.	�!湛���!W�	���I��2�e���wB��� SI�U9f�Ī�%�E�Έ��id������'�3�P0�	�`�aTvg�Eb-�Z�T֭`�F9�V�q&6���0+��us����*7j��K"Ad�q)K��������@���)(�:lLtoe^��7<o�����uK��m%h�9X�9!�g��Ύ�p�k��1�{�J/ԏ�h�ˀ��<3�������7HS�ά��9iا�a�3�%�e�=�8��x�����M�p�x��!�؈I�ԍcBo�qΐ;�s�����N\��n'9&94	q�Q6�D<,��4WTR��3���|��q^�M2`慕�Y�>?��X&c;L##i9�G,C�&��4FV�!�Պ���E��K�>;�<&��>��L�,��[@9R�D
i�{��W���܊��G)qa�C��|C�	DJ+��8��v:�L��CG��sۗJx/�eOg��Z).��NsT��¸1�0u��;�LL?�ͭ2Iܼu֬Y����LJp+���s����}U��4�x�}�I+�n=7�"a��:���������^z)J譄�DU�}@�ev�8cq�&�k�s|ѫ��gJ���0r2Y��؇�"��D4�4y&�Q��Y�o?���?S�b�O��o��^X��d{IӠ��l
�rea��{vlCs�a�3�&�Q_[����2v�1Y}c=�����pW���/<w;9�c�ߟ(�¢D]�%�;L�\י����AΧ[�!��}{����&�|���� c��A��z�T�,-�����g�[�Qq��g�z~�دQYW�W��7�Z��M=��R����>w�X/�M����
.��D�9����x�O(����;q��#
b�������JF?�Yg�����Ξ���QP��4T���^,^��Z�݃Q�u���-׉���K����q�s�l��T����&���?p7�/8C�4�%,{M�����y�����_���C��Pp-}��^}k�ϋ�K���R��C���V��>|����Z����#R�5W����3s��O~o��&J�G������?g�~
ʋ�H�p�p��y�(r��I� ��i3>�l?z�~�]%2����b�3��Y�u�ȼ(��XЇ�{�z� �C=h(���@���hۿ�v��#��IS-<� ʫ�QY]��d�=-�2u���J\0o��BȤ�ر}+�|�R��$��7F$,�����ۋ�h=��b�_|�8��yzB"�y�>_<g¤����@�5�}ͭ-8��&���)S$�G�K.dL|X����G��xb97�I��WW`���(G�b�D����.=h~���~�A7�˃�o�����AwS����[�D4\�ʍ\��M�s|g5����j�+
4��ˮ �;i�S8\�9��s/�G�G;[�!0Ҕ�?3%���w-c'�2l�;VdH7��Y�$Z����GU��@�	O.�\:i*w��h
�m�3�٪V�ؘ���
���b �[�S\V����O�Y�'��$;'�O �m����W^��dd8� �$�m%kZ���@Ql��`��Z��P�Z��dL�ѷ�"�ֿ�	3��snv�۪�RԒI5����u�J�,��O#=UǏs(�����@�Qѝ�=X��%3ʾ��x�FɈ�s\1ˆ)�����Cb`��rL2P��dp��ň	`JQ��~��$ikY�2;A�q���j�)W�b��*�q/[����o�Dy�:K㜉`4�/x��	0�ټ:_|�fC���V����չ��@�(�ء�� ������r��b��z�jl��L��/��(Q�������q��kw�l�Lb,�LV�� \�Ҫ����{�Z����tP&wv7�x�݆&�5��cun�����9q��SR�cဢ�s�����Es.�5�/���c����@�$�C�a��'�l�	�����4H�L+��)��Sǜc�w�}]p�R][�TV����v%7E��j7�z��� >k�Ӆ|&��H0	:8�rÕ����1��V���y����2.,-�Ĕ)�p��9��I���,RkL2���R��0��$���K��(��`d}��rN=e&�i��ի�*L/?SP;¸D�6�JRF o}�C��oH��+�궁���Ĺ�N&�����Ž�~ӦMG6S��e���W_ő�G)��=�b�y���!��K#U�ǌ�Ƒ��>ڰyg�M�n�t'�C���igL�7�s�%�U��>�sU�4�3ӣI�	�"
HH"��%�1������8���Y���`���L0IB	( ��2J�0�<��9V����{W���|��^KK�QwW���o��}��������VVQ��9ɭ��>����15��*e��c�voO?�=�\Q����2%���ߛ�ԜڷÇ_A�V�����d(��Ţڙ��ׇ�C&�/��^{����&V���N@L
�A!��x��{�Y!���7nx�u��2v��r �/U�}���Ï>	���i���\���������wމo�r;���~�y(/��Z���2�O����+����܎��/���!x���!��O{߸�6���`meU���+/�{���w���DK˫������;�م4>�[�'>t#j��v���݇�s�u�U�`��f���w��g>�	\z�k�R��k߾w�}o�P�?���.����Ͽ|�T0    IDAT����O�!���;���G������V�?��ɮK33Z�,�C�8�tu�B~d�|��p��<����ރ��4�	�Shwlx o��2\q�E�E�d�L��n�g��t���E���A,��hz�h��5%�-*N%l_h��g��a-��r1+���R����1w�9 ���c#�=��!��C�� B�(�V0>1�7\�:\~��8crL6��f�=�N�:�ՕeE���Jf�L���Ռx�t,x�ފ����aju��i�ڔ�i-鞴�1A #�}��C���$�#_�}��P������t�>|w����-���#>8.G��h���|�AU!/�� �1
����
t|(-dqꥃh.NM����t�ڵXkSD��i
E3T1�2�:�t��&`'��'e�t*��/�DNC���֖Q���L���I�� 0@Ͽ���H��`q�s�o6<��ak��1��[$7��>�kjUG�N�(�&:bt��:mjrT1���R�F`CA Q�-|�,X�4�FB� ���>ǭ��6<�!p߳�sꀷ6��~�kd����v���4DX��(���<��1��l(�~��g��Љ��c�bBZ��n
j(0暻߳^��z�7 �!�"݆�f8��Vd�bvTV���R%��*`�Es膺�,6A���h;�ZSn#���3�Ü�0fQ(HL� c*���N<Lrm�L.L�{h�LJ��1)E�B��V@��4��*����l�s|fy�ҝ��6-��m3���b�JA��{����+�MC��u���e'����d%t�p'U�il]�_��m,��	��!pC�u��Wwo |�B���W���Y�,����V��E��,�Pǲ��HJ����a�0q��Y0ʹ�.��E��CpM�i|��6D}���2����oK��dsP,�LD�.�m]�e^�k��n�FX��n�=ϫ㲍���u����3j�Jbx��(�u\��Jp]q V/�طu�O�/����UD�0Բ׏�ỲǤ9s�ƽ����J�$�!|���>p��*ܬ���_��5|��_�����I��{6�Ln��6���S����T�a1�p(%53W�z&�=�z_�X�\q9vLnE�g��EfI3�*�g�����K�J�z
��X;wO���s�R�١��+��m�u�^�w��@'���O��_F�TB<�Y����L�ߋ���Ӏ��g``���<p���?y�z�;�2�<.��|��g睵"Z��&����N�z�qrfI.C�P�ZK�������s�٧��8�p�k��pЋ��Q� �]�2�0I�&g�����k�K�.Rij����w�ܭ���?u�l�H*��$�߿?��~��������k�p�t,��&
�y��x�l���?������D�������x��s���������gC��ՀV�ٳ����p�����[�����5�|���uo��H?�����w�P��&�����nx�����n���~'ݶX�1��ޟ�����}��'>�i\�v���w��K'f�"2�k�c�Xۋb:��/�����q��c!Sė�z+�}���Jz���.��O��������=|8��y�?����	F{����`��F�OnF_��ǁ� �cd�_p�>/y�a���K�����	�����׽o{�5��A�L8�)V��8|� �M��'����c�BY9�O$��%5�.a�Sze�H�5W�!�c|d��*fOB�S����©�(M�S�jZe$B���6�#��"�ka۶1\x�Y8�Ha��14U�i�>r���߇�Qd2e�޻�x�;p��stඨ��Q�|׀?�J�����Y<@|Y���jF��;&e�ǃ%�c�^m�ӎ�\�u�cx��X��P�&��7�D��<).��%�ۢ�O h��@�EB��A�������C�Ν��Y�ذ���Nn��6N�ޚI/��=�m1a��)*�tJ�{S��Ej"I,dVQiVe��Ô>�r[��4+ޥ�k��a^�?*�jdh?֎���e����)�J�}-V䤲��/�`�@r�m�����q��gu� {s��}�������4*�'��l�u�'�'��N��Y��7_0� ;u����D������Ы?YN��������\�|^��\��u!j�sŻ@w�XZ������66@�]7D�Xskp�8�x�6@�D�g���4�/����o�#o�R00>�%�m�ᶺ��\&���*�
BkE��_z�9I�����L�bd ���d)c!���z�����4gY5��	y�����g�i��yQ
I�cG*Č	����l]#��2��HK�ͭצ�6e����'�lB���k@��p����	0�8�v�x�b6![zl2��Y�\�ހY��EO>\�Ca1�3��u+n]u��͈\��z�u���1i���*чl�s>�P���Hw4T<�����uǤ�M��}����|+σ�˼��84�.�a���8��Mۆ�5�Q�2k��|��z�b��~FRQ�f%*�峈���a��Fq��C�6�t`#��QA>��T2��|����{�0�
m����O
/���ر�L�ر���� �����e:�6_����B
G
)����,�RD�#�i6�\Kl���ׇ������3��Y�j�����hMm���
YKBKhM�{35u�|F�T:%Q�� �h�����
�T_J����aQ�(��T}ppmo�]�܃�Ba-�()
��,.yݹ��?�,�ٳ�=��6����㶻���rQ���T�bzz�H\.C�x�<��Ve���q��UGuX��}��pl=���0~�k��}�R@�*iXb���Ie��Ф�"
�٤-��
!��y˖͸��{t�>���㒋.D<F�\F"�� [�5e�/���ȳW�W�ޑu�_�����^�B1�'�z
�P{��Ț��Lz��&�\y�e�u�>��fq�w�{�}_�C������>�쉗����˘_��^v�m�r�99����o��F���hc5�QB�?{S���w������������㕩9�8 ��]�����Û��fl�9��l_��]��?/�.����7��O����=�ݣ���?!x��ӽ��;�����?����b�~��m�ţx݅���wD��#/��󷨖JZy�X�����AŒ�6�)N�/:w?�|�58c�fM"��&��B0�?�Z	���)<v`��(���fn�&n�p�t�yR
|��N�f�f�C��:>*q��F���h����i��!�e�B�Wm�(���(z�\ULn��=�14؃�?G�Z�@J\�c��ŗ�ñ�1=u
�l������9$5᳼W�P�P��P���,pR�M��h�P����S8����%��{���o��ڹs��%���g���|;��􏟅B;�N0�6'9�6�3�i'�|���|55D�C,�*��W�p�$�s'�&7}��FRv�]����i
���m��{e=�¢L�k4zU������W��^s%=q#*��z�>z������ɈS��\�g�5�:N��с�\��qf�EA�?:�4n��b&���ą���U���,[�����(w�?Q���y�2��\��ޛ���u�Y�
d��\s�bd�ּ����n�\w��U�,bAC4r�m!�ɰ���"�z�������[��|v���FUb���Z��~��Y�[q��C�����Q>֛�.EҺ���v�Š���Ϫ.�����Sa7-������J"�3��;�!E�|}+,4�cu]�J6���kݮ&;�2�
�6��r��&C4�p���R^��!xS,�"��=�O.JJ��@�h�Yz��J��O:
�B��SnuΪ�W"�S�;�AW=�ƈ����s+�y�[TvcA뮗�k�:r��M�M!l�u\ӹ�9�^맭�a��7���w�4�*ǵ�A�)�r�jNC��k�=�K�8�#S�.4%� �'6�����knE�v�r���lZ��5>f/s���{0����p��ה�/��FP��QZ����4	���}X>}\A��E��E�T���X�2��W,���Т�r� �F)����>���}7]�͛D��s���}_�ڷ�$(��������&�.8�8zz{O�Pm6�+��{ﴥ��O�y�vP�eՐqP�g4�wt��{�037���R�	�iiF�eSvύEe���s"CM��J/QgA�|��$���:�{�z��4�H���	��)�Tg������z�ʱSx��d}�YZB�ZVH\�^�ŗ��?���b���4�BX]]�wo�7�q'�Wr�S�@�Z���S�9�h���{�����"2�j�:ф"�V��B��:������	ˍ���*-N�}�?9�O"���*�=A��j��� <�<��8�7��شiX��U��}.���wʹ1�/c%��/~��
_kyȕX����މ����`d4���U�/.��&���HH_2���Ѣ�e�́���?���y^L��|�{p�uoC4�Ľ�>���_��|^Oo�lQo�\q��g;&{Mh�j?�1�w�8q|
�{�M��܄�x��Cx��#X�N)�m��Zj�.���vn�a���Ï�~<�Hin��׿��?�������>����!��������O�y��O�l��5g��AO4��y5��bz���o_@v����^�� ,�+�2r������d�K<C_�gl�*��Bk�|C�PA��	̧�x��x��
r��/ʥ�
3:�p � )D��چ�UJ�ZC��I��Ϥ1}���E�=U�y���P�-��2��*�0xz}O0�R�V,�P����>��]{�U��ګ16Sg���n#�_��O?��o����7�x��GWo�)�kMDC~��P�mX�ZXn�bK0�sϿ����Q-�Ъ6������4W��w���K.��{Q* _��;���%�Fv"20�J'�"���<"�|PPʩZ�����H* O��B�Sm�!��d�|�˳�4�d���3�Ąd��ɔ��1N?`��W�a��<�EoaA����Z���I����������9�u���M¸<��8����eU�`"�6��In�W)�s�U&vC}L�RZ����2��F���F��nD�Jb%�m��F���,2���[<��y�4�4y�<�c�:=I��|�F�h���ˋi2�tԐ�L��r�v�f���9�FBԏn7��m��"�rI]����&�N��S���&���fZr�qT�Td�P�~gժ�M���e�?�~�Ud�!0�װ8פ�;�!;E�M�l.-w���Y�v�o��˙�7��+>X�7uDER�I�愐u�z���]�5�H�6�7�q�p�K�u\�H�]�Hb��i|�ke]�4��-![������� F��DZ�P8�
y6��p��s2����� 6 ̬q�
p0` kg���E%��rt^��w��n�`�{�Ap?ǽNZ5u����_����-2���g�k�G-���P"��t�(��̾blo�3V��Y��o� [�06�������6\hX�`wH���zm�����;:�k���t{����5 �Y��)}���ϳ!0�;�m5>a�C^��N��Cem>".,��,�7�C�(�KjՂ�A{��O�&n�����/��?�_���ar�C(W]��⠾��e!����'��NQ3ғx��*:�:"L������F
F�����.8_�Z<������XI�ɉ�띃&5��y}H����3j;f����D�kA�|.�s@�Ki�����׊߇D*��Q���ӊc�@Q��e�波fQ���(e��4p�E���ػ�}ޘ?���,n��v|�������꬚�Yz�062�}�iL�:�F�"�����X�J�J�����^GKS�7:@qߡ�
Q6o�y��b�� Ɗ��1���k����1U����G=��Z�4O�w��{oz���<���<}�y<��a�I������Op͵�G_?�.���F����{<�6*�2>��� |�1!}�)���?��{+���a|�[��J��f'��7��bc�Q���w�C��$�����?���{/�+�x����>�A�1ڧ�U�mH�]k���ͬbhp���>���s��S���������ţO��]�������^��i�{����}�{y�S/~�g�d4�A����ҋv�w\�M����)|��^9p��z��Mo��PB�:�+�U��a�%(�8}|�J�^����0*0��Xb=X̚��c��7z�����x�I��hW�Y��p��h2E���J>�|@����shU��k�-����Eu�@�N�y;(��G��O�>���Ɠ�Gp��a�]���t �<<:�P�w�Źe	��d�O�]��j�H ��<��P%�ڤ0%-T`ye�A!����<� �W������EL�TB�E�����mx��Ch��݁���&���r7ufX6���[B:!
��#��js��z�4:�Ex�LϬ�!`:��h����yaaUC"�lt.�I�^;R�R��h����o�������:89Z����:z��\y����Mw��+
�c��V���Yί��7p�:��h ��'=��~��G�)	r�qV���Q
h�j~v�����'g�aj*�.��)�{�uY/T�f�����rAFn�t*��l mC���U�ʐ�T#��\��/�_���ES���5@,�MQ΂�_]��� ����J�r�����t���A,������4��H��j��q��˭O�I] ���LS;`P!��� �i�,I[Ʒ��!򾽖�a0z��BD:���0��t`�fZk�,�DTp0��כ��Y�r,�b"(�(�b�M���\?\��$�5i8::���>5A�N�&$>t�i��TQLlhtj�"äYg���=C��Zfm<����W����)}������j�,��BN�:U���V�4D�
�m����C��d�
;�߈���f�͎C�������#u�\zVt�4`�=�f�Ar�(���}[�k�u���Ʈ_!�a5��n&�K���/ol��>�(]�yx����j���L��`_�|>�lQ�`�5$��А��h	�F��*�<��(�R����̰@�F��F�TQ�ٮ��F=��ާ~7���1>ү�f�ߐ�Pn1m�؁�Va�c�`7͐��zx�O��#X���&*x�҉�\&ԩdZ5���1�B����|v��-[ә�y�ZD�:�H �T١�耆�G���+v���b�I�WS��}�ӑ8�5�&��2�@?�F=@,��k uA�3asʡA��G0чP���W����i�5�9朻�����ۃ@��<X^���������:>��DRMN.�E$�UW��#�x��p��!�+Q`d�_|Z��у��#���g�J�6��!�A�K�]Q�;^c�+�I�JH#S3ժ��J����	�&�s��n!�5_9_G4�<���Iϕ��G�h! ��B� T*��ګ���W��R���� �k�af,��ԓ<�����Ï����h+H೟��}�;���⎟<�\�O0�H�G{&��jagl���S��׀/��o�+~���Q)0:2��~�ݸ�u�a�?
�,�"�����ͤ�����K���'�E6����Jem����᭿�����_����_�2�����������Ƃ��N�#�2F��\p�&��Cx���{Ŏ������#�>��BsP#=F&����O�	i �7�3$�o��|L7m�#?o(�\͇�:�G_��Z9�b+�[-�������5�&��_4[�����1K�9�����9dW�P�̢�_C=����QTWf�JѴr�@1I��?(nn,҂br%_��;�k���#� �'Fq�Gk�    IDATÂ�<�����DLLL`߾=*���qॗ1���b��VֲBX��
er=x�A����lx��ʞ������m�Ė�{���P����A���	S��A���LQ
�{��Jn�@�'�0���%�8r3�@n	�F�4^n���s�fSpol�ͣk�ĂN���:m��<@jhH��W]�FЃ�K���+U��vиKFeC�����Fʅ��-�_(�)�D�V���t�&��"���p$(��]nR�
�@���*'`L'eA�l�\���Dt�Ri�V(��B���x@�~dy]j�}��d�фL�b��~����n�)��7S��k�m�Ҧ�Y�c�kp6Ѵ�c�J1�q���QR�,��D�B<��i	���6�݅.M�6ۖɼ+^��JW�V��i�/���`4�;Hf=p�٩�j����;�E�i�u��˦���fUM��N�b((|�*����;[G�(+��EE���k�_<����L"�4jR�x+|�7�k��g��ŨiN�]Z������]a��]����r!�V+ISD=Lќ,E~87]6>|�������+�?�~شf52v����bUG�q���u�Nos��]Q�͵pz~f�����b�6J��H�[�눁��p(�-�F�5,��ߎ���T�
)sRss=J`֊A��IC���y�v/�M���X���3��b�hKa�b�*�?���?�>�iZ�G��V����>g�L�Gm`& Q�]
x��F�^��E��t���j��;��VUUY?�!����U!��w����R_Լ�zHѲ�Z�&m�gUЪ��{��O~7���<1"�r��G~_��o���i�t��)�@h"�J��(?dԬ%��%D�45��&�|_��) e�z�����g��3/��
3|��'�	<���`1	F�3�����ب�z3ף�`<j��:BX6���.V�Ѿ���5K��̸�� � ��U��B	�R���� �YFqaθ����}x�U����w��D�^������wo�M.CWy�k��C�\E�'�+_9FF���O��WЬUT�0�Iz�:���+Y��Z��i��7o�~�5��o]�I46a���ڭ[��Z��JSZ��^3+E�B����~x��jU�NKUm]�r�Z#������
�
P��	��K/�5W�۷�B4��z,~E#!�,,��_�/�=��Ss�z��@8����o��R!?y�!<9�v�� �MT�����r�fW^y�y�[��������/E��&���x-�;g?Fb)�ǒ��IY�4td_#�ZË��Y<��A<~�=�4z��Xo��z��~�g���O?���<��������_��^_�w!O�H}�6�l��uo9��;�\�>�<|�0�9�N�P�@! �VK�ey ����5L����g����;��d*b��C���`�?��7���r?}�(�4�	0b�|��oZ��ׄO���@�?��(���]Ά�ը��,��^TXY#����q�LCym(f�d����ޝ0��N����I)�2ݱ$�Ѷ��ؼIH��v�Ã�D"!M	�F�q��N��b5�CG��1^"A��
Ut�1E��b~yU���Ilڼ��aK-�[~�R#(�(4=���Hģ��˨R#a�kv�lhB� r�,��*�����bX�^�̋S(-.��2+�����j�7�&�<@����\%�4n�F�&��P7��.8:�}��2t��/E'�����ͺ4F��.T4���kr��Í7M��&/mӋ�2�"���9���7�욒�Ñ�x�##C��P(���Q,5.M<p����A4���˴,5
�7C2��e�ҘA��V����'�vl�ύ�5�~�#��<reo��d�g&��E���w�w�SǫI3�k��1i�(Y��)�T�u�a����uC�( �OU�f�ɯ�m����6㦙�s1��,��l
.g�h���b1�(=J�����r���J�N����=6��6�>sC�FS��QCc���.�Ѫ�H�k��%S7E�-bI :�b��_��v��m��'����h*�(����X䄔�~�x��3���b�;�~�c}�Ɂ&rf�s_�Lνe��
A����h	g!%��&��An��Զx�)p��_�ø�lG92������FKϫkY�Y�4l�r\q��w2�5
n��m�]�WNVG�YoƝ�)_��V��ܾ��m��XMg��(Xm�gQ����Ѯ�>��Ym�}�.@bm!}�n�k�&��#5�r�2{�9f�����V�>'���1H�	'4��z��&�r����m�GBr�/��Op�4b���Qwd+��\i�&I�{ =��B���w��vLNn�n�hi��?�$��Ew"i�f.��v�|߲��L�_�#d�L�-/�
O![�_�h�L�LZH;�k��+۳y��M��@�Z�����������{ H��x���y�tl���Ů]�q��-z�ڝ�
h�8�dB���鼳ϥ�p�"WP��~�HI�KyRg8H
�� ��aM�i�m4�9$ca���}��{IIެ�:�a-��-�߁o|���_&��Ui�1��K044�G{�|Y�T"�@o��n�r�r�[����H����4{������;��Ќ�0G�Yr{��HR����=��9(*��H�$�z�}�BZoD$�ggt}z�G������sExAt*E��>Lnٌ��!C'�h&�:� ��2f��Ih�(��A��$vm۬=ujv9%��h�8@�ˢ7ʡN��z�l�=g�C$�ZzǏ��Jf�v��}�FԹ��2b� �z�������H*u/��<w���VPny���ͷ��'���W�[���3�6�]�4�7߸��x�����1�/���B2B*�ǖ�8��p7>|��HR~���]�+���i�ԩS��3Ocnn���G<փs�:W\z%zS��8�6n����a�<���q���P� �ބ�$�(`ż�B6�"g�*Dڈ�M1�E�ŦC�UC��A*B~m	�Diu�R�)t�V�vh����4��GSa!
mȵ� KS9�lKh�4&bR@ٓ�G*��M5��d4T
��� ��1���B���o���!���i�Q.���oɞA��[|a��w6F�7+�P����P_ z�2-7gB�L��I�!�D��� ]�(��!����CS(�̡����QF�C����i:���<�;���ʟ3jG���+ca�/�9�I*�Ӄ�/��}���r*ԫ����Ħu��֮QG���"�c1%`j����fo���'���/�A8A1�E�UE<D<���q��1	����9,�dp���V�G���?)�G��Zc�C�<@$���� ���.t�k~z~�B�z�kjltYǺ릹�O�m��f��9�S�r�iSYCS6�~U�4\e>|om�r!N�B�E�4CI�����p�r��|&tG���D�\4u�ڲ�[�eP�4���x�� q!Z�ڤ��S'ֺ�����4=�bh�}J%%�O���$J:����h8��I��
+R|A�y��x �}Gc��C�M4Tp`܃����k��i�7>U�=�\�c�H+"�����F@Ȁְ���3'������H�,�t�l�)5Jzn��I����Z�뿮@'RX�G#1�r�����Mp�hB�0���}�FC�[R��Y/r��x�l6&�¶�ʽ_�4�����UMQEPf��S�e�b�V�� n|M6�>Ni-�,2;�VB����{�"�a%���<���0��`������1M���-��1��#W:e:tfP��Akok'�ZK|ߴ+���4�ؖ���&I�\k�
����!�aG&�ۆ�Y�aC�j��1ٕ4�Z>k\���i�b���� O���3�qꐠB��8�٠�4���ƦgB:"L�Nv���ВZ�&�.PMȔ��5�xZ�Ƶ޳���䱩7��X8~��u�����O6�ȏ̢4\'�#��m�������KNC���*�q�U�"(���CT�����T��E�Ը4%&כ!�b
X�z_o�z	~��V��+�3c _@._�iG�	�,,�?�=�4D&����>I�K��'�)�J��qx2Ʈ[p�%����ئ��q݉VR���˦�Ke��ƺ��X,+l��%]�:�ᠦ�J��Z�?CDC�sh�a�Ո[r����l� iE/���W���-��ͷ}���t�~i��
E�k�p�����g8q�X�Ac�a"�}�:�l!#�h���4E���xM\�+C�!���y(V�{ɺV��.p]+(РTל�GtMLsGףx(,-���f�P���76�P4�ӳ+(�k@�Lv�<��j��U,{�S�ϡ?�j�)�y"\�q��=��6��2����Ec�V�?֣�s�H����^Z�?��Ƞ��XO��%�baL�8�p K��j�X�p0�(3@3���A��F�Vњ���4�i�ҳϾ�͗~����{���i�x�-��������ٷ��6#��:���|������ކ�&R��pr����"ۨ*2�B٥Ez��P�U��oۊ;v!��1���@�@�Q��!8���e:�{S�xC�	�`����]�)�'�z�^�!Q��&`g�1�͡����8y���C�UC��D-����,*S�w8�(i�c1χ3���4՛�S 7RN�+�`.S�;����0`�A8Ef�C��� Z��9R(:^��!N���^�#K"K"I �7�J�p��D�@�RC�����i�| X���ll>���Q��r3y�m��(�!,X^�"}rk'N��[��Y�h�4��5+N]��s<I���2BbM�Xh8<�d�$ܹ)u|�z�p��W�+.C�,e�Pcp��� �4_�Ym5"<$�*���CJ&b�u��d�OF�xQ���Y�ͽZ� I �c`K�*ӟ�8c�VLn�@__BM��J��W�M���Yx=!m��|^vzlz#�$�
L���b�X/&'6iBQ*�������
�VP�(:����v�-��G���f�ˆ!Dn?Q�F�H=�q�%�m��<>3�$xPV�p�fخ#�c&�>�N�z���jG�lG�*m�k����_�X��(r����=ɔ^[HM�%+@o��g�"���Ȝ%���c��܇���:�O��y�T���+(3s��D �3Y�5�(���e&�L�#��m�h ��9Y�sa�>LC@{A��H�
��d����X7�VIlg\�7wM��M��Ն
�F�]�C�|���L�b�A����J�c�Di��'q,�L������'���n<��3Ң�	�)μ>�}�׌�k �T�FS	��D�Zcjz�[d���r�C��?f6'"fѪi��K��)�XT��&zl�����z������7�M��ll�F��>6nS7&lBh
R'�7���2�v����ma��jz�:��c�,� ��,�Ig5�~;�����%r,=�-�y(e# t0H�Ѡք� q��	�I6����R;��iK-P�j(c,��ZV����]H��	>�A���UGd(q.qYT'��@�O�c���2�F�ql��҉#���[Q�d
�9�P=�Wr}�R����ڪ��ˈ%B��} z�H�Q)���R�:G85�vݘ�qHc㧉�"�Ex�Z� ���Q��G�-f@,d�/f�z���CS�k��n��.|���ıc���\ ��#at��>�u��������s��#y�=�Ll���w6�B�8��}�TzN�Zs�В۳�c����a��`E���d�0���E��Brpb>���P8��ͷ܆�o�3+i!�jv�MsY����k�<�aiyA�/���e������b���_,]��Br�q���4ו�㬀��a�!�a�=��jp�:e��������rKՊ����2!r+����}��,���6�Z4;��M�9Ҿ��{>v�Bi��U�b#�5E�3d~F6М!G#��$�&�����T�e�i��~��%@S�j>'[^�*���ZR,3ǡ����5.\���E� ��?;����̳7������_�����yb�n��?8�����&��	�y�u�ba�=L����o�o��L4*U������I�w5�"�λ��F׬u��0wzAm2�2�PQ!�s�^�a���4�|�y�[�h�R��#Z��L�-/+A�#@.��8�}Hp������?���d�h�Oaen�R�zY�Q�����9�fŸt�8�Q�?�ǆ�xȍ�֡�<�PK+k�4qz��Zr��������<�4ĎP�b��w�D�|u+���n�.5���g�w`�Hm��6Iu`�ghQ\�b�+ѹ��}1�͈y����Ʀ�`"�`4�⤚�#7��գG�ɯ��!�$S��[�.��[�lEmC�Z�$���Ɔ@�<��3�	o|��p��"[+cvyQ�,,i=ǃ��&�u�0�F����gsAc�NKLoJ鐡09�5}�l��cG��ϔ��TL������ܳ�(�u��|����Vs�7$a����5�]7��q��E�"^l��p��kjW:^L�/�0������qj"q���d�:9�!�����H�\RZ4��w��?'�,@�h���>t�z��a̯�9���]�A��>)�5NЇF�t=���i
����
N����J�JYt�h �T0�h0�����y#<�:�4k81uJ��,XY��s$z{4����
żx�>o�@�7����|aY�-�7��@h�^1s8�e1�� t�Á�h8<���5M'}�N���E��!��:ņ$��\N��ZUN~)(���o8$������В��͖��{<�yX���B@[�H�ڄ�y�t�!
D�	Q9}[˘f����Q�L��$K�mMC�R�WǤ�j�Ɖt��\.����;=n�C[��X���b��߇MSmi7�����d��VC�t��;�&u�%H�z ��B	�r�j�hk�""�����4+�5T0�.X���)$ח?`t#
x�?MҀCG|�s
L�E�;����+D�;i5j��~y<oD� ݔ��F'To�T �3�io��3k��	��zY[+:7E!V�����P �}�q�ZU�jpy�щ���-�2t�g����.���m .k�8������4�1�r�ʹI�9'Mf��v�<���DB�2�Bz�����*¡�������z���!�a~qN��-[�c!��ߍ���{�uS�ɕ�L��\z���&-�����ֈY��L�\�i_���9�0��"f���+�Tqx͚�F����}ߓ���'<���#3/��C�I�u!�#�w�i>��\�f���wm׽Q�T��Cg��$�7͜���GF�n�$���쮷�h����ǃA��8=I�C��w��V�-Df��G��+��[ο~���ͷa%[4�:!�@.����^�tû�ӓĽ?�����-�%cIY��xMi�\/�9]K�h��f���Z��3�5��!�R@-5Q�M��RsmB�|�"D�y���L݁ix�B����pO�땐?����p-SD���^t��K�꜄l�f��}rc��N[j�a�Ў11�$�fW��I�d�X>"�(Z
�5�<�U��ҾI$�YC��C=�������	M��H.�e�-����L���!x\]����7]�'o��>��C��}O~�?���'�ڤ�b�&}j�:��U���ُ��l����?<���-�[�w�YHF(�1Zӥ�
��ů����T+�z�w?��� �{l���,r������=��ٚ�I%�Z��p`��*Ӎm��D*5��< R�8��<���X�?-�z�d�NbꥧPJ/�Y���q�#2� ��W�d�8���%R��:���-X^]��'4�
�a�Ý �K��4�����<,y�E��;�X�K��Y� ><�g�C$ދZ˃t���xZL�s��b1�		�D�'O�Rz7ڶ�'j�c!5�09o���'i�	�    IDATO�%�8���k�ƴ�8�3�"��D64��7 �!غoy�u���X+�1�� Q1�3r����l�)���@cm*^7'~��z�כ���6�#����է������0}j�HB~̡P�wL`��]��%��o�Z[-��$�m��Qv-���A�|�ٴp��&3�m�/����ą�����J���\���V`����e���ڻ HD������PЃ���n��� �Yn�-T*ᐦF�^o��_���	��زig�ށ�����>5J~�����[J�<|�(�?��m��(�ش�=}j�}q��@�+M�8q�33j�x���a�]�����0�8t�ZM/R�a����f��in�^T����qyR��/�Aς�h�'�?pzɅ�1�/!�-�FEw��[K�B��ü�<���0{K%EO��܎�ӳ�. /@п��ds%�--�J����(�sP�h��Aڢ�	��b�k�y���I9�⵨j�����CM}�O���H<5��j�Q2.O�kJ�Φ��k5Eժ)bCA�&�rh�7M���"ժ�ժeT9�k7���HX�-S�V��[|Th�ĩ��$���'_��]�^��k�ʎ��{"�s|�*ބ�m��i�+��߳�ea��ǻ<g6�����?(|�hTB����	cں\�~�jd�Y]��>�"��I���+����I^g~V5�B0IY5|�ԩ���ɽ
�.�g
E~VҺ�i��cr"�AW��Bf�dT�����+�?I[H]��"�i<\?4��� d�g�T�;�Ɇdn�q,�]N��'�OW�i�m6fbk�o�/��|�}D�ZH��0���>J��f2m?'u=NG�uE�(�wW֖�b�Q�	5�2��6n��mx�E�c���$K1N�Im5�?R�8,���^��dK��i���g�)mR��d�4�̝���������S�ͦ�T�@���Rw�s����㥃��ǵ��>�A@��m&t���p�^���\���䇱w�vD�^���d.8L�趨!F+D�g�&+N�r͈�K�2L���)���A�!��A�I.Ąe@H���jA������X�6��fC�B%�E�� >�ɏcǎ3���݂�����I��	�u��YN�2z�0p�����<�Epv���h��$�����x�g�q�gQ7@"�g� ،/i�-i�G�Ѭ�0=u�؜���#(�<(׉*�iH��I���tfCĸ�yY�9+ӚU�hB�I��k5��C�!�J�������"�)��(x�VA%�
y�=}�?z�8`����=��o��2L*e0"�@�{T��zn����>��?�ȯB������·��ҁ��D��@fC�i��+jVs8w�v���.F�p�]?��?��NO���[�n�y睏�����G��vp��q�r����%'R"Qn42)����O,����G��\>���U��5�P��b�r/��+W H]���[��ћL�B���UTrk��3��En6���,
��Ȯ��*�K��b����R-"�X�����j�6�oA:WD�B���H�4J�4�8�
U���MU��oaph#�[��4P����7��M� ���;�Q��	�A9x��;�ٲX�����d��C�qP��M���W�@ ���
f^<���<�����!��(Cf:�6, ��Fʐ2ℐ���l�ѷy׼�x�ůE�Q���*ʭ�I�dҫ���cS4����.n�"ޖ��F12ԏ���ka/�aP��<��Ȯ�ėd���5�y�(�'F�;Oe��x��� �����
����M�BؑBϱ�l���`
�HH|�h2��q������
�Y^+�!�"�K8���-H"��)m�lX��4֏���(8|���p��]�������Y/��O~HԶ�۷��s���h��r��r-�2
�
��E���+8~�<(��s���ޝ������D�hz�b���f򘛝�����&�L`����ݡQ7�
���N �@����:"��l�Ǿ�;0<D�9<��G����*���-c�ܶY�o�}�`i9�^:���%M���� @nO>�kK��12��9g��c
��7���*6�Q�3L�� S)� �KDυ�����i�1ב�L�:��W�c<\9��"�$pOS�9���-�zzz�"GytD<ja6*jf8	�:�a?�׫��|�݇b�"��j4���RJ�TC@�G��2�ŃrBȽwnn�j�d�&�|&��¦6Fr [��F����a�T:���'M�H��-��P�T�(��؈�Xt�Z(9�7SkY9�*����YB�*��B��z�D�6���l�l�} ��F�^��X�>���&�����N\(��6z�G��T)�̠7���C%��Ȁ����X���8�y��>YHFb)��E�VK�1	��;�~0��d3�ω�챙d*g2�!KU��j��]��{EL�,�#�Z݊���]�s����tǡΉ� Rg�稵6�,�����}G�E4�41�
��0����!J�4��3��XSf�o�bJ�tS~���2<�ʟ��{��ޥ�r6��`���}:�Y@��V�H*���`�H���Yi��&6#�ߧϕ/�0?;'����(S�qV%���)�8�0��tO=�<�i�39�<3b�}h�`�F�$S	�$��ƶ�Mص{�m�d,2�]ON�I]M��
�=!�I����ԩXZ_(7����9H�П�U��
"� ��FԚ60Đ���AQ��Q{��C��wo�=�?�pT5��!`����0������2�v��x��g104�-['Eu��3Y%	�-�i�M$��-��M�6iҮ�{G��k���LC@tJ4_Q�l��+����oֱcs��w�vZk�:N��JCq��Tj��s��R�_�)��k�ͳ��&����a�8�:�>�� �T;GBc���-��y�%�p]��K�A��F�y�j�<�ٌb��D����n���ϲ�נ��Kg�L�V����Õ��k�|�G�}�[?��cso`�0(�̅�iW�M�ć�w���u
��җ��g�{N�������Ǿ3�Ƶ׼Q�����<�pƖ3�!E���6GP�z��K���T�a5��(j_��� �0��8QTHq�ڤ�� �1�|[(����"�����Ԕ*��t�i��v!?���e,��`��14�VL0�8��p�O�1j̍���^� �;�Õ�)��墧��dڧQl���TC:�D�h�;�bǞ��
EP�3�(&x�Dt�IC�0FZS��X��!P@V�pr�h�)�a��oq��JO�X���x� j�-���P23�������f×�iVT��*'.�"6��n=^`h�V5�.� �fMA�VQC�F�
 9��l��r�%�*�x�it ��:��GctT�H4v���<%�}r�I�;L��W��zӧ�����TO?��<�h��+
��B�!�=��h�E?�99��vn�P*B]>/��6҅��#�,���Mڗ��Vd(!<7N+������@_o�������x�sz$%�VV2J��3�b���c���Pss�k�㒋/@_��F;Y��k���i>�Z
ʛ�Y���G����c϶1��f�U��5��e�o��)�10:�3�ڧ���\#�9r�$��2�79����B�EX�U��=۰{�V��$�=}z/�t��Hb����<1�D2�&�gW�cO���'��GOD�SY�j�XG9�������_����
Ł@>W��\�"6�@�XF��Ǒ�S89�d���vچ{���R0ds�P;#���d��5�)�����*��bU=cr3�S��P�1�����Oaa%?��Q"!:��W'�ǰu�V��p)�
�����9<���ͯ"�@ 3�d���V�@����>l���5=3���9diL������t�����v���}ƭ3S�L�e��B�G�/>�uC�k6�=V�s$*hsc����5dҤİJ��҂��.b�7�-[T�բ+騳KK�9
�Iu���#�c~%��E
���"�<�����d��8�l��̊8豈Ec�M����A?Qܒ�x�N�h�k�Ƥ�����=�{q��I4�2ņ��zE�A����	��"�T���,������x�a�S=ƴ����4(:�"uv�k�M���0�B���-c�-��5�X7-
)���t��y=(WK2"�z�N�P���c�#�t�H�ؓ}�mt�Z�R�x.������RfU&iEa��x):ޅ��CZ+�]�WP�D�~�6b}�<���shx|���D��Wã\���E$�QL� L��ty:��*j8��ľ��B�1E�Ͷ\��8�����"r#r�
1޼y���,�Mk@�i|�d��Kjb�mۆA�VuC{4֟��>�i�3��.KȖ�ZF�͢�B\?��e�p���1&cQq�stn��=?�!IU��'�������Ө�f�ם��F��p�����n��z��N�[n����0:4�5���82<V�֔M�""zDX�p0655��6d�j��{�Msh��5���f�Z섞t.'v7�z�k����s�P6�7/.̩����oG��SϾ��'fQk�4�a���N�Y���q�2�5/Ǻ�)�ʚ��k�����e@�:<�P&N���ɉΰv����K��E40�Y�g���8���h�aW���܊@@�N��Vn���������?�����������Ǿ��#;��;w�?�+���ܳ�7ЛD���,��=��� z��������E��G?����V���A�0~�Cƙ;����^��Wa׮3�wיƻ;JI����1C���O�ŏ:���X�%gX��T
B�M��:h[K5�hŕ��)f�]��&��7�1ݼل�G����U�x<uQi����_Y�@2�x ���9L��
VfO��]E��E�����@�\\�?��/erI2I}�_g�vn�w�K�l��R�I�p��(v���;�D�����$��JNt[
C����0�u�o�y*��D���~y%�'?��4�U�z�QX�`��a����k���nt2�J��~���-�i'�dq��/�M|��w��[~�:�y޹X+�1���L��"U>�6H��27qM�h��&ҏx$�T<��TQ?06ڏDԧ@��y(�gW�92��j	�f��y8m�7�X"�Mze-�����,6�M���/��X/2�&�٬�L�ϥ W�f=�(��܆�۷"��O��k�^)_�ca-���,�L�b~)��7�h��4t�fSB7�/K��5I}k`p8���&01ޏ@��%V�(�Z��V�Ea�o�z�$=�䳢�l�y��32�\f1ST#ݠ���F���k95�k�Ul�2�K.8[ƒz�:L�b	�J�b==��w<:8N��� ۷��̽g���]�y��6�Mo�2+��|u��AH BHhF,��a'6��;�_vv�O�΢I�Fȴ��խ6�ږ�Y齻��n���Rkbc?|P�tuUf�{��y���1a}��U*�O���<���(Vx��e��.�>��o�#�E/I$��8�O��MЇ�zq��$b]Q5x|@QN����*�ϯ�0��!��'�v��az��Go,��G���?Op|.�YzJ�$̻Pk�ƽܼ��2��!�xV&��������m�7��5���	�%}N]��maI�<n��	RM��*޼z��օ��E<�^YJy��������� ����u9Af6���*^|�g��_G ��ˠ#땼B�o�z���jC_'b1���VW�y{�[��4<p��N3�!b)�������f�$&�A���I��^ش����X{;zzz��̴�E��1=���k����mayiM����@ �����p���bC�Tb�h���X�_�����(�X���(bvu��Ϋa�Q�{U$�dWV�T̝=3��[.�RP��rB8L(��F�g��4�W�â�}*o(�h��K��t)��QV&N%�B�hݝQ\�tgO�#�,��/���s�:m6js�˸7�Z�N����(�O�J�3�'>��8ԆF�)��6�I�m�VC�ϭP,�x ]iy�89��NŉC�nAOċ���|�G�䲺���d^OS6e�ff	�6V<�`��f�hpQ��4��)�䆉`n��PK���0iKC�|��nܾ ��=���hs�M�\I@eK�2�	* U��80k���Q܂q�L���cT泔E+%&
�lf�0X���=�]��RX_[F6�ԵB�T"q�?���.93�-T3�r�	�ǩ��̻��悹:ST*H0�Y4@��(��Q�#�ΠQ*i[jmTQ`N@>k|D�fP�Xյwt�^��Ck�����������i��g����2ٶH�~vj���T�(o��ʙ�4�4�����p��n��7	8~��$I�,C+a�<�Z��V�l�f�ͦ�"���R�?ӊ��w���|k[q�͗���w�Q�sJO��������Lp�h�V�b"č�������uS�7���s�5I���q�Nz��"Y<��%btI�UE��{O/��(���GW(7ٔ�����s��ĨZ�չ���S������3J��l����J��+�L�������#�����MO��(�!h!�4����B��B�RF�PB:�eeww���?!���ӟ�c�����yV��'�NN#�L)R\_�E9y����X��V�O?�A�T �\3��#�k6N�i4d1.?H�]�7�49�`a�u���
�Xw�n%�EK�&7�3#�0�^��X�Rhr�%�H�lb{}E�����,�D_��C*l��k�iza=�.��'�x�cxQ�]cm�~Db������,����.�%jr6T���)7�{���5{k���eQ^�|c���v)7�J�������\C�Z>�:J�U�MۭN�2ؙYFb~H�57����2)�\�����_͟�o&�(Cz�4j�ǯ�7q��i�g�j������tRAuMZ�:<�8=!����XG#�]{���
賶Z�(�rҔ�(�_\���v?&Ƨ4��2��Z�/h�������p��֗6tp?��#�SJ"���ں&����Fq��	c��z;#P�O9��&.i;�)l�'������#T����~P?�W�.q�,�jeDڜ?1���^P6[��QΕ������E����0vlH��� y}^\�1��k��N��P/8dB6�w�P�o���d�f�|frO�@$�F�d��Xm�� 򭳽�Qjn����lo �օ�!�zԨ�Sx��Uܸ=�j����Ń>BWW�}�c<H%�(f3e\�~_~���n�??��� �N&)W�g��1�����T�.؜>TI�P���P_�������I	|@.SE�����b6o�4[�v��f���~�ʛ����V��x�����7eG&��Z7zw� &w�h���<��*�-�����+Dwg�j^1�ę�o_����ؽ>8�,L*�
�1:ԯi#ϻt2!���U��9��+��W�Ж���j����uH��O4�\����N��討��ܸy��\� N?j\r2���|7�o�{���Ґ^JitD��XP�16�/�?S��B ғ_�Ϣt�n/�:,.�����X��B(�.��ԉ�ho�p@��(W�DKu8<.dJU�mm��9m��ǎ��1t��(�ٕ���5��%��GQ�rBgP��3�o����S'd�.�/=99N�7�s�S��E&��'[���3�2���RX������"m=��RH�Q��c���(����<�F�`���t�Fg�ω���No߼���u5�@e���6���!p�]�~:,�\Kr��D�E_�������J^�ܔ;�� 6ŷ�R^�V�!�v�!8X[RR1�-�U���
'4aeƟ���?�J�J���B6����hN����kV�4�*�$=1M�L�T�<p��K�a�\
��[M�Y���l�TH;��s�,��    IDATŉb��C">����5�H�����K�l�!�E_;��JF�cH�
U�
W�qq[���(R�|-v>��4��x~F�t9=>��mh8H1��=���dճ)`���2�e�h0B���K[4�acT-��D�#�."�Y|Q-�	y�{��;����1�A���_������/�`�PϢH(�����!�T�\[��a�nZx����5����r���<��#L2�J�^\1�jn<Z��P.s~��:���x=����t�?��.>�g�{_��3�r����v�O���ϧ�G������6@�ϩ[Bz׈6�S�⽨�	G>�$CV��f#�� 
J������	^Ǖ����]��,��dP]��F�A�����J���h ��Q)��ޞ��_{�3�����e�/\�eE��Ȇ�/�����?�BW�����󟳝��jZ�6�	ݳ�(�-"�'ll��4�����D6S�����l��?������1q|\F.�Y}�}��� R5+~��
���Tm1�8]C�P�#։�#5��i�S�\uױזB�D�Q�G���S%���P���!��hj�5��\Es�K�I�XD�i���J�T�z��,�/`mq�tN�;MWҞV�:��s�:��}/*��._�ɳ��׏D���,6��J-�����pƄ��� ���C�!�*&M��o�2��y߰
�ƕ��:zn	l\'3d��>�]�
�r�$����YY�va!���'����j�|C�	��͛��fB�~˸�d"�Yl�
"CC��'>�s�?���!�6֐����uܾ�����vc�hBA/z�06؍�('����m�q�|��^��;w���D080���Ǵ��ح�%_�֭X[�c~~;[;�����sg���&���+kX]����^�CS���A�t�F�)�zN�O�b݊�����po~�IN�c������N�e���;��]eǄE��p���f��p�>ҩ#��G�D�8�$����I�Ӆٹ5��ڛ�h����/���k��.����5M�ؔp�BC;K�t*�����pj|	1Y�l��#ܙ]��^��1�:u
�v?�i������
�:&''0���	d�5ܸ{��.�0QD�N�O�%���x�{C8d��nJ��\��;wp���tG111")��Nb����R��3�g�dC�d8%'�:*8y�S�`t���PW��א��sT��F�g���� F���3��E._��ۗo�q	�
D����h�-cjIŭ�ӄ!=`��|��c�=�a��$@�#���d�@��Prce=�;밺���9�*az��c�2�J�vx�H$,�+�A^�	,�3������m$sd�wj�n��:d[ma���K��?І@�`j��������puh�����&gܬ�p�07�%i��U�Y�g���<��%tF�ȧz���zݚ�Ո��e�u�n�f�g���:��W����	���#� �'��*)���l	 �ˡ��&���0wo�N���sgPB ��p����Y�#�'|H0�V8�� ߏ�N�(�=fQJCe H?�=�K&Ӓ��mJZ�v���L	3��1?����}�1]'�ܑ2{&F�1�ۉ0�]ng��0&K���9�*���`f}��Fn �aj7�_���id�K�KC�7�\�9lfZd�w&a*��І��V'���തDĶ���ZE�eG�׎�YI�P,��Ӣ#U�	�,�%i��l~��aqY����|nz��,�V���Mɡ
s�r���|��&l�67�`܌J1�*�!��rU� L�p!���>*%�ahm�8��7������O~�d�{�f�S(�U�Ѡ���|;��&/�$�7L��
�,��8�in!i�Đ�����F����A�X@��*��5X+ ���jY��);(A�ՉP���n#c1�u#ݡ$�gn¸!(gS���o?�g������5�q����/ൟ��3�������� ����K�Tƭ %]y���C�-BY�P�b�k�e4��������b��6��Mn+ݛ��N�m�^ÓO?�������Ƿ��|�+�h;�/���	��!)�?���|����[��&ZT�}H�FN�;�x��>[a�	����$�)�(���N�,�M���!���Mхa����g�$g��#���(�U�QJ���?RJ���O�ٷ��~�_�����i����Ǿ���}�n�>���_[�>���'����� �.�Z��c؊׍D���_~��'5���x���?{�4z�{�R$k�M��D��\�[x�'K���/�!(��p21��Ҕ[+F�U����g������7�%m �����<��9�2�J�l��N�J�."��"CP�7`�U5�aHH%�j5���*�����wy�=�HJ3��� ¡�X�,��t���(���'�8bL��!7�`���UB+fN�>忓����Zaa�rj�x��f�z�b!�ٮ���kY�f�STԹ�ce��iH�����V�27��a���DJ��.k��j��\x-ِl��Z�bB�!O&���Ga!��}}��G?��O=�d1���u�Kd��-M{-�8?#K�LT�2�GC^�t�K*D?��C�f�I����*~��7��ρ��:�c�;jH$T��Խ���[7fD����(\��a��Eo؍�O�8��]x���w�ڔ�&$�<�#�d����#�_XG"]����TN��Vc�f°L@�}K�]a�����U�ְ4����Q@,Ȣ=�É�R(��s+�~��::p��Yt��! �._���u���1�Ƌ|���E[��σ��Mb�� l�M?���=ܝ[����BC��N���X���9$se��a�#�P����}Xw
�ُ�%�������h}�BA�!*H�������M��GG����#���/�:>�lE����#'H	����@�g����06�	���u}�f��~��,����I�p���泄@ȇ�''1qj��:~��elo��t�t}��+ņ�Ԗٔ4�T\q"RFoOF���"� �B��F�*��vP�r `��;����i"U�W��Yp�X/F{� S�������_������hu=��3��;ʁQ(�|vknJ`�.5ݽQI��a��^�$4�o`~a�lEÖZݦ��𜚦�1[,���V�-�����Ŭ�MadЃ\��<"V��(�8��ʐ�Uʉx�qz��~iyC�c�x�H]60�(ݬ&��,�T��e�,�*�����߾�ޮ^��>��6�κ\��������R�*�V����+���Q�wj���Hk6�,���Y�Ͼ���ϩ�? 9�����p��"
5�HM�Zc�x��菅Q��4]��:�t�XhJ-�\�k���b����aW.����*l6?�.n5��{$i)��f)	F�0�^x�D"���)%i���5�/I ��]1y"|�C��xm�Y�ӆ�Q�k��BJI�J�o��Rg�������HS-�(�0>0n��Ӗ'̜{�	�n� I؞&���=>�H�
�4�%P�N�h�!�|�R��S�!�v���t�u���������oG��ͮgu��':��Us���?��
v䦟�4�PJc+�P^S��X�60�2��HM%=���=7�p�����������bwK��M���r����L�Q� ū+W��Θ�ϖͥӤO�������"J����w��~�_�:q�,.��_�"^��+�X[�$=�cbbB-�A�� D6�l荴��>D

@���2��țB�dʩ���ූQ_�'�C�i�г�8���k�F[{�ȇ�{����������7��Ym��
Ez@x>�"���6�Me���3R�Mӿ`Hqv�\y~J���%l�9P�{���[c�'"tU+������ ����`�tB�}&.���%��x��M�u$Շ�-�.� >k,�����O|���|����~i�ZY��?|�/�ݸ��������'�ddƀ��"�NvH��F��`�����y�[��/~Y���|泸x����)�|tx�PP�!��"ժh8m(Y�(:l�ދ+��．�-��%,�9o�P؇t&!|'/`6��H�`��u����`i"��Q����5x�4f�u_UBF+!JCH�vb
oNL�+����e8,L9��"�ͮT=�*qZ�Ց+du�p��%CNs�0+�����@L]T�o''�l��(k�⪐ &/��F�qS_ɡ2�s�+r��������?��<l&�� drm���*�$y}����f
؞]���"J�kz�_J��ʅ���A[y'�Tg�F�!9�h�Hk����}��XO�}x�=�F�Z�����J���CB���6M�NNA؍T�
/��d�m����h�� �r]�m��O��_��̂��S''��#9d+j(��X^�����51B,���;����G�P���v��P������@�z�([�RA�q�=����T�� ����v�2�7\�X9�3f��x��sj�T���I�H"�{�(��ۈ�Z��ccm�~;ޏ��!D�V(��W�I�ԉ	LN�5 S��*z�9RX�s�;�0o|���N<ya
������,�7/���^�I�mp��	L��9sK��ב]�jas{e�~��mlmH�A��R���>\�x��$������z�6���Li�'��9��cCGgT*�4,.���\�yՆ�����>�:���Y�<1$�>~[�9\������G.�l�>�n�(�J��`���&__���hH��e ��&����dnK>� -ª�Doobr���&��a�����į�m��[3(T��J6�Utw�pz���vd
%�W�74�f�*ϯ���9sFM��AK���>�A�<�=�88-����p
�544��j����t7o�be=�
�r�M0��� )��׭��g���XtB��ݎ��!�>هz��"�B^����El���X������α��Cܝ����&��Gp��C�:��{x$���
R�b]}�8���.*nm�q�˰�\?6���6�~�����*��_���>�6���:1K�-�����ɉNd3>���Y�C^D�^��fNL	v᣽�s��{�,x}�����-H��Ś���E\�����3�ù�����)DCV�y]��d8 ��&�q�{�(��� ˦��*�ݘC:]���#��J�Z��W�)*GM)�M>#u�0ܭ�",t���Xk$�FB$�cS�ϳ��nK��h��_�׆��Y
�@,����P��MA��BF35�w��>�?��Q�l4bi0�jD��K��j���)���v��NO@��i����0o�XD>����$h�k����%��v���TJ�`3O����P�
���9m�4�.Ր�a��$���"�X���!?���}����af�!j�+���Ϗ�˃2�{*P	1� �
2�8�U %U �tk�s�͝��=J�!�C#�
�#D#~����>���T�:�ޯ�|�+��~���E4JUX\v�={�]����h��+M�2�'}��:Ww*�M�MM�9���l~�&м,鰦��A��4����^�I0va��0>���~��(�k���=��~�y�m�T�
�ͤL+'���Uo�b�\{������V)���i�4�V�L���P�H�67�8�<;ʵ����!pZ�Y<�T/7ݽ1���X2؎������i�YɎ~>��,J������>�����_���F�����_|����i.qh����@�/����F?K�͵����ߏK�<�@0����÷��H[>�[���$VW֑<Jall]mQ�䥫x�󋇙Ӎ�ło=7��?���~؜�Zx�[�t�?�U�:0�'�\"�/)I,։��Xx��UhX�Ӧ�I�m�.(=^eN\�nbp�?�|�����!�$pJ�鉌������n��j�}x�P3ȤV���ժ�5I�QѮ4��ć� nL�ltlV�,�M*`��E���7�щ�1�P\�	�G9�a�.<J�x�rE�i���E'r�"��
�X��|KW�a�� ��l�q���0l���jF��������T��CpC ���ߋpg'~�Sx���B�e�F|�\N�o:>T�`c��|��AyL���˻� Z��c��`����v�:b] t���č�E�:ur�>�P�!B"Q����X]�UcKiGԃ��v�u�����pa���ʠ����I<z���c��73�	����pq*ICdX^�cii[�t��T��Ԝ�rZ"��[+F��s�a�KՉJ����p�3�J#�F%�X^�������LNM�P�OK�]��l����eI�
�{�~_���@L$��|��W���Pʧ��Cx��8N��"1���T���Gow/�(6v����/�`?�k��I����~LNG{W�TU[N|���p�<NM����h[4��l2���Awo3�	�w�Gp{\��VGoč�'hp�@��K�zk�o�a+�Ն�Y$^�M"���f��=����m��"����gC��2'���eУ�ѕa�|D	��	��^�v����a��R/1|yI
�eVV��qgukH������ ��;��݁J͊�dF�-q��r�12܏�}}}���b}s_zU���k�#}P@�qܬR6
G
G���p��"���H�Pf��͉
i!�a,TL�^o�lf�#`�����\8;!�%�ɣvwv��0�T�@&����i��S#���!w܂t��0y��C~�}$�n�U�����'N���p�2G��r��R���s�$!�R_�v�3�{	�P��
�١^D�m�S�_��d�<%{{�ً#�+bp�}�AT+LǶ`}s;;I��(o"$��`�fL�O�>��W��R��յ���Ur�k�+���만��],�l	����Ї���'�pvz�7�Vȷ�JTe��ys����	���΁K3��Ŏ)jLc�$�fa����S�5�龦���D�V�!���gM�����PC���`6���m%�Q7O�7�9���Yg��ƃ�s"��E¬5�)��1r4e[/�JW����De��B	�۫�)�f��Xb�R�WK
$�~>�q!t��gF0��ĉ�������6ko�LZ�*C#�ڰooo��`0W8Ԧ)��z[�G�x|�3�Kj�eifJ4ͤ�7ZFt^#�B��8��q���a�3�\�6�?����h�S��9�y��e	���#}͡m�ڜ�{H"b�������O��L������~���+�bee�<}u��< �c�k��:�;$)�5�<"���Z�M����5�5���3�tV�����d୛?ϯI��ֶ`Ʒ�±�Q|�����}����|�Y|�k�����Rɸ��ҡ�%``��Ɛ|�&6)��&[ͨ$D-�s�<��
�c�D8w8*"_�!�LL�c�M%�;���ys��GT�<N��v�6U���M�g6B��m�����������_�5���_�����^��'��z��O�ҩq�}nƴ�4o*�s,Vmv�wv m�������ܝ�������޺yG	�;wcC��sm�$ZP�Rw8P��pX���߿����6��a�=�h4�
��ڬR�(¾��}�@��|&�N�s�O�|�؝�S�{��@g{Tk�%)%�0�ީ���|2�j��DU&�r"C�J�alN���3M����H�k����6ӌi:���a/��p��Z2ׅ�1�36#�y4����-��D��Pi�%}~�gq�ˤ�I%u3��n\G;H%�D�``3��/��X�v�6<H���66	nd�X�����e� k9/�7���A��<��]�@3�J,|�����{Џ��z�8��(;,�9<D*�7Rŗ�K#�knd���l0殪����F����������ԗ^~[�+r��z�!��~JU�88�bs���{��M�@i_gcc}G|Hd�X�����2��I��v�x��i���g�oyu7��Ӵ������"?P�Ģmnn��1CY&��d��=6�${��(��6    IDAT��Z��=c(�����g���ˋH�������iP�i��V6�T���crbB׻M�
�ٌ���p�\+����a�8�mg������ݦ����`c7��^�V6���|���$����Y���]M�'G02ԧ�7��Q/��S��"
Ӟ��XトDB2G�r��kWp���� ���S�>5�4�%P*�5���ch���Hg���},.mbaqE����8?���&7$m�'�꛷p{>��ŧ����R@9��.���4&{A=��<Ә&L~='cSq��o�hѽ��%W�#�3�(�|�ʠ��2����G��簳SD����D���@oPj�-N/�9\�ys󋚸3d���ΝB[$�	^�b�V�s�H&�:�-2�k���"����!iG���faqe+�ԵѢC2�fւi�MC��N~9�Jt�KoC���h�����bVXZ[�R����:� 1@ο05y}���lXt���a/~�p4���^x�V��d
yܺ;���+�t�w���NO��G���2�7v�D1>9����|kIm��ߚ�7�y�sە��k���!�wG�Ig������%�r�:y�F��k�X�XZ������e�M����}z/�-=�z�"4�E��m���Y��"��4�q1L�Xwq��mg�5l4@�jJWgfȩ�S�vA��Tx��2^{�&r�Qjhр��ʴT*\�Y�j
�c��?'��D�kN煫
� 1[�'�8����t��,hCP��F�&C^�f3�b�9eU�z3��5/�̵�:l��ՖD�u���)���_xq��������m$CT��`5S�R�R�b5��-h�	�rf,���_��ӓ�$S��ڔ���P�n2�骻�N�!�D�mh�`�@�_���|�y������@X�5��+`��+���pSρ�H���v����J�<4:��g�<�4r?�G�%�v�e�V ���_C�#Y�Z�)��K�����A�\Ѱ�4��$l4���z��<�^y�4l��2N�;����tOB��&������2���Ď�8�{�@<�G|���!�AWW��	6����z�2�KTl�0E���(�ğ���C�>�ׇg�"���o�ƭY�J�d:a�d�S}�[Z���(�*T5��V��.��2�F뚓쎅���<�(���h�����J�-k�:�+e��Lz��gho���䐚�}meU5�6z�(Rzd3rT�c��J����'~���~�/~�������翈��kW�N�?��������C�N�_��GpfbTd N<-V�M+��T�R7ig�T5�,�3�l�����^�)�z�2|?{�1�����
��|(S;N�É������o,����ى�4�c�A�p�׆�X�V���]��y8�^�Ua��m�ڲ!���.<��Qb_4 ���O���)�|1�:��1W�$�n����L�~?�*$l�`mnJ�7�Z�p�T�=><@ü��C>��pju�*P��p�'���Ѱ�k ��Mg��4�h�̈́�*�_0@�پ�\oQ�X�v�*Cs�������>��-V��9���&
[{(o��!hm8M0�!�!��_���/5�T����~k5&��j���;<�'��^L�;�L��x"�l���XM�śSH9��)�4Jē�Gji��T1趢�͇��>Cm���d����Z��r��'.���g%�� �,ck3�����]~/�F�hj@�= 2��֮��G�I���pf�8�>���7�0�����ɓ'��$�0������,�V��į��^�!�3����:�&��u������h�,�x<h:���FW�=݆��U��������Vd�<q��C��@�Dԕ��-�5�H�9e"4�͵M�8�d`?�C�w�7p���%v񺶠+��vL���������=��:q��iD:���Nf��v�6gWP,�1�é���B�V����e?{�0�׃��zcc�җ�Frr��M����Gpb�\���h6�����W$�ů>v=�n]?̄�����E\���Lن�.R`�	ΠV6Ee'���d<a�4��7������㵬�X�2W���v*+]��B�u'C
�x��)�#�2I�����/!��+L���al��Fb�Eð88�p��],.��~��ڂ��n��԰p������;8�?����H?eE�h�R���t�� .	�7DO� ��+X\���;���;�u��ǉ&�$�H�۔=�Q�\��;�T�IhbM�1�(s�S_o ��+��EogGC�*�3����[;;���bd�_�E^�2��-`u�@��Xg7���b�x?�n��17�$:�"'ϟ���)�H��6�����7�!W�!���Ǡ��NL��O�� ��#��H;���ҥ�8�'�9��4n�^�Q�<�$6A�� �u����qD.�H�#U���'�xH�4�͹<.��x᧯cviVg NoH@nR�b��� ��Ch�h�p��{��Nh��I(�=n���"+�Ԡ�5!��+�t}������R]�&��Ak�X���͢�`wy������*��8�3�N�3��K��-9�f�e>_�y����8=C$~G�c��m�FlprLg�An54��+}�\��h��r�v3�u(���f�
~�Wޅ}���h"u��<�M1���qD�"�������8n���tbo�������o=��e�!�y�P�����j���{�7d�6�k�f�BH��kq{%Tͩ�	+B>�ڸ��R*	{S������@4����Ã���4����ZS��-���?�G����� <VkC�֯~��x�籲���=�yGW�NMk��a*�$�pI�"e0+++j�+����狺~�K��c��l�l�]T��Ә����a�����Y,/.a;����5�/=�?�>���+����n���6ů�'iS&*�ZZ�y<�z"`�E�C�b�(�T��E�UC)kW�M:�-����Y�8��0��k�t���~OX��pr G�%7%{񸨔�YГҬ�4�̱��s(��>���>�������i4��_����+'������x��ⅳS�����}��2j��y��d3P�^��bӃ�:)m��k�y����|�mqo[Qd|h0���F���~/��|�Żx����!���2 ��4�`g{��!�>;�ռ�47���h��cM��!A��:��Y�i�L)N� �j�Qb�ȋ	��f5�Q������`2҉��k���F��@!�	������;��o6���dh:T�z���Hē8`�r�`̵���ʼ!3�4�D���:�:ۢ2R96<��#�u{�S�ce5���m���P!O�ON�x ����H�!>��)CĜ����}���7�C���
~s
g:M�0�����͂��	��G?�c��8(d��L>h��'�����A|`jb�Q��v�TJ$ a����%��#��r�|��uM~�.>wv?|FӢ��Cd�5loe�4�� ��۝�ƺ1:C$ꕌhe�@��s���ՍsS�:6L\�8��"{�(	�׏�X���u]%�Y���J�}xT���)�_#��4h�lX�Ħ��5�a���R�c���!�}��v���D"'��XZ<D�(��tN:���~�	��N�kV(�j44)fS�S�@:�����p'Ƈ��E\cM&♕8f�v��9��z�q[��ab8��'�`o�03����6���8�:�ȣ�102(�7�D�޽uG�}�����$=�� 1dus��y]�3�c�x��:L��raq������ǧ�����������M��g�K�qvb����;
d�e�SY�[����&≼���(7j���W�z��gpX��Ճ�'���2�)fX��͗6 ��>6��FQyv��5��m��=��ް
N�g��bn�@?';[g����=8������%�Wn�`ecK?���@g[ �C���0b���o���[wQ�������8��&`���*#�I`aqV��P$���Sh��JJ��r����D�0	�7���9�x�7�&]��e�&�9��o���դ��&��۽�.���
D��[wxt�x|�K�*N��V�-M,.Vvv��=�F�B���=875�����4��𳷮k�~|z�/�E_wX'Q<Q�ݙ��B3��eI>تe��n�Y�܊˴��c�x�Ho�|˫{x��%�492,�vw�Q+eqzj�ΞBIX֪��ܝӄ��^�I+�i�{	���M����֋�գ�6��ͱU�1S��lUX|p���ho���Rg�tⲞÒA�Q�&K�}�󠶿Y��QMͷIG6������(�T̆`{q?{�@�����hZ��rj@9�/��j@zSf|�!���&@�$$xϞ�t
6�ʺ�ܔ�z@o3L1�3"�3Q��"���+J�H�K�<7��%�k�^��� ����p��Y]W�~5v�C�,X�n��nL�v8<���������G/���4�v�R�ai���2�:4�^�w��𬠜��:����n3%>�a���D������B)��@��A�����#���N�{	2D���j (s)����������tm}_�җ��|��r���zǍ��a>����V-�"||\a�-)/
�s�G��=���3�A�M���V�a-C��0����w�P���kv����X�X��G/�>��9~L����o���޺��"���-��7�AÄ�E�����ͦ�l(Gk���~�\+^�u^l��	��T���R������ZbTK O#�^�يЯņ���=�G2nyy��z"͍~�ԩ�qy�!SM�>���>�̿�%j��/���׿��T.w���㣃���b�S	�&	*��*�-/��?��C#hF�wx�L���X?|!/^��x��˚f<r�a��I�Q03��EZ�-���.���Cf|(;j� @�S%G=�����.� �9�+P+hb��)��S>�5Q� �[md�MK�N��4&�Rfo���ݝ�p�h�����j��2T��W1j��ACfeX,�P�2!�'�I:�6�5�hv�t�J�ԇo8�4%��{E�*W�d��kr�̤�r�gK�)i��cՍ�-�[:�C�'��Ӌ��u�P���c����p�p�- ����چ�A۳+��-²φ �Mؔ
ٸFf����	���_h@�;c!񎇁�hl��"������9����O`����	�'�dx%���V���4�4�.

o\N�؄�Z��3��X_a?������.���b��#~L�Źs'�t�t��s��jC@�e�ZD�-�������j�!�`�8����r|d�����������~��L��/��U���&q��]��m��
��� ��8NW�0mM���kwN��$V9=85>�XԫаX��jI,���-���a���f>F1���twu�\�a/�0J��P8���^�4�)�ΗAgl�7�}�����Y�ŭ{�8̖����������G��<Jbyi��q�ol��3�����a�"fss�����^�'O`r���	��q��,._��U���pb|�U]v�|����O^���*��G��#O*M�����:^z�UMg�O��'?�^����L������\�Y��~/ie���T����0�=J(�������y���Ws�k���)�&�� �z��L##��-Ւ�����
j������"��h�|(S���:�����B�l�W�`ckna�]��j�:8�j׆������z����喧_�*��G��~����~��G��?��.��ͫ����Z����@�\�4���;7ഌ���N75��vEd"�9�cp��]�p��P�+u���Z����{:�(#===���[f���M\�1+
e�>�G:�875���`���ǋ/����m���!��#S(cqyK+����&�Pt1bu��;�q�8GRU�;{"�<�ԣx�l��v�K"8�umV�9��qxs��!��c}x��S����L���.���M$7����֍{H-��b(T��ȋwJޒ:<@����U�����f  ��5�,��57���+*Mj�I1n&�d�M���ޓ�Y9� ��V�+�Ѕ\Vt�؜��O��>l���ML����<0��!6�b�棹9oM[�cA"Z�{�;�̚$�5u��z��4'�V�ߐ���W#�ձAa��`CYʤ���48N�{{:����^���Q��駔���$��b�aDmbc�B�E��[0��5������=�+��		�`�N�*�c�:�RI51
�YP�e���5i�!�U�@X��*Q��9Pc.���B���L��m��I���K��,(T���#mj>3��9n'x�����J!�Z��]���������B�S����/�!�XY��E�?��O��W~���I]�;vL�����5r!� Uj��1[g��M"9��X���to�OT-Q�*��,+�P ��a
�n�B�V�G>���G?b��j5���+��/|�n��~����d�[uM6�!����~�X,FY�rɚ	��n��ٔ6eN��T�[A���fC`��qϞ���a9��<0��t:�`{j6E�g��Db�M�z@D�3�#���[x�K2������o�m�X>�����͂r��`V�Y�y\\�X�9k���Z��^���,�I�������.���?)Z����k2d�C�y��i9����[y���:��9�^څB�#���i��RC�Z�����;{����)�l�,�L�� A�=O�c�Կ��3��&������g�K��ЦL�t⭴҆pw��+̃)���x�.�����2���j��2Q�������s��[7}X��IKvXu��Z�p�K(��+���S$�t��=���:�x����4�6��Ȕp���y�7P˒��!(�f��*L\��U����r^��`y,�h�+f�#O�����)|�����ӓ��88ܓ_�����R�u�6%G�5�|?���)&R7;<�H_D�Q~^�W�ͮ��7/���h|��I<t�$��Je��Nk+"?Qk���ر~�X8ȼ�@2��̝�nn����B,F�0�]�JՆ�˃n8�&=1��h
���+�{wQ�ѻ�FQ�t�� U�W/5E�U۵r)���c�8>܃H�����tևG\����3$1��%i���ѝ�-N>����a�Ϧ������G�rX�a�y�8:�U�-�4劚l���+�'��3�8>ܫ��L��ٹ%M�YE�N`d�8����:�V��$1%!���� z�{u�om����W5M966�_y�1�,`�9=n5���������p+�ukk������
����w=��c(T �Q���x������&7|��$�^1I�E.�!iZis!���(��)!m�Yܐ�e�,fͬ����F���K�pa�S���� bm
�;<�a#^��f�{i���*mC,Ѐ�nA ڃD���._���:�?�����Q~U�P;���y��]� �����W����L3��b{sS�������pe3���}\�YG��LBpF��V{�Y���7�(��
K��Lq���@�ư��6ż�b�mDgg7�,��ҶW�y���`og�Ϟé�,�\B
�����El�;w�ΨO��ҹID�.V��_��{j��Ϝ� ![*��������	�p��$.]8�\��H��z��^��@(�}�x��Q��[y\���{��8��`qF���l�r���0��t}�`�2FR�������YX�U�y}���_� \�����LA�7!V�2�,5���Ņ�鐳2f-�&'�Ҥ71�|�r[��<�[���P�%�� E �����S3�0�hr������Hw;�3x�ߑQ�zzt�Sޣ�>��+���-������$�s�h�\���*�˘���dv�!^?�uE��)@ᚤθ��/���v�	�s��8J�!���    IDAT��yCUv*�����ꔃ�14د GN�w��a��q����>�铓pY��Be*h�V��G�S����ug?��WE���ϠPj�!�k�{��$
�|��߫X������bq
e�r����P�"U���Je�# /����L���S)��2K�p+Iw�h_�e��pJ�
%Vf�^����K�+e����S$s��=�s�H�����5�rK��P3�������`����C��I�VR�Ӊ��#���{nml�!f�̕��0�+��YN�yVpk�Me������n��?�,Ǝ��{A��w�<����)����?�{����n���eά>[y�s���Ys�k"��u��6xn�-pP��g>'�nX�~�C�(��!��\��(]w{%ie�Q�4pV��<�ʥ��3�3!�Y ��oXل;d'Y���MŃُ����~����;����7.~�k���J�~���A�=u�~⒘��2����9'�􂫺F���+�&��_��7��?��᳟�oP�����?UCp顇14ЇZ���~�ˉ�Ӂ��2�}q�]��~Ƌ������o�{�k3o �v��!0]8��N'O��7�F�җ����n�Ԭ�l6M�[���-��ea�cv��hyZ�B!#W_bN�.��������dU�)G�D�7�~�dh���'/f�Ѻ��?;oLfo�А��WC�烝��C��I$ꇤ����7ڍG�z{�G��۰��Bie�p(�l��������7,EԸ���I!Y�|�h"�{����R`��J:�8����|��7QCxt ���`���&���#5C�x3�Vʭ��/�<lLC@+����1�߁��0~j�(���Z����E��x�P�>qbv��G����VV�����g�ctl ����F���x�g�O�pfz������hB��M�.$Q���i�v�YL�^\��[oݖ4)����t�ZF���д9�K� )!p�=�E��a�DP.$�)��}}�7n�aq� �E*H�wQ�0��ax�,h��A^��D,�<'4�E�A�����z����D��A�\A�(���x]2��h�� ���148��� r�f���J��l�*��p��$b��(�����B*��{e`x �h;�.��iܿ7��S$�{��$��:��At+�2�;z�����ۧƀ�{�ܸq�o�F������Ft�3h�����^��x��D��p��d
l(�9�"�8��τ�q���!2�����6��y����bN�m�xj%l33�[Vd�<.���81؏��6-��)�5l䕬�MQ(��g|r�~��`�Lů��6�V�Q���ׁPЇp�'�_{$��n
׮�D&��X��}��P�b�??1���-t��q��q�hf�Z݃�lw㸽�.|)�ԡk:�������w���`������G<w�
������N1���$�x}���҂Օ�ܹ��Յ�g:����7noȀ-iAvѠO=zR>J=���Wp��,� ��O�ы����&���Wqx�����E_oD�$�L_���윶���������N�D	w��p��
�"��n��W�0�.�\zǆ;���itE�!"�-`e'���������=�K�����mtt� U�i�g���0U^����h	���@)�]��g��P=(�U��YE	WU�2�����w��zF��<�!�/s�%�u�>�s����'�03��"1"!�� ��(ﮬ�]yW�l���Z�D�6�H �A&�t�L眫�+�������o��sp�&���������$)�4� 6�d��B6	S%�]=m؜��K���T6�"�G�T59��t<3������jh	x�Ha�q�Iu�i�㸮D�'�J�$�Q������؀�W\���{���]QQ��� nq|Ϯ�.�%$b1��.`yyUt�MM>��岉/���M1��hm��?�a|�GGk�4��P.��މ,���e���୷/alr�H
�
�NZ�k��2Pap�����ň\>)���$�2¬j�hdbG�<�
�^7�^?r#�6\���H-�!��c��f�[,Q6�4�ؖ �����[N�mlP�g�$����#��������㏢�g����˯����FX�����q���U�@YY�۬J̆�����\N�'i��~qi�v(9��ó[�ԙ�d��F���k�^�DJ�5�=�k����Z�����x�/ICƠIRn]���[��qR��E�i�A��9��	��	Ko�Y,Ek(q�[�0�|�wQ5�bE�M��d攃���Y���0P����\Xm���Q�Y-���u�wZ��� ���j�&���Zm�W�(�W�~��7���o���S���"*���=s�O����J�=���g?�	�s�9�x���1�tb��$U�ʎ�q�x�g��+��`~�7��т�.^�i���+�E���*��:T�A�l�ݨ���q��2�7`r�̉�pU��o-`u�=d6oAW����`2%g�EK�'�J]��j�&,��5r�Tl�D��s��&!om�Rc+"'�q��l�{C�Ƣ�]њh��V"'Rq��^�P�U45}���e�e�6��`�O���	/��wUE��=I���LE� �C�:�8t�^��T�,�S���)��p3�cHO� LZ{�*U6[j�Ϡ7^��2���{$��!�[���'���^�F-��O�����%���*�Gn�x���9�����6$��.�]�ū�&�rX�!�Z��w�5n*����&f�W��E6���6�9Y�A��e�9,έcfv��:{:0��ͭX�vAj�70}k�Zw9(�`v�Q��(�ne�Gx1�B5�Ո�������7߼$4.��n@��e6rP�غ�E���?��ݏ`��v8�W���z#csX^��P2�h�˴6����Ƀm۶���H�\PR���P,�B���]"�#ݪT("Z���B0��d��-�N㭷����o�������m�\3��BO�@T�/��n�w@�0C�
1`�8����[�r���V��ъ�'�c�`������)�yҒz��4:r�i�Kh6��bzzV�l*��Nǁ}���֢,4�CE���%�si&g,���j��� ->&�Z�-%(�Y$���ɪ03Bk
8���ϥ	��>X�KR�%��d`�UpYp`h }m2 يg�豴��7��o��k��ۅD8��!�^����e���h�hA��&�Z���-alt\ޛ������D�����i��\��iŎ�n�)�
��B"_��jo\���LQ^/a��H�?ٻT1ǽ�,�yMnW�pq���R��r�\e2�Q,�Žj7�#^�����G��������p�LH�"���[+�dU�W2����{N��]�p�X߈��/HƇ�⒂p��n����K��[3�96%t����y�Q�RK����Ņ5�c9)���8s���nq�47W�7q���"8<m�:=R����WX��éc���䁁��|3KK2�س{�������obv5����U:���|�ZV���
���`1pk*���י�����G��B�d�>H�=�-u^5N&ox<����*dG9j�5yf۔2h���pc�����3��bpx�r��L��T!k��-��iѬFUCeV(13?�BA��h��EA8�q�s_6��j����ӎ{N݁�����h��s�?KL�Z��Y���z�nMH
6��ZZE��47���il�/I�Щ���W�v"��}��6#|�#[[���ūo]��K7�A��ѷ��)���R��m��Ao_;������]��-B+��\3!K#�c���MO���<��px�a���Q�ĐY^�YI����nT}#��	+��S�;J�O�˧���T��日! ]꽋�q��y1���Ht���P8���)��7I��h <lP) ��܌\Q�
R��P��(E���G�Y��<�u��O�C���9��U�188�Ǿ�(�臡�Y����O���t�`Q�R�X�����9)v��K�2u���T7�$F�re����7O��
,N+
d 8=09�(Sd,e�^��l\mn?\� ��*�4L(�0����I��sO�J�g�vlHs���\�8�*哴{�C�������w�)�@�g�Y��|��CO����uƽ�����#�CsqvZ��e^$��L�5���b'�Z�}��O��˯���_|��p:=�t�lpg�>��D�#M�l�	e�Sk%���\�jf����z�uLc��y$7'`�F���v�U�E	5d��q��`j#�yv��h]���lL�����qՌL�E	B�E�{MR��N�Q��h�h��N�&�\���X5K��v��*�E��~u��3�l���FJ�h�Ֆ�'5��T�L��8�}w܋�ˏ�D�bM,�t5�k!��Ca~^�E��SD.��5�<��IR+��W�hI�����6N��4S���MY�B�__�m�`+�BdsC��(�2�=�x�t�PL��$]��5eجftw���aC��+������1<%A&N'7>=��mt��a��I��ı���xr�Rxq*�⛼ϙ�YL�O��pុO`h(�J��X,!���)Z�eQ�Ä��ǌ�i@Z��"H�怛7�ƛ�P����D�^ձ�R�>�Ζ�y��q��^�����r1
yē	ܚ���J�"E�tqK�V����ׅ;�>�kka��,a}m�-ݪQO��=(�fCJ����2:[ZD8f�D�h���022,����.��6�����ʾriy�،F��٠u�E$l�	E��j�rQ�.�7 �ĵ�1����=]m��P���Z�z��A7�r��T2�d&-��r���!��R,z�f�O�U���tt��E�\�H"�w��K�]1����H!��������.��v���O�bbf�RM�E��[d �l"��)W�D��F l4��

�8��<z�8�k�ۚQ-�K尕�ar1�щ� ��:0��mp�)d��R����[X\^A2Mo�\���&x=.���%����� �o�AoW�p�C�-q���H�ak+]9'�\}�$E{�P�Z4��P�\C�b�Ѧ�h��2r��MMD��3MYL�FTJ*=��˚��|��L��S,�����Â��>����=��#�$J4.0�V�R$r�1����u+�zo���v'O�Ǒ�%_cvn�޹�P,'��j�@��w �����$��gj�;��꓀���Yܺ9�R�.�v`��9��ߊ��u3&����a�ce�ݭ��qldԗ��Ρ�Ɇ�G`����N(C�vВ��a9�\�Rei&f7`v����H�Y|��{.K( �.�@ǩ,9��x-e�O$�{��ƹ��XMt5��aPmp���g�& ʗ��}e�,:jHe����hs��ԗ1�
�/�C%�����ڔ�I���h�Ҫ1�â�D�,�*֢��S9
:D{G�YA�qRl��3��M�]�+bQ��O��>(�<_+����3E9��Z~O�É�%���{��	��l�1?7���R�-8,&Is��ÿ��;wI4�<�r��������x���$!wm3�V9�*WE|/�F��w�ß��;��	_�����އ.��\E�E��
��y�u�*�:�"��6P��`u�a�bb�O��RY�w<x�2���<C�7�Q��:��E�yqY��n�����#c��q�/(���$�#l��^�|Y����1#%��������!)��V((:��  f�e4� �l��i���Q��Ҏ�� �j6*2�Q=�+�G
E6�m� >�Gq��\�>��~�:��N�\%-W1l��h(8�cv)m�����QxL$��?l��F����yJ�2jْ�--�9P%���\�;��&�f�V��Sh��X�D9��$2���C|X��%��׃���TII��z�! ���M �č�}�����{�<�3/z�'��nkk۾��U���z�?�H(�|�(�~3E6� �ln�tv��'������g~�v�އ'���bO��ko	z��;���rI:�� �͎������n��Dpv
兛��XG���Bx+co#�:�C0�r.3$��m��#�%2��Z��ps���d#��:���A�����
�1�ol��B��=��F�Oԁ�b��������KWS���|*�N��W�|V=Q��W������&��_ţg�"ŃCw��g>�����h�����bM�͙y$��QK'�3r!P����4ʐ�[U���R��iX��K�n�ZZ#&;Sꑯ�оo'���'�هH&�<=��U�$�U�M-[7���u��K{IN�&�t���σ&���mX[+��w����p
-[Z=ص�GlE봬�G�>�M��P7513�R��M�#���������#�����n�B4����� ����*�M��1���G2Q�+���X<'�Y��)�5��2=���9t}8z`'�:���^�A*����V�["8d@K8��$c^3�̈́`k {���U�9I�[[_���M��D��^�|>yƦ��0;3���6q������`������Qq�ٷcz����"�I7���-lFRB�(�B�f�;���������:�2�2V���0��X���ؿg>�Y>/�G1�z3��Jr/'Wtㄪ�=��-�YR"�-\�r�l
>xv��G*�E�"�R7��q��-����x`6�`�W��s��!��҉z'�}6p��DcI���������}"�n��/
�h�ɘ8�(�p���ۇpp{/�����Y�o�16��x��
�i�����!p��LƢ��A�˫bH��@{��A�\��O�qs|\��L�#���LNnu"� #���+�KF��w��c��7��"�)b#����ElDsbyJ���tsͷ��[ziP���#g��5h��+-��fo@�5E�D�*b�@㝻�I�lwq�X�<���Ui�z%�&�+c|r3s!�*��k�GWlf3~���ɵ�yk.� ��[�[F6�^���-ڇ..�"�N��I_o�4�l��*!m��\�"��'1��b&,��K8��{Hf��CB��|���٘F[���y{�m������ξ��~��sZ�SN�^~�]��/��l��D�F�!�D5P@��sR�:&m��/�7�Et*��9<Pϟ�ݯeH�Q�J(V ���5��ze1��F!l�3/��t�":QC��s%���L�\E&{�ƙ��F�\hA�	�Fb1-����������ɰF�9��=�kK���.kں�BQ-$px�v���>�{O�@2U�&��E��*�t+Kz1�_�wo����g177��	3m��DC(����l=�Ǐb�А�#����B����n�������K#�����J�l�IE�K��]G��;�����KOڪPYLz�*E�&�Qm#�Dg����RO�=�k���jH��x��@<Fm}EQx��Sh����YP���2�:T(�=��L�*⛫h����;2������_��?"���yW�^��6Db�/t[�pTҩ��D�+s.J�V�/�#�^
��7X��b��Y�B�)�|	-�� pc&S����edQt�؉��K(Vu�046>�}d�5�a��TR�nh�a���Nh<Ԫ��D-�A+�c��4�0֊T�=�a����݅�ю2�mRF���v�ZD\��!�*���*� ����r]�LF2��r�-�z�	�%=����ԄR; L�'*�R2z��|�?��_��K���3g�>����w��=_��cf�ۀKo��[#�傳p#�A�X/U���@O{'�9"�~�C<��Y���?�,6'^~�Uy�������@�
ü�Ӟ�\�LHCpc:���U�M6�����$��4zNiJ!��yY�b9J�B�.��j|w)`9�Bܠ����p9�ĆM�?8�W�7�F2��U���q�рjU7�6`�ř��Ȩ�C�f����M����hX6?��j"�@'x\3�M<dH�����    IDAT���(��r`y¢�����߁��rz+��I�M���(f
���_YAfq�XHlG�ey�X\�@A����6�	e�:v��&�*Օ��i��*E�އ{?�1��[��e#��hn#3�.ioݠ_��c�#(�=n�]u��u�`����8��Q�[o_��jL6d~�ӄ�:���P.�a��j
�~�G��뢉Y]Z���^t��y�pi׮�k�D�oS;���A�P��k�Ў!m>c&�w�p�
7t%s1�5�Dw�3:�>l�oE��	N�zI��x6�l�
��)	�L�\�bcmM&2�v�ܵ�U�t���r�������I�A�ˠ(�v���#����ڂ;����6|���(�V��Ϧ��ю` (�D<�G4^kǭxN
x6S�\�8���G!�v�V-���aG:U­[�~����C=���@o>F1�.W���u
�Kkr��s������D�9l6A	ο�6�q�{p��1TJy��� +@Կa5���O��
��������6�f�:��˫�����V\�O,�8!b�/@�xkk��v���Y�Ǵ��2�/#�V}������>x�z���sE̯&pyt�\y*�س�;�Z�9a�ې˗0:2���i�����ıg��m��\���XY[����f�4�������BE��Zhu�&�KD�p�ОAX8�O��܊D�����ά�\W�d�w����ܖn�Ty��5�Y ps�W��:��j���͍���MϨ�T
J�Utt������ x��8bш&c������
nM,"�&g�D��߁�w�۩|�'��q����)�l^����س���o�զ�/���]�i�fn�/��{���[��3h�l�=��c{_�jxL��+���+�Q(�k�&�Z�Hx��*���ýw�`w�h������d������a0�
'���Q\�����8.D����h*�$J��n���$�RD��I9��䂨�v>4�W5�Q�4��k�-�����!�r���$U��f��ʟ�TD�C���.C+cø~���X�����B�SC'�i����~�L$����@~��&hs�|�����h�h�?�C����:j�Nߏ����q��6��]7R���_X�m7�=;��W��ܛobeiQ��Z� ���L"&~�;���g�.	qܿk� ����5�x��7���M"���R7�>��D{f��fh��=�F��݆���/�cy ���W2��ב+D,�s��3]�����$^���q�5,2'���9Ąە��sN�����t6t|dXC���Ei:��,tҋn��ك�����݊���C!�B__��+"��3�lzz�d\v������nw���p���dA1?C#�Q�2?$��*<��gcP3��<�E�`�J ���>�9l�8v�nt�auu7�g�M��%���CO_����sb ȥYQ�DMרb^���ڄ�[7���&���g!�K�}�w���<��^A�4G*��鐡vMg��k#b!L�F�VO�c%69id"!��p����lk�!�U����(&���I��y�vk�����~�#O��O~���O��/��OG����կ}���h��je��-W��>�诛�`��On�/ξ���~]}��?��?n��n���m�A��2�������t�6���g�qm*��)�WCf]�Vj�5��C~q�' ]^&Ŵ�$��vw��6±tJX�����H?,F!�T�7�Yj�kL��G�h�O¡e�*��p��M�͆���}�>$NJs@.&����*���_l7��Y�+!|~�jE�A���B��:u�>�w�8|XO �zv¹6�6YX@au��8��@�S���:��n�	ɗUb���A����EM�TCP���4�P��]�x;IE�7�[ÍV̈n7LQ�̚�֎PK!�-���t����jEk�%��|I���ܸ1�lA'M��u]--x�C�������N%=U�kkE�`���V\Ёc���) ��M%�l z���N ���lm��VK�d��������т�u����Q�契Ի2Fn�ԫz�z��j���ō6?E\F��M�c��u劸C1x�lb&�����WĲ��ptliiq�4�t���&�y4���+66|�,������HDc�mo��m��WO�����O�P)�r:�s{D$�B'����d�,#Z�es)�l���΁��,�0)ۅZŀ�o�7������S��7���"�,2���N��KØ[Z���R�&���b� �k|.�8#qS�|�
&f��w�n�:q:��P@�XA�j���f&�m�������C���L̀�x
k�a��q��'�eL��C"_MH�'��4'c"J&:VB��A=���8�c-^�.�0�����F�W'o��Z���mMp�������Ka������}����8<�`~yM����떄m"�,��069����MI��W*��6��s�rǑ����s+\���L�.��� %%Fkf%┽��`��^1�϶��vt��# ���bcSX]]�����>�@�`7�.ҩff'��f$a�#�.��مMIi^ZY�f
�?��{qp�)\c�f�h�<��p&�Oe���m��8xhP�@Z�2��]��I�/�w�.������C2�ǯ�='�aO�
˴ ����7�C�8��0ۈ.l�TL��1��{�g� ��T��%��ﾍ��5�9s7���h�;>�����]��VX>i��J���"�|n���T?�Q03�$��T:/��D+�F���h���Ҽ	������4R)�!bs�ns��E�4���u=vlF�]���_z�dT��:k.C��kv�U�sV���:��� ! b,�7i�����MJU�-y�]�4#O[���u9<t�	��>�];���G���e��Gi�g�Z3!�͋1�s3��uo���ZB6G)��բCoW;:�mعcN�y�hPx�D97����i���9�L�;��[��S �S*uX-HgR���h6��ѽ���S���ŔL���ᔴZ�x�6l��8�*ƗWP&Bbv�i�����*f����E<� �"Ɋ�B�WT2I���v�㎄v�x��ڱg�v������&�"!����t�ac<K�P�!S�BQ��V%"��N'���uww�����(}�����Jľ�g�\'J�%�ƣр%�8NS��t{]r/,�����h�؍2�&�������>z?���x��7�(�I�\�l��/Ur��FgO;���Ǳk�.<��g��Kg��ʬ+��}�_z�Ӹ�̽�t�m9s�XgP �uD��͙%�t�"F'g��B6_}�b��P�����#���%��R.-hu��,�E�ƅ�x��(��%ԍV$��r9��O~����׮}�����?�Y4l�}�տݹ���/=���+肓3���h%�Å�bE��¨�KM g�%`dl����`8���	�{m%���lV������B�h�dQ�����kӸt+�xՅ:S]Yx����YQM�a���,��of ��e0��<5&�W���-ǹF�1R��i �i�/LU�
SSih���0R��Hl�M��Gm�:�"E>����0X%��f-w�����?V4�	7f1�"�G󿭪	��)[U�����N�l:�r�ފĂ�Όz�&���`�a=�GQB2�bY�����++��B@�nK�!h������dr@�$e���p��!BҌMׂB�6TS0��/K`Uˮ!����ѾoB�-$�����)���̆[��׷a���&+��u��t�t&��ce%$eKK�m^�)��������&����N�͑��l��Y�@�����ꕪ��܁��vi�����7BX]�@._���W���4�~3�M6�#tu��U��L�s���)?��<��±�f
�hm���n�w���$}�zz3Ց(�M�Q�[�h��Lh�nq�ڰ�D��s����y�ZXQ9��k� S�X��13=���1����u`���fifˊk]7D���H8���(,V7bȗj���HhSW�ݢ=��m�欫�`����W�N��@{G'�>�@�V���v��<������bc+_SP���� �ž�;l�K��+8�9w�
�~/N=��}]��E0M4��9��X݌HQ�9p�����@�0���`umC6Tt�`�,��������L��&WW�Y��E�ri�����R�;�FXĲ��zo�7�H"�r-�C��;;��x��Z2�����6¢������1�bfa3��hn	����>�L�B�!98���-�������mª���݇�o� �KвA�+c�����-	ו�H���mi�G�+��2s`A�/���tw5a������Tč����H��d�����n�ua���������{�a{�vx�N��9������-I��7y�G~�mB��|jn	�ˈ$r0�=��ZLla{o3��؁m�ڑ�%����=^D"5�;wW�M!Ь�W��:�2�?u��P-�g\��7&q���SEq5a͌���w����=�r��e�OL�������,x�~�#���f�y>aS����x�Q,ą�`*��ӏ#G����q<Ҹ��.`dt
	R-.��5&����CljZ�H4@��:e��a��A�)bdAKr�r�a�{f}6]�A�ˣ���˿@)�]�,L���m^�����1��f��A��2Ӽ�~͢�הg�8ꅜ��R�&�6[���Z��:��=�Y�w��^���_�|��9�h��!=tc�PI��)�%Z�W%e�`>��tF]��Z�q����ȇZ˴8�y�&~��K����N�#�! �Q�
�v��QCa2��*���g�����H'CJ��z�e�3������x/��:�.�����S�a4���|�*6�4I����P���/
��/��l���Q��J�:J-�Pl�i�]D��\o�$������nh>Q��n� 	⠅��wH��1mH��d���Uz4���ag��	⠆��|N-��b��
�XGF �c���u���:���ƽm���k��Ɩ�lv����5N�s���xᥗ���.<6�l�x6�2I ���A<��7��_9�<�,����^�sF�7�/~�?��[[@?;Je�VK��_�	���X�%�+���R��S���<�}{�bL�0Q��o��:��������� l��J�T����7�Ǐ��4��3G��k�m
�?q�q�y�0��v�D�G�Ɣ8������:=`��g��ML����tvt�;�����p �6W7QȤ���ms(��<T�&�`mr��W.����������%�X�1��?����K�<�p	NZ���EE��/���	�G�&�䬑ʠ�?*X��u���dit9\X���H�@B�)�J$�܇HM����t������:�tg�j�>�Ǆ'Z�x����J4�"�bi�6�a�يp�?K3^#����п՚�aϱ��s��U�!��ą|���f��gf��a�;��-��(�C�����'�,7\q# mIkJ��uecC�
��4~`MMw�FT�u��߅ӿ�t؉X.�͍y_��*�!rT\T����dqjbl�N��H'���\\v�v��+�b���[�[䄑ְ�
s�X)_�h���&'��L9�`� �<9u�Gx+&N�bA��V���f��y-�0��H�łJ���Y��5d`s����*6�t+��2�1#�Dt�e�%�3q*�g9����>���Ď�\FFM=*W�#Y,H����	H&�*V%_���F�'ŝ�붣��S�{\^��4�~�o�^���'��x�*�B>Lx�twv`�A����i	A�j���E�1�/m�6#�(0L6�G6�B�6�u�w6c�@�fz��&��P��6B���ƶ�}r�(J1B���P\Rhg�ezMz���B�B���EO'~Z	��o�ٳ���78��N�ޡq?�e��N��"�FzZ~���Tsj���O���	fE��B3C�迯֧�f��W�II���Ct$+��+��I@_.b���ػMNZ6A��/���/�aqu���#��.7�i�)kޤ7!��ʡDH���KtیD�1�ɢ��Et!�&���+K��1���9�*z�Z��/Ҩ�3h�Zp����lU:��b�rs�!��`�;Q�V%���R�li�LkC��K��rB��8Mع��?<v����8nݜ:'s=}=0����hn�Cx��W��'p׉ؿc� [�Lͬ��ĸdT03���hmn[�T*���ez��Ed�ԗP��ఖp��p��>�3���;�s�Q���B[y��^�2�������#bhҵ��11���pL�CX𲁸��aѼ�	_�X]b��(^�=��u�!|術h
8a��Q�����a0�����&/��ײ��W�r9�
�y�1BC��i�"GPEZ�jnO,�X\�{АB*U-��x��̩@%nUb���'|-'�Be W!�͈N���Y����(��2�c��bM�@.:�4��60�fB~��������C�Q��_�����4A��_�(瑊�@_L����/}�RP?���ɟ<�����1����+% i����f�������u��$$8��Oc��G��{�Q�U� D�Q\|�2^{�_��۶���5�/c)Zq�s��!��kǼ�t^Y�{�.�|�ە�o��C{{+>�ȯ�#g���駟���?`fi3Q|\�.�}���W�l?{�E��/#�B&G-]d6��L��ȵ����Yϐ�]ʉSy�ܻ�oԜ�E����es�$P��/�N�E�ً�ih�4lj�*�%���z�X���h���-��'���H4I)��z�<�'5;���e���Z�Hg2�����燍t�"]֚���"M��Eٓ��?���(�|��x��W����t��B�D2E�,��?���G�����M|�c���k������`bbB8����|�_|��n����I`!ia�LJ�ڐ���Ǫ��j?~�g�r�*�2�N:�'~����	���X6��!�"�sPLOX�n��7.㩟���\IgF����~�
!`0��:��d�����6?�tK�cL�.�Gl(+���;���/\2
�c�����g��ѣ'��/M��8�\V|����bG�7��ׁq%�����"^�0����!���aA	�.3L�(��}	��q��i�A�i:m�
�K+�=W�f�&BU�詅$�N�IC`�0Q�N`T����	dՠ )�&���]%�b�5���U�<1�R�sc��NQ4Ž��t͎M�A� aU8J!@����r#`�b�<E� B�K'e���R��L���c`��:v,� b�:B�,A��'#qD����
��I`��*qA{�>�;(�_xq�P�_��D�WS���!��sEq��>�W��=C�h���*�!���9��r`aɄR��gC�h��v�����M�DƧ&��Rf�N�W�SE��_�@�a	ƣ3�#v�LC�������fz(��t`�S�)���N%�ҙ`�{Ul{5�C�={��kw;��*������2tu�=�A��hj��
XwZ�2Q�%���:�|�\�]~���T"��&�
�f�T����MeU�B��+Z�Z��R)L�,Hx�p��a6Q>�K
�րO,Ը��TTJ%����e��fKrh��+�]r�s��e#0�ӆ��&	��3\�ױ����b�$��Z�sW-N�@h-����2�|���9x�Za4��`RɄX߽s�:}"��Z��!�������N޹�]W��;�t@$����-�#Z� �.���&g������lQ������հ�����&��'yM8��J	�]�8�s ��8�� �T���-�{�&±�tKk���}�K�,���BO��D8��""������Lv;�D(��Q1    IDAT�%�p�S3��p	��1���nx��l��WQ�F�� ��ߋ�N��gRx�Q���(W����-��V:c(K�!��2�*&-������GoO����rzӉ�dP���Ĕ�o�l3��~}Dh��}}8�w/�Z�	����-�gX|q�5xȫ��1���-�hC���t�R�>����}�@�����>llf��ۣ��	�^s��H�e�G{�	��:�ަf�r�3��H�F�(�kiF��/��< Z�`}��.\E$�t�:z�x���1��+M�P2�qLO- N �ʔu�`?v�DS��-:� ��	���a,�D`4 e�Z2��7������~QƢCa�jb/z/��XM��XB&��c�S��V�^�sSx��O�^λ��BGj��(d��I3u���V�2-V�t���5��p��v�w��i )�F�V��b��U��9|��	|㫏�}�"��9T(�����M�ݥ
W>��&�Z�h���H��f��/�^%^c��{��ѷǏ��hP��jvf�?�~�����!����H�e@ų��X��kHg�H�Ҁ���x$YN�������'���<�),NM���ۿ�3�=/Ti��!((�ѱ� ~����о=�55+��#��29�R"�(����F��j��`R�C
�9�$O^�3qo�z�0A�v�Z[��t�����52�����RQ;Y�+��ަ=��QQ�DXÜ�rQ9D�.�<y�F5T�VV�����A+��x����#h
���pK����D6S���Pf��_��8~��x��g��K/au5�l��r��g�q31Գ[8vl~����#�/�q����I�tu��_������n�cy5��naf~Qj("��l.��؇p��	�,��R���E\�x	��v����<��wb�Bɼ�u�O�B"�%��K[g��q�w�zpa"�����+._�Z��rc������ׯ\�ڼҿ�Y(C��|�G/|o=�=h��D���1�PىQ�C(�`*���v;�n��y���F�n}��Ò�ZL�@��]�aW*�'F�~���l�a%��i���8
F?�t�*��&ԓ���22��W�W���h�*=h�0��q�7����S��\��!`�(���E����ȴ�! ��\���)'!� �8�Ҍ��T@�����ZxM�Ŗ�1-��7i	��A�q����s��f�����yHK�49��Y	ɒ���6�>��'�=ІD���L�lQ����b��/,�f)ǒ�{��+�Aq5P��[�#�5��� <Su,��I��*K��?��|�h�Տ�XX��8޶ٓ8ru�a+�`*҂��P(��:���T�!X'߷Z���Ƈ���[��*tU�PU�b#j��E(d61.��5�y5�)��0�M �.�cE���Wk
�b(��TEg�@��#��v9����˂&��ѓ���h=�JbQ�0���f�)czN�.M6�ן���{/mO3E%8���2�g>=�Mf�p�"v����d�)�şѠ�sڳ�q�vv�J��il��D� �t��V��t��0O�h����,(��ً� ~�"����"�
ŲXwwx4��L�K�[3X\Y�����,�F*.Eq�|^�Z��Q ��G1��.��^��dFoK@�C����V�Ji��<,��U�"I�O� ��B,�C,���d��*�ޒ�N� jOQSJ6�s_����F_��u��y�g��]nй�,��M���a��K�u�zc�=Ai��D��r�T�U���iE:15�D&�@��w�BWO��\�F\�x��7��@ǌ��"��lD�@dT,Z��ߍή&�٧B�6:��HR�X:���IB=ӂ�De�p�Չd�r�s��z�]�-��j��N[BR�r���i��&S�B��_��jq�a���mC��	�` n��Y�0x�n��XVqk|k�0
4	7�D#��a���bh�;��Hj9�x����y���0�9���,R���8qtz[�ddݳ���Q�L>qEj��([Y�q�ŀ��0.�{�+[0�Z��3�8z|����0)�fM�
H�2�PJ_y�O{<6INgA\d:y�t�&�|�]ds5��Ai��[N�3(�P��)�69s��{N�=s����N�_�l�	:T�[�/e�}���P����fA�ˌ��-��ܳ@,
��&E3�5��D�Z6��
/Iy�)�Q��ĽN
X���J��#q�1�D�\M=��
�0���h���Oa϶^i2I�I����ٗ��K�`#A�n@2��E�C��':�g�BQ�
"�$k�	Idg���G����q��y.i�I�Nb���~�Y|��G2�Aw� �'���Ь�+O:�t`d�%dIueHu(�3�\g*������~��/byf���{�h����G8����:��v<�_ÑSw#��`an#�cjt��-���1����,z"�L�V�I�
��6���et���D�q�����6�I��|?�_���3K��F���$ϝ��C
5m ���|ѭG���%�jq8U�k����>�|��_��I��l#���XW�|����������e`H}uo.��o����S�>4(���U� e}@��%�-��~����=t/�����_�)��c�у���~>p?���{�^y�"6�	�5,��"�u����ß�N�{
ӳ�x��Wq��w�݊���{�����u��fp��E�{�=�ܼ%N��;y�Їpσ���.,�������λ��ri��~��������q��~��޿��O����q[P7�$�������R�P �"��V�U�4v�\<�;::��x#��V�z�k�|
w�/>�
a�*��B�\G�`@8<��i����5j&��dn+Z��6�0y�U�Cs��"6&7�����}$w���#vu�SԐ ����@6(�վ|J�wr*���	���A	(�R/b�������,�AA8O	��e��>ŉC�����4�{l"$>[�eqſ������Uʤ[ُZ�vI��A��J
��g�a�8�a��K���$r�,6W�XZ�W�T�,:���)-�Л��'͈j䋮&R˾�_�_������7,j�<�ُ�>�q����ŭЦР��6e�*������M�?��� 	l��!W\���|fe��G���3��%	Q�A��Y*ݚȏN\^X��� E��K+.G�E��9�#�|6l�]�]kN��'�MM-�ZhYA�oE�E���:�yoMu �ΠZ��	f��,^�0[l
�����!��i��,`�(����CR���}>�V�Sb^�|Q=?V
���$�۲LԼ�ޭ�{=&:@���Y3"gT�nT(�6�dRE/f��$�%��(��x2#6��r�jE����f�9q/�oBo��M�%�uf�æ��i�4��[=�^Ah�'��q�^���:<Ru�hx�+��'���M�wW6��Ax+�b�"Sy�[��L5��1i��E��3�6I�S�ӈ�
D;�4V����j�Ey~O-EDdJ�3,V:���B�h*y�>��=�r�^�B�����1;��HtK�(F�wv�%؎`['�VW11zS+��雭3;�	5A{u��.��߱�f���cq9�X2�<�w�,��r��^�{�X����B�h�#�c��y��5�]�u���#�$��
��(�8�i��ffV�������&�E:�	�׆�}ؽg �"]G2�6I���R
�n����ˋB�C�4���Ut-ط�W�W&��Lbf�ϕ��.�!$����V+vlkCok��5
���`y $+^J&r���\��lyq��Ǳ������.V��B-A�:��79�`��>b�&x�~��PP%�L�TB��e���WFp����&�����\0[����	�}堅o$�W��R��Ybݍ�u�A��yf����{���1�E��J��f�&�f������$�Ne)٠�ؼZC0؂�;�K����4�Q,0y�H�Ii�$I��J����g#��qF�Ѵ�Bd��Tǝ�w�؁]��Ȧ2�px|r�s��q��A��>�V	�4��<��t0T�8��b1�=���}�Q[[ՐΨ$��xB���z�T��V�=>��A��ģ�	�+�$����B��"<���E��r���7���?�YTsy������߅�탻��X�h��#_�5��013���0'0=:���Q-I�%���Ј��Os�s�Ć���Fs���6�W�̩�Ƽ��%:.j�h��g�_G?��.f4���X'F��:)DH�gP=���f]�F��"��r)�Ώ>�|��ay��f�}Ӫ�t��w/_�w��?���|^?Lz��i�Q<��/��p��qi�~��p�֤��Ya�%-��l�LǏ�Ʒ~�wp��3x�+�����q���9��{_ǃ>(z��^|��s%�$��m��ݔZ�n���ѝw�%�����o�@6���>�1���~V�����?����E�H��*�g��Ϡkh;;�m{��f0�=
˧&�Lf�G>����_R�?��!��#���w�ݫSw9Z�0ڭ(WrR��HW�&���TJ������+Y)�yx0	�����I���=;��O'��G)���@9������.��2<���8wu�L
p1��iF6�(.C��"PKJ(h�E�5D��*-�M%�dQ�H1�&xh���o}%��L^��7_O'�w6��Ft����3`�"��WSŁ���2�{N.X�K�]]���{Ni(��MQR��2I����$\4�^P��r���*b@�L89Q"[.�a�{�=��<��قx�(".�3�$"��������.i��zA	��, ��AqaR�FC�>�
E�^<�T��3<T�pU=X��}8�鏠cϐ�.R�/]Y���>�"��a;�I����z���X�eI'0� ���L&�]"�P!�Ȏ:.u:�"�ͩ���oA�H�G�$>�174���%#`�YTE0����mK_S�6'�,�gM�&베�?�to��q=R�O"i����>�B�8�d}�O8�.r���1�Grڙ�i��W2����U\Y��U�C��(p7�ܨDcC��N#2Y� ��H;p��ؐf8�7��.�Ox$*�C���g���rr�C�Š���A���]�r¦�h���,�;�SRق4�3 �A��#)�D��*��R�u(��4�rU�!&N����t�X��'e��"WB
b�V@PB�`Ӓ�q����Č�i���(kr��FHgd��	zY�aC`"���Ǫ�l"x�X�kQd
�Qۡ3T����^/�����/�&�,$��o�m��]D��B�8�7	����!��!�ɳN��*L�Y���^"��$,�"�.T�5[ܘ�ץ����(6�����4Z8`U�V���c=�[��q�`2Vhr��w"���!u	l
7CId2��l��dfF&��z-���6��4��8�^�3\�6�d.#6�,l���i'�ǜ��y�l�^u�$uc3�յ4�
�[Q,0���X��:��	�-y�o�\�Ju$h���
�`fr�Qح��DC5G</�l6:�x���G_7Z��&o��
9e�ۘR��Fˡ-	mF�&Q%"o�Z��pC+����缑�9��U�C�sC �JKH�kĉ�m���2e�Nb6]m.�N�4��;s�&�Y���Ӿo���l_�]uY�-w���8W��1��IH���$�痄�pr 	� �``���^$[V��UV���w��7���o$��w�9��˗�-��~�y��ۿ� ��",�R�=��CI�RťW^�{�y'�o܀'�|�}��r�"��$�a��j�D�V��Nt�h��x((��穧���U-���a�s#�,�#�AZ��"jk��6Y5�݌r|w�6�|.NH�� Kd��LfE���o��ׯ��2�Wݝ������c'u~�]���ʎc�:+�ƕ�nD�-A$;S�Ht�3�)�����q9�<�w�{ߥ��]/���|��q��Qл����Տoy+�t�m�]X�d��2�siL�C9�-��ȼ�F�a�g��Φ
��Zرc;�m߂ٹI����j�i�g��#��%/�SUS�g���nQ��6@C#���#���csF�O��@�%\���V������lހz��1����I�\�[|&�>����?�^8ѐ�H,aaa����˿�4�]����#���?���������'��Jn
�،�����oy��?��O����ؾ}+>��_�w܂c�f���>���Eݎ��c%_D��S?������������`f�4|��q���� b?^�s������cs�6m��`������#Չp<+�p��f�����{n��g!�;���o=����o/�,X	�Q;�S�D -x��~'{���v�P�\y\K�ZnY~���f�ܱNz�Z� T�A+`#O��_��^>�E3< _l:��ަ
��(��8�za'��/$��a�Ž�D\/��VTz������`#��	`1���CI��(d���7�?w�

c���3Ԁ��Gw+Âa ��"�n]ʍ>S�ؠ�8S�g�r["��,Yl7����^䊶�=w��m���:� /���@V,�T���N�����z�!�R�]9���Դ(C��)�j��QD�F�@#V� ��O|��!j�F]�.���D����������{�6\��7a���X.�^Zԟ�͗����Ռe�h0��M����69r"��CC�����@�����hW)�����<����C��V�?�A�$RGE�37��L��tq�k�6+f[��~��C	�:=�ikZj���h0[=6�>�Q����hM8(��Kژ_�7����)��R�,�.U{*#���Y��Ay�Xx���,�Yf6��9�n8�Z��g]�4�b�i*@�����D/�3o��5��@�`A�2B�PJ�٠����C1`�&����O��bW��5�5P��͜o�Z�Lضy�Լ��!�o�{�:lft(�χE���hX��fiB���z|Q�Z)r��TQ%�ؤۇPb�R4�u�e�h֋Z��Qi��s���D���h��
<�Һ��{s�g�am�+Z w���
�a�7�h
���jF"j��K��B����T�'ت���`2��/%����A�9,M��� �}�HZz�,i5�w�p��&=�r	���P�v0�N���
��9�ZPL#�c��%�k+K��ٙe�Ѱ�.ʤ��DAp.M�Z6|�z	���������T��ߝ��N�aBi�+���YA4��:���PS%݊����J=���o]�l�$Â�؀�/��6�[=Kjn�iY^��2�����WVLNN+�Ո&�X��E�]f�p�$����
�j�8�
)����(��f3n�<��0�פ���(O�%*��dL�}������@PZY�Eu�����U.�k���|��y�V<��K��/|'O����&6�j�܁��aG#��eD��E~N��Ʊ��K��z6�Ә9?j���ֻ�s��t��)"�B��YN�%�O��Ԫ���a."���'Rf�Oa�S���M�OcrrR�i(Q���P.M�fqI�P`�+$���K���^�vѺ�[ai+�f�Pv
�����E\y��(
x��O�[?���et�^���ĺ�硣 ���̯�_�cf|5n�_DH5s�jN�'��̥IA���p�mo����������ߓ-4�wHEL&��H�+/�Q���12I���Ya�MD��"Ƭ�<T���ڪ�/K�H��u���/|��x��G�
�X.��ze'�V�ϩ�����ǃ�x�N��>���Ht�Q�7�~�4�l�7��]|经`zv�2s,��~��"J�)\�c>����w�O�x��G��_Ņ���G~����[���k��?~�GP�P�EQ�5�[�ܴ�?؃    IDAT�¢������\��������.|���C���?�2>���\��*�ƪ�u��l�Y�����!����6��̾w����ȵ�>��'�K��9v����9�y����7�>��|�2���ux@D"���j!�������7�;�߂Z.��-�!�j<���-�/?��s-�b��l8Պ�+]� �A$�M���-�r������&���]����Ã��M1�fڕ �㑘�����^�,A�|i**@����h;<�OW����F$;�$Ŀ���� �J�rQ�RKx�
�$��jf�D�~/�6d̢'�FOf�F�F�H�Q�R�B^/2����7<~,��r����$5��D����,&�Cyn�8�D���lhm^�	n3�i�9������m7-SM2i*�g��=������ʛ����M�V�Ȯ,�����HF��j)�nR�;�u����7h��6�-�]�����?Bj������OG*�zdE�&T�P�l5Wr���,5ޖl/��S��tP30 *@տ�Q%sr[C�9aT&Z�	��{�}�3St�	�ͼ�A2u5_�,y�������ὨU
J�֟%_���p5p�58��
?�&�̈́�������9��<�]uǸ��j��iX�6�����9�Z<0�Ǝ���61���2�7�7��:��A��f�V)�J���/�w��&�t��FL�2�B.����Y4�#	�9ģA5�eMDY@:Tͪ�pR�8��oy�%��2T�J� �kR��U�d���FjŇf i됌N�-*&ݎ?'[d"R�yZ������K�W/jlm�4R=	���+GMן�)z՗K��D�u��C�0?��^�&�����K%c#IosO �~4&����"+�j���I�(�ѩ�� "���U�+@�;�79��Z����0��PY��I�Jut`aiY֤P�H>�-�of.}$_�B7�,�in|� Ʀ���~��`v1)"9ʁ!�Z2��#���F�l�s�����iA[�@V����D'��� b�!���S4�����^i^������:���ޕ`�)�D{��kŌR�6�[��.�HM��p�GGG��m�\?�
�i�h�3��'��ҹ��!��=�Y�\s�Қ���i����p��p�s���gn���Q�I�i�>;tZ��#x�9�"�o�IW���@@ǯM�6�o�}�x�������͛���W~�� �\���"`	٪ɦ��gw��j�Z��Q�@�x�ב��@~y�����2�q�,�lй -S(���`���9� �p����-9������u(��������9Q�]Z'� -q|�9�ynK�@@�c��1���SD���E;�����^y��8�ry<��nL/g��X�����
�;��#g�]�ayf˳�(+��5��@��˯FӤH�5oX���މn��h�|��x��Ȏ��0ؖ���-����<�^�g����Δ����E���]:/tI�=.+z{�e�*������jUsN|����o�	:�q�O#�!�4���8�����?��#��hI���˽�)U�}�7n�����b���x������>f�P.q "�k ��WP�O���Ç?�x˭7��G���
���5���`�ރ�ߟ�J^,�}p�a�h�"3R�BY�B����Ό�vJ��]w�>���~���~���OK��G���y�#�K�#-���*ٽ���}��8xv��/��e�S���ӿ�����ɮ7{:R ���³�*B�e�����D�AH>��X��/���j�,��&��}w܂+�ߊf1?�l�hoǭH(�b���<���W0��b� _��Y��>��~���舲�sW���1��Q�,
l>XM�e��>1���R�ϰ�%��%=)��:mA]ᨉ ��酅��V:4�m0��C>�f{��^bB��5M2����8��T�qs�-�æ�֋��FtC֜��%�j F�PE���m��6�G�g��4�VMf}�|�B����ۏ�҂I�j9J��zk��Y�wؼ��D�ܠsf�;�4�ܴL>+�Ʉ6QCд�ܶ���:����ZI�$�)�Y��60�)�Q(���`T;���Wu��������G�� t�`Z%�<JW���l2���L�	�&�N@t&�AA�{�5x)�m�q��ѬU
���Ó(/� J�6؈����nW�M%���pN��y>)���(�2|�G =�2�s�.u��E���4�d�D)�dR���f������-n��F��t�
��/nQ��ƶJG!
��s��v#�� ��8{ˇr���6���?�6�Q�)*f<����1�RC�Y��J�!�G���6�<��昴lY�#����a$�ğ�&�G�!���Dzl��!�M0C&D�|u�||r�hh2���N�mӔ�TqK$G�6�\��׽f|�9PH���F���*����,�3:SQT��0�%d�M��IX����8�g�ͽqә�1t%L���=#-(�H�"I�%��DQ-��8M�?u!~ګj�!r�B�t�2�RB�d�ƻ��e�T,}~ۼ�u�8�R�c(gy��h�Z�]5�Y�#/j�Ic�P�)Jd��������7�U
�� �~��2�z�j�Ac�h�D�F>��J��VN����o�����/�֘�QU͓^�N�s~�]�.��c���jrP�� L�%g�4R��1�&*�jLc%݅���r6��@�:)Z��Ս�-FUc����G. �Vr�#�.包5���B�F����.����T�F�X��le"-��� ���:,`��a<���b�PH5���6��R^=����Z쭤���s��|����w�i�c��jlY���FXMf
|_��2"ޚB����4lߺ7!�YJÚ�a�u���;��; z�	qcݥ����BKf���f{yæ���ަ)�}gM�3Q#b(�̠�BJ�N�X@��{4*��϶Pp�XX��%��w�}���:�t��� ���cf9�t�.���r��&pjdss�H/d�O�!���<wGW'��D#�\���T��Ƚ�o�Ϋ����jى~�{��'�W>�t��aˏx<*��-(�FL,��[>/�Ѹ�a^S��D4�H<���3J	����M��$(�g"e��E�����{q�[o��5�ܐ�*�zz���gy�*x�'��?���t�Md'�X0*�����m܀����b`�*|���#?x+�<�%.$�{B�(*^F�4�+/;��ɏ���Ɠ�����������Ν���e\y��xn����	5�
*�`�P�YĺD��ɜ֖��&i6��߁�����x�����Ñ�y8M?�%G?�L�4x^r���	s�h�J�Vzf߽������怳��e ��}������<�o�o����P�mį|qՌ����.��/k��pIh�A����K��ý�܄k.ڦ�r*�e��1SbkMT��|��#84�E=����%$-�ZF�I{ <myEQ"��M[��\��BJ�r���E�A�mg�e8�-�F����~�N��4���	`!��M!���X��OD2�|n�R��-�K;��4����i��a�4Dq~��@��t.4�C�� �bLbW6ʌ����͇��ؐ:�@ej�\w$�a
���� ������C�����FDcnRi�l"�m�� /"C��]/y�/-*��V$z��7�cP$5w��Cv����[�2Եi-������m���W�#�%<��8k��4�E�Y@�y�&��D���}�f�����с�M�(o���0`�GII��2����/a��h��6_����E�
�3q���Dl$ƴ�`3xE�����jñ2�
¡����\�����s�g��/�r��w�g܍�l��ś>�L妵^-�Q�[.���d�5j�p�fЖ�����'�^���D��D�q�#��Y�}�EU�������j�Ԕ��7}z����cM]:� �Ґ�]ұ���M���������2r�� �_RY�G� �0)�D��8��b[�]5�VÂq&E�U���� n
e��ƛ��*�"���O�,BFkb���50+	��}j5��wL�B�e���O���7Ä��P�`1�G�
-r���L@	%TK�T���hu)��=#���Mɪ%����"=�iBP1�U���.�բ�il.:G���E�8���"e��9J�o�	�E9��z� :9Z�6�~r�)�� j{�/����Y�Y�09Lb9Yb?U�O�5ekɤ]��J��\�2����N�FAz-_�,��&:�
�����ZS2Z�5}O6�^ݢ�pT3(���:);<t,�0� >�Ǚ L���0�<j�jՊ���`(�H��_��6�%>i?�»�M�~Y��^�nO<~.&F�B�y�hv�1�d��m�U�]a�X�^c`C����ĥ�D��$,&������C5�F8е�uh�Q�~�py��B�I*Wv$�A�c[�J��Zm1�������OV�>w�݂�Q��aZp�RV�%�o��[Dve���,��{�ƚj~NC�j2T�}~�@�"�ڌ���A�BX�u6�w�j��C��2�kg���1��o�SNXv:@]4��ͥ�Y\{�e�붷�K.Eo� j��Ɖ�S�_�tΑ�r6W���2&�g$j����%N(w��Z�hB�H-siW���ǭ�݁ށ~o�M$cx���c?��,Ź�d�O�6�|��٬���4 �����}}}:G�]izD�;u�$fffdMg4"q��m�sV��7N�:�^���|#��ηa��u��Q	����O�Ңv��x��w���x�Ԉ44<�B�޵J�t�e}����OcÆx�����o>�م�B�P����5�[�B��᪝;�@p�U
����;��/�����k��Sϼ���×�o�1���P�逇C��l(M��	oÁ��Cqz
�f�r�����z?��&��{����82�,jhY�[.�嚋1�<=~�|�s�
���{�]�㫿��#?3��~�;���G?�T�m����j�RP�m�e��U��-k��bq�YL�`�A�@P��rp������7`�-h�����6�<��&0�m��?z/�A3؋���Z�ÄU��
q�fD|�yz�k����3�%CC+�~؄�gh����i'G����ni�ς�B�M(�Tf'03���k:I�eG�B(�M4�9&�S7�<�,�W6��@��B{R��M��-���V��S�i"�����)g!�A��1#��Km�4�fkğ���6���&e�NDvA��j����I�=�����N̂�V5�N�̽�/"R꿙&���6畍���t
����q�]��c� ri�K���e5.?&q�g�U9��g�-�(ݢ>�q�����/b���-_(W�Y�Àd�8�	�!���h$���k��w�i���T�<Z!��M��t���-�(Έ�9����CK�#�`�l���Q,�]s��J��͘�`�&���������,��%��-�	l�،r�d1��L	��@��Hػ�M�a�����(ɘ۠8�r�;Ք3p�T����BÁ�0�6���pT�!b�!� ��e&12����y8T�0iZt"e�Pn ���C]
t�j��<:�Pv2
� ��ߢ�ֈ��F�X�D�h��=�������X�5Ի*GhQ���4Dl�j�.���C���#�rCm�����3��
�"-Kt\�-�}Q�x._��<��5Ю]V�u��D���p�OQ�����e��P.ԋ[~�Z�~~n��P���t/>��A�:Ҍ���+Q9 �C��e+��>���{Y�kV�#�e�f��Ơ����U�+�C��;�>j$�`���"�D��Z]BL�ظ���AO�O˧����(�p U"rr�e�f���W�F�M:�ʭ:�#~m��`��f
4 J����?��Q��55k�45�&�rAx<uR|Ҁ�}5����Hq9�:��zC���:�BЌ����l��=.����k��eRp�DʀY��9�^��H����	��#*��[�Zfx��0����ni8faq�`t&�\�_=��z蘁 ¡���hP�d�G���sOʊ:	��s����-2jR�ye��d��J$4��+G��{6P��h!�%-c[�T
�䳨2JՎ�\+ �]@��Aw7֬Y����lX�w>��$�P��,l� t.��6�tv	�6����YR���~�w����Z� ��|FAD��6�A��p��-x��������r0x><|Ͻ�'��`��D�Ğ��|���RA)�o/ay���u���VQ�=6-�cA�^�+w�$Y���شa/�z�<�(B4X��j��V��"U�b�f�D�Y:4���r@�(Ut��H�3�������I�\V���Eijj���{ϻp��;���%D��ċ���{.�l�>s?����].�����������̧�oz�8v���_�SϿ�R��b�_+ m[>����8������ÖM�x������F�'���я�]q9�۽����Tn"[k�iZ�X	����0/�,P�
W)�W-��4�`���{'���7��#O����(��X)�3��홅�q�F';�A�P�|n��,-���{o���|������o��7���|���D�M����oӈ��_f��IA�om����1Y�ZD�U��7�o��m݈f!��y6�I�h��򂡧ˎ���~<�w�� |�N����-
%-����;̦҆����[>��_�L5Ww P�:�F�NN�o�P&��.2���q���.'�&�X�E���\mDCQ}/B�,��S�E]l���T��X.����$�L�ж��>,:Ylk乚	�nֶ'��6H��IS���Dű��%7k�>�!#������;5����&y�Z!�����5��G^�g��@��B)�m1�,Z�h��4�����;oEt��ˋpʴ�d!w��\�d��������S�\q*x�Q�{�}(U�5j�g\Y)aa1�f�R�'n�I7����>���[JD�G8L{�rYK+yC�� j���203}����.�� �E����%,,eP�q�ِ��[.#?=�_�9����"���������V�Nߠ���3�eɿg2uM�Rt�6�8�X��+�'���'%(}aa	�|	�B�b�\A�|n�
p�%B����ۍ�N��ְ�N�{�g4���>і���p�@�vlb�ό���y,���v�.�%�?@
�^��7�@�A�
*	���Cޠ-�B&+���r�=�j8eb��j���ry];�ъvh�+!��[/������p�Mݦ5��m�[�е�L�m_�\TN�Xmږ��,�D!jB,dO� kۚ�H4 ��=�_�(fs�ؖ�RY�)�P�旃�Ϙ�CG"rQIǐ��I�B.��,��C��?3+������3��q�i���|YK�Vԥb
�(5ԇ��!<҈��� ��aN&�]��H� IHȡ�KA�P!�Z���	�}��WZ��!�M�(c?*�*JԼ��6��2��K 9��U3�i�����49��iRg6�<_�t�i&�^R68fK+�����:æ�K%:�q����uBD̟��1�"6u�K�N�6F�//��P/D4Q�*�C���j�Ԁ��'� ����@�f��?g_�@�o�Wa��u��1p-BWď�SG����0:�s�g�J-�(�e3�e�h�^�C!��v4�`<�2�txF+�� JZ"��RK>٧��7GzGN�C�A�2����R~����Im�
�2��-�4h"�Ƕ�Zϔ��@T� f�5蜡��A�I�	�!���}874U����s�e�]K����	������{��N$�](ׁ�{^�W��6�B���8����Ơ���9\���&U]a��뇰z�Q�:�f�n�:�ؾ��R��    IDAT�O=��DXZ�r1�r!+����Un���'E�=P��ש�҂fa���8 R�H����0����,M7m^�o��0��X�zz{�$��".����!�aai�_~	�Sҗ,�s�aE#t��C����	�s��ճ=���k=��GN`a>�/n����x�ݷ���CCC���{?����?ę�q\��J|��~W\u�{�����#fV�(4�f ������p�%��o{eO��|��hd�x�]���>� =�_�֏�\
�P%jO��J�"Hi�;��,��"M7W��w�w�-��3����|ᖯ|��ϕ}�5v� �,���A��6B@�(�y>��<��Ig�� %����c���͸��mRg�5َ�AَV=X,��#{�̾Q����l�`�!Z*u���P�0�V�g�6|^�f��9Y���)BԻ���,ѫ^"M�|,�,�����Nӎ�'i
A���Uٜ1����P���k)tS���QY��ӛP6!0�l��\��\�1��AY��)6� �� ��F�/&�K�R�)�B;̀�CE�qE��^�M
6��J�%ߘ7v)(����/a��)̝>���	%c�����n��g�鹁@��V��@ ~�ִ�QI�;!��7�}�k�1�8�M�,E]t��1��3ĨPT��M6Y�*��tD��G2F(l	=bS���	`y��ӣ3�d!"�0|�:��X��)n�yH0y����<���dJ��[<I=
�5�,�R?�{��ۋ�nF��G0�U����
&g�w�+���M�6�!8k���I6�-#(�@��Md9/>.��"�t�I��G&159�期?[�"c�@��ukz�Q{��_(4P,;J��gZXZRW����lQ�;:��NX>5[6?|�l&y{��'�(���c۶��������!��`�c8~jT�.��b�Sw!����6��� ��*��
Oc��IubU_��z��5,�������	�"�a5��I0K�'�x|H&btm��I�Drx͹��a��,�.�X������*"��i�I�!o[� sJ��i��n; �nZ77�R���3FgGTHd�X�[�R�A$�a��nxP����M�\A*GwW�6�E��J��ȸ��4�
!�~���S
 [���Ɲt/�N�Ye�':
i�`-!��6�"ǥ
��&�\�,�0uGB@C�2�X��TK�����{ܐF���a���A�ؗq�a!DM��Bht&��7"q~)deJ8jw�p*���e&h��kk��%�Q�bFN��@�e�%��b���s��5)���f�^�	��>+��z��IdJ�M��l�	��%�d)f��z�����]T	]�3��hK���P�H���t�PO)
�&�K"�58Б�Ntܧ�h���p+�!�æ�H��<'�� B\'<c�a��Y6���L,�MY�&m/RA/�'G������tg�I��cQU_{- h�����`�d�PK�:w�����/j U$M�ҋ��r u�P+"!z���8��ˮ�.Y7�Y7�5�|��;�^��	���@`�_s����n`i�>�kt���h�����>g���j��`Uj�P,�1?;�����?��~t��}�K��S�Y�9pT6�t��3�3��
RC�i�U���t��'���up�uo����p���z��z�{6m\�M���=8��n$�ADI	-d�-zH.rD"H�#Zh����NkU>��A�<)��Ւ�.����m�ؘ׆�3�����r6ڰaz�Rj����γx��4�#�H"��ʋ��9�;���rZ��y�%&=�U^��E(�}�z�s߻qх�05��3�?��=���>��Uwg
w��v���wc��a+�y|��G�/����p��;����5\�����գ���g;3�\�!�{�g���LGK� �ݛҲ8Ш)c�����;n�'~���<��c/����m�e������1E�V��斅�F:;d��EU��w|���w�v�o�Li~�����=�����UV�yN�l�m&��� ����R|^�#N�ⒺQ�;9l��{�o��RX��J�<�=��kY���[ �����)-+j��-����=R����p��:�hjN�\�a��	���;%�W���@�X�2� ʹ�M�����b�B+��X���S.鰩)��� ړF��$������G8�@,�B<��(�m6e+�
�̀6ܸ�^�l��cN�NM6���:[r>��q�|�k+A�4�<̔�C��,���������'1u�Z�
�bJ��u�]JԠ�_�K0A8<b�ρ��4IŦ��� tN��Pۏ�;/��o��ս83?#M����4� �~ �����h�MD��6�BWR�������Ё#GO)|J��V�0�����;�f�$�)D�aD�@���
r9���`l|
s��j�9TPP�ᗗ#� ��D�N���B_��l�@��B��9�M���^D�v�?} �m,� ���RU���SDg<��kp�%c�'��癜���ѓ���UBAu*�Ė��~x-�QK�\:����Ĉn��"W(��ֱ��"��7թ�c�@�1Z^fHj6K&����C�O��СCr�ڴy#���da�XX^)��Gq��8���B�J� R�'�cx��V��[Y*adt����^��|��Fw�Wԫ��<}�YLL-�����[ab�;Q��TJ(9i�/:�<D�6*��{�vu7A
�9�zQ(8�dȮ0!3�Ņe��@$�D4�� �Ŏ�<�N��=�Fn4
adc��C�"9Ф �wJ��{{;0��_M=�GGgpjt��_��6�@6��H�����:�qY�+lByƧf12>��SG��O��
�m&)d�N
�������m(%�1���B)c�mn�xІ�� I���@(�����@ 5\�n��6_�%��V�D+R�'��v2�R>��:hy�.8⢋&����:��4*ED��6�Xɮ耎$�BMrقI����SB�b��H��!Fa;*����WS`\*�I�F��8M4�M�i5��xL��Z�P���^^���3Pdˁ?�蔃��l�is�4bkj�b���i�[O�ZꏂZ"��6���5�(:�=б�Q��c�-�(����U�Dr 3'`{�M��Y7?�<iF�En�A��r1ۏ*��'��'���8G�]Kх,jZh�`6�DUxﭐ�$�l��5S�`�DEj�d�{	�kDݘ��d�N1�q�K���V����A��2�b]})Q����0k�hl�"h��B�
��@k��3HM�ԡ=�7 B�R���C�;����9�!I�]��6S�qD���-��b)�\nK�sz���^|�T/İ��q��}
/�rDBu!B���!{$�P@]��I:�;|�֭�e�\��`߫�g�^7�%w�u�W���W1v�B4�`ѬWt�)���鍾�l1y�s��AW�k�k������\��@����h�P��B6�F�RVƃ�j5�K�Sd�[�?��ՇF��L�����R>+�l�y:�L虛��G�qp���y���`f~���2�~���7�[nƎ;t���x��]x�'�������V|�����{�u����W��M�����/�na�~Y/8�_|ť���+�th��:t�j���V��/�_K�]/���}��p��8���S�mY۲3\I/ ֑���.D�V�����,V��Үw�r���^��������EŭV�����̝���K�A�g0�هۈP)���ف���QO@��(��ڜk��f1�u}=x��7�査aN�6��s�����Ș�ރ}��� ���^��"�c��n849{�Zh��p!8ׅu���6�j�9y�p�d���(��^�(�w�p2�*(e�1sf�'��Y-�UuТ�Z�d�.D-�7]�n6�Ąe��ۂ�v�`�d
����n�t��G>,,�ZA��Wu�ׅ�6�2�����jk(�fڷZ��`Z�q�ǈo����^�?�ܖx���p�yQ��>�����a���h���Pk�S��i��t��k���p���4ˇ;/��~;��@��.1�;�Oh²<(���!ҙ(�ꊪ�*���z�"SG$dÒ�;s3���"zc�3��D�66�Ī�x=55��H�@P\T�QT1�аTffVpz|JA(l�I��cB�^r��L��דĪ�P�G$�T��
896�#jtHu!�l���T��rų���6���l��U��X?D˽$��{�Z�PǑc'p��i8��z�fh5�ߺ�D�BY�U��ss3�}ʲ2�G&�G&�hzfN"�������硧�S(ii���q���SiG��c(��oڸ������:<���z\�m(�B�it�-��D��!�t'u�
�&N�k'O!�Oc��\z�6�R��5�+��~�;1�F�BG�_��|��U*g1;7�5�{������N��%	��In�}B�r�U�e8e�b{����+�*ہ)T��a.���vp���c @퇱5$��6�`¶]�8�z;�ۓ@���E�U��-���I���"�! G��΄�p�'�]�^8��T���]crcSS�n�{��O��������k��N��+���*kl�����$��$�c&���Pn�1�\��^G`j��djwH25ե�ᗕ��{���Tu8\)ע���Hؒ��;e�IW`o[�V%���_R�u�/`˸�Q��+ ==	D��T��Gb(�+�����bZ]��V�F_o7l���,�FƐ^)"M"��@�b�QA"ɍ���p)6��"���uY�n=]j��l�3S�a�5�#��0:1�z3�p�[(�'Qn��NsE�� �<��#';l2gHK�A�C��N���ӣpJ"�&}Kj9�5���=H��:#�����c4Y��p@p���ցH��D�2��ao	O�������(j4�#�B8�U)�K�-n�#A�����b�b�J�n����Po����	����w�B	
b����᥎��0uAoC��R!�5ëq��m�D�>�1�5�f�>�p��À�ؚ>����.�� }�@C��\5x}?v�"t6��]H2_��y�PH�<�r�dV��i�w�u��}J?�[Q8�����
�_:([��}>[��D���	ѫ`8�?�%g�Htubpx���.-`rbJv�<W6�J�׃S�cf��ৣ���'D!X�NW�lQ��効�V��'b����@�z�N���I�V��-����A���2wD��y��g��s�E����kW��\j��!��	�oP�/{Z/���ȯd���q�v�u�]���/�r1/����g����L�si<�����/�����\vmX����_��o��r/��2~��sx~��/�-#)mA�l�]�x���LL���//>�,<�v� ��O`hU7f�s���?���4F�g�J����5�ᵃ�꺫���+���	|���199^�6�/�s�M�������@����w=�Ȯ�x"���^��1@�=��L:7�� ��4�Q��p.ں�i���S�֡A��-7�k/FPj��W5��Uiz���p�t�y�0^�(HT�@D�J#%4(�~cIȁ 0[Q�x(kc���;�b*��%$N�-�/�Y��΄����)L�����$��4j�,*�����`��c�Í !d�J��0M99�2�� `����΀|�G�\�[�n���mH#o0�"�a��҉����x��)m�kHkІ�+���`hqI?gn�0�5���z��!T�E̎�c��a��T̆Bn꺿D=���ꢢi(��|bQ��O�O��qI���p�%��;���ITJ���SuhY+R��z����-Zs���BG<���B*Aog�3+����o�`���~��8�ɉ9]S�P��:����S6�������$��4�׬���0<���%�.����Q��|�x8�d<��x�h]���I��a��40=���㣘�YA�gÎ��?�����m0Z�s����<Ş�p ����w�+���:\����UN�����Ǳ���`2��/<[7�G���%�܌151��L�"R��YA&���1m��o=lێD"�r�dj��/,��l"M��^^&�jN�(�Х�\�Ճ}������#�xn�>,,�M��gŤ��&����\p�FD�(�y���9=�m��P/6nP�1_#:�U~���Fg�-�2����7P.�Q(,��wಋv�+�Sl����=���KC&�a9� ����ML��a�L�@��>����(��w f����DZ{61>��vaxu?��b���HA1��&3x��=XX� ޑ@ �A"D_g�09MTOg�P(~�rE�o��pt|�����B�����Hz� ���U�X?<��Ta�8������Q���2����"�P��c���� ��]����2��P"����7'H?K%��yzz;��L"�#����+�B����E��,abr�tQt�x8���.l���ߨ��Pw��0���4������2
�_t>�nR~Mz!����O�o���wu=%��cy14؍�֯AG,���<p 5���l���5z�X�I� J�{M;�Bcc8=6�ӣ9�|1Q�X���U���q�A�=�V���/�@o
����p�u�:{����0��v����<B���nXv\��%��x���1+���)sO��y��U�Ap@r�1��6J`����zV�q�l�QO��WX���UHόc�]H�0lͯ��L����׃˯���l�����Ǧ�P����]t�����scC�_z��J����ڪ*t�/�4<��6�l8B�׮[��
��=%�V*6�h�msho��0��ҩ-*n�}�kƳS��m�k�����=<��wQ���e�B�s�.�:��˩��1O�,�;Չ�n����^tu�ѓ�ç>�7xa�^-���	�H?�.�s7��z�fCC�Qt
�Ӗ<�B F3�G3hK�H�����mވ�D�ęcG�t򰘐m��;m����95a���:U!�����f�H[i���:�y�>�}�|A���cD��h���N��(��@�pW:5�4D���\޻JC,〟YU&��	�LV��A�;�y�V�҇އ�n�ytt�Uo�ʒb��+���_�?~c�SȤK��g2K�ǃx�}w�������w�����/��3�:+��zzq��nĥW^�T��k3���?}�>�Y����>��o�>���3x�ɧ���]�	�d�50Џ믻��p#�~��Q|������Ѫ��;o��/�gh x�_~�·�糯�����M9EFm�m�_�ӫ׈C��z��B5\�e#�鍸�����A�:�c��4[�8~]�����lU
u�I�/��������
Yqm���&X�I�R�'��q�}�\E�Q��a�p �VS#8|`�O*9�^6�J�:�p�0��H��\x9��U ���Ь���->y���gg�j�jh�יB��k�]�U�!�٣�+��]_��->:_R�d�H�R��������k@�a��b�*d#�4�OI޼>D�1��z�"�Lc��a���.��@��s��sC�O*���4�OQ�8LP�@�:ۋW].ʐ�׉SS�
a��!E�J%��P\G;Yc�bM�ذѨ_A_*�ޮ��R��Zu.�0=�����6�Bvc�A�ZՉd����Ï`��#��66mތM[�#��%��l�QA���G.Wҵ�DЛJ�� DwW�	~=n��p�^�/�5�,���3��Β�O[$�zV�i�s��J�$�ѝ�chu�!4ky��)p���S6��O�b|v�D;�މu����An%�l:��S�鑓�
�aӦMHu�D{��`߁�
�"�h��M*�m�|ay	�3jp�r��h�­�	�k��7\�����$�QL�-��16��N��TPY��6m���;���g�]� ���ɓ��oٲ��q4y��F�T����bj6���,�u�	=j�|���o5p�[n�@�h |����0�~��    IDAT�/�1�m��]�����v�=�eo+�To��R��wW!u# 3��|��eF^)�)��Յ4��?���R���9�j��BAds�ɑE<����+Hv&�}�H�����n�@%�Qt��zF��QA �z�62�]/��|Fn(��}1uV��j����X���(�����,�y�%LN.k��1�ϢE.�	�;���&��p0�)SS�Ng���\��t�)SoÇ��w�ƪ�nl�5!�� ����8�B��L���:�9����h�A����1����,�<J�Ä� k?���>�b%�K.��\2,*���˻�b����5C�$�d:@G!�[GW2���å�� ��ػ��;.؆���x�l~�p�ŒZR�e�"�f�b'N�`9M��q�[�G&��J��ZY!_�Y6���ѰGׁ��b�A��A(D.�ǩS�p��&�g��'�z�z��NIbM��h�{�q*c항��@R0�B�E��v���TIϨ(�5��_�ci�8�B^���~���~����
Q��t�� /@п֑�i�Cظyn��-���K����� �R� ���Yg,RǪD�~�{j�E2"B��=h�:Z.]5���L"m��CCk�&�mf1@y�Q7I���g�G[n�l�\�!�8c��z��1�omj�����'W0����sLց;��:SW"��A�Xw������;��@�j���"���g���/��498q�~Fu���f�:"6�=\љ0F� ��>,����Ɵ�}R�A$�r�#���C�(<�"hzV�"3�M���0@jڋ�R�$��� c���F��K���L</���2�y�X ��a����@��5�F.�R�D��>�!6`+{���*h��'��1�3�/aq~I�zL�E�Y�x������_5�IF4
 f��x���؏���c��<B�s��Q��q�.�{�{'�t��!ly0�/�����tx��W��{��M��T��v_�ڷ���ݨ�*B����k�g���hg<1���N�F��T�!��`�.8�)L.7����;�>�c'OU����w�~ӯ|���u�ݸ�����A����������w��#҉�T��h\o�D��M#��6=��%����Ӕ]g�� a[ظ����\}�H�Z�&K��]oT�-UQl�X)���{�V���� wڿ	frc�h�&*:��6ȌZո���q�K�V��b�:m`U���>d�ǰ���171���ÎT��1M��iB�\�(�e(h�)���ᚠ2) AmVX��%�kx�&5C�&ov�Z�S�X�z=�_t9����m��һ�EaG�ߺ�rr����,�l\�rR��룭��pW���vt��k(��J��I���e!��ǃ���s�J�Bn��9����8(�Ȁ$
SQzh�X�r͕x��o��ߍ��Y�
e��ܐ�Ӭ{��� Ű*Y�z ��򠳓� 6�bU�V� }����E�-fP�02��W��w��k�4�uG��Sa{���|j�E�XH��u�ѩ������9|�)(Ys���}_bazR	���tߵM�z�/50zf'Ʀe/���k�>�H�a3��X��QUB�[WW����J�Ь�Q)��҉�?�ۇ�?��<N����F�`͵�V˹�U���/`��&�Ǆ��R�����~�*��J����XZZ���شa���|�X�_ye/N�%��DJ�(�Y$�~w����L!�+v�6�8ufϿx��I{���Q�p��q�CB�?3��S�XZ(b�*�O�1��v��54@���brz��ڏ\�Q��F��F}\݅m[7 ��XY^Μ9���qN<� �ǚ�==�(���$:��L��q��}�Ɗ����Ӡ�Z/�Rq��-B>�a?ГJb��]Q�|V�6�.L�022��Oc9C?z?J6x��-l\Ӈ�ke-k�~_Yѻ�C��W�Z��bS��B��_bp�e���Aф�����"
�!��P(�R��K���{��DO��ִ��6(JeC�dN:��-r�2nE�K�ɢm���>7�46`sDKf�oD�ZUXؼi֭�Ҷ:ҙ򅌆�h"
��]���/�3g���}�狸�������|("��r�̲���C�e�������'���p�5�chh����E_=xL�=�o����O������	\�c#���=ur���f���#Ea%y�&?���Ť"!R�h����'��ɩiL�M�\ɣ�ʡ�/�[�|R�8�BU��"�)�E�@с�1C�9u���r�OΠ�z�mv�4*^s25&�g��7��1��M*��jp�>]+	����֜��J6#W�hЇjf+�'0�
��~�#ز6�}������+�~�idV��.s��$֭��o��\v)�y~>��@�PC(�)�>w�sa�g�!�H��@���h�ׄm�o��1�����8�z@Kj
�����������`me?��ݭ�@�X9�H�m�����#jn�������"x�Mb��4��ɍJ�*CO�ז�MC�~���]w��|׽H��K�����/�'�y���YVv(�)H>��Ss̥#u?v4�@$��&����M~S?���U~`�1�z�P #�bi|4\��9ixd�*P.�,�ݶ(f�A�����4Al����U�6�˩.�b/b�]���+�́��R��(}�

��EͤO��y�P,"_*��g �V@���G��[P�����Eh�+�`���p��oEgwƧ��k��x��gq��	Tk������ �_@8���;/�G~�Wq�e	k��5_��$A�i4J<qf�����O<��^��w��jo���{p���`x(��������#8��ޱM[X�a���}�����d�Y����=w���~�?IŤ��W�|�W���������ݶ�'X�:r2���zx(L1�pqֹA��^A"hc��a\�e8�0�a��s�`bi9�K�cH����gO�ɗNb�D�����!=A���`�⹁������a�ZC�n��N���v �C+�H�豁X�����8��Ә>y(�h���2t?�V>�
�!�� �cnI
7ZH�:M��n#�X4�C(�9&T�ƥ��Q�;J�<A�H�v\��;���F��G��@�1օ^+$G�S������d�Ñ����
WC kFZ\�.E~�_�KX�����(�͡��{�`Y��Jou�9�нsN'GD� D� )�$��#���l�l_L�/\e�G㱲,��� �� @"���sv�9u�ݻs���~� x᪩��*�sv������}�zV9+#Z��iLlbV|��_^�Df�h�L��!���>���QL&d�S�##Z�l9.�P@rT]Lv4$(�t�s���s����素�ÃF����(OR�j,؏�����b��̈́���&{�淊������	�]{��щ'�V�u�����`��n򰺸�,9r�@�Ë�pP:�6����z�T�"��4X\���`g7&��Z�N츪�@2=�gi��B�h�A����oB�8���̺BAB���C�������f�*�tyD�Ƀz�' E���2VW�ఙ�z��)t�}rm#�4~v�m��1LL���K�iJ�R���W����d� ��!��er�KUI�jSg����o���̀�l��+�l���]�s��15D��.�ccu�1�*&�u�#�F����Zh�p��p�XX��?�	
����uF��L�}�v�-��9E�1?���IR��<�X�����K(D�N�`h����]��������|�,�=�����y`�����S�:\z���i�U��r:P�g._��0����>�Gi���k��P��`����x��p��m����&966���~�ku"�$ֶO��Y��o�`7D������X�v��NJQUhg4"�-��g?�g].J��4��h�e[W���I�k� P���*��q68�k�l��J2�=N+N����|
�Yx`�`{g�RF�6�&�N�v�{�1�|���Ο:���1f.���������k�@ww?�����l�c/r���n��uɡ�f��$��+/����l�����)bl�_�D[P�T2���%�g(ݚ:5����l�l���eE�Ti��f��a�s*Q�q,�\��ͭmll�¹�ˍ��~�=3�F��\�,����34���u[���v�Z&��'w���!�p ���(T<9Z	����f^&X���xM�%m�	�Ev�9)���5vky LdSR(�-h�)$v�v�o�����QҩV������K/�X��a��:;��c#x��O����x��W�g��ć�vBg��'2���9��R2Ħ�L8�&z��Uv�+��s�Qz!��g
Ї��^) r��R0�<d��}�����9V%9�<O�ϲ 7%�L#���X�K����;x�E�qӐ�&h|�~N�����9� /6?���෿���lC������?�K1�r:��:��0�A���hP�l��$����g�5�I���`�YI%����g�f�΀6��4���
�f<V���U�$��\��3�b��fWi��PӖ���LdJ$�����{u+�^�M�5`!���_˰6���Ry�z1TU/9�i��P㟆��A��C�X���L�㣄LJ)���<�jU���?�4&�L���}���5i��O���I�R��3N:�&h Ԏ���Q|�����ĄH�9Qk���ǒi1�n�Ń{���؅�jD.y�\� =�~<���מ��Л�3[�V�X�71�s�_��n4���8���K�|��?�k�����s���o7��ɗ����?�ڭ��(Tf�]�H��u!ګI�t9NV�2v��R��a2���8����`w'�P|L[��8.�ɫft!U2��7��- Q2h,ߛ�7�w*?��
�t̌hTQ��$���&:�+b��0PR�e�F�F�t��,L�pyhD"ĉ�-
Y�I���4Ȃ*�UAj$��j�Ɇ��v&�R[, �O�!��W�</�h��"1b2n	(�k(&�ӏ���=�@xP��B�T��)�H4u�͗��A�6�^65v�՘T�z
sJ	���Nv%���%��L���"��S����W6�A� G��M����fA (����ރ�?��6��₣dQЄ��TL��L�zD���*�rJ�l/������P?tu:�SȔ�4�X�<���6�<.�;]�������9��)ܸ5/D!j�9���lww���W���5,�-Jx��@^�#�Zd�R8Z6�Xk�f2��+ֱ�v A<U���)���^#Ӧ%ۂ�O5�.��"7��q��:ۀX$���e�j9��~�~�2eU�%��w�� =�b2G�p�]�|�j�E��89��e��`� �V���#Qܹw_6܉�~��E��t�%	�I&�8If�J�L�P*�@��������`��0��l`?ǭ;+89�.�	���sEBb�G����@&I��*�V7����795?���H$c�A�wv��?����//"S(+]����hkwcx���<��P�j%�����E3o��w����4��0���Ϗã��wq�
��H�1q�F�跛dQ�!&UL�%�W%%<NL��;�B�RC����>��8��9�/걱u���C�JU��lZ�m:�t�^��"G<��_��ߗ5hhh ����j���ű����hWiu��@S+���'R!��&������N����9����pt\�����+�e��:eT�����4��H-�J�!b��@m��1�k��Y1>6"U�F�M}��.�t`]��N�L#��YoC�0�Ņ	,����bԈ1weq��ޖ5���abl�����������Y9�\�rA�O(A��_�>����|�ٽ8���a���d.�G�M���4�,aeeU��S���1;��W�ʄ��*������Ӟ�V�7���������OȞH���A���X�[[8<����f����z����D��W~�6^�v�f�S�����F�b\JCN�Cʸ�:��:/a�J.ЍfN�t�9X-�%<�W�+�Id������/����iS���o���\���_�I�����~�>�s/��Ͽ���O_��7���i>��4�kYpO�rrL��y<O�Z""R���	���:��~IA�W�Jq�z)�lu���[�4<�AS�g�"�����>����J,��ʦ�;���*:D�՜��� 0�`8�i�k�XYY^���G?����Ϣ�o{�������_�5�7:��D��!-� �h�ިe�7��i��}�,L,l8r�\�>	z6��(屵4�'�l`2P��D2�K����af��I�R�@� PCRy-Y��-̫�R-��M��t�&�j"��_�3~=�������&��'�NN0��R�1�p�!�+��()�sk
C+�o�j#�C�"��@��K$J�Hd��j5B�+#�"a/#�5��W�`��½}�))�z#�b���7#��Б�b�	h���dS{hSLx��G��c�A[G��r��zq?�����p�!�/�8�G6�-������>����]��J�����%C,���o~�[Ͽ��ԍ�>8�(�٤Ԇ�TZ0��)j��*�d>v���f7��&לt��Á�����pO7��;�ҕU�N�$�A��#Q1��?Y�K����`dѤ��'�����T��
<2�90ƲZ��#�:jתE1ji��'P8����<�V�ЈG��4��j�c/�Ui5�eq%bMO}�G���KI�l��h��}xģƓ�G�d����¹����j�h�8��j�05Hα!�� ��@k�3<�ޱ3v��3�(����d��u�AT�14��cJ�F������n�C��(����P�R���O� ����pT����mH�Nb���h�
Tf�����*��Z����{��U�s~O������;>a��H��**߇<rꦫ��{O�"D�F
.;�'�(dO����p� bY��-�5&<����^o���@'�{���
͸w�3o�\��ƞ���vt�hkgGڋT2����5�!���s�NWF&A6u$�Av�(Kku���@"Q���A��{2:�6]�S]�]��V=-����6�lʢ��2�R���>��XG�焇&=���F�#k�Q%R���e���S$�$�(��<t��݉�vv<�H��0r���8=Ot��;(]�|6#�k�l��0�8�c^@��LT�>��N��`_#�r��ݟ�V0=����(�Eދ8\Zt���#�D6S���6��pr�@������p{������ڲl�CC�u ���νi1 ��I銱k�n��h'\.;J�*��g�t������EѠ�|�͎S��zm��� <n��i��*T:�Zi��#�N�YfB�F�x�XH��R��6	���/�B�H</z]]��v{jvw�Ba��`����"��mCOwH~w��E����#��02:��+�zT6wP�ac�I���,�,r����"TE6)����,�۷���l��`��Q��Qa��bf3�5���t��>��5�M~�d��6�N��I&��������3$�]�d"��o����%Xh,�����嫗���Ij�ȉ4(�u�K����%�L�3*	J�N��ٳg�ibg�2�;���+~���R���ul��p��<��$�8��$���ù����k�p�ނL��>3����6���ݝ���UٹU	ӝ!Ν��X��N�'2;���Y�]�2)E'h���j��~���C$Ri�	ٟ�����p��)���T�r������9��bwAk$��!i8MU�7ʆZ�/�!���d-���Þ�cVP$�@�zI<�����������م�c$RW��K/�_��7���"����q|�K���="�?~�ۈga��`4X$����a    IDATZRu%O��Pn��Q��:J8���8j�WM�jʑH����R6�D2��Ha F�tZ�ܳ�A~S��½%�ly T��$V��"��r�(A���E�aD35�6
Z]t�bI8ZC�	0�`��k�0�,����	�N���@$����bq�U���	&L�SA�6�C&� ��DԚ��P�Y���1��	�,)�cs�QA�ߏ�P�T�ӷQ`A�#v�\��dm����Ţ�ϫ��2����hu��ڤITR2�֤�U8�k�żZ'������,����g�J5��q��ǂ��@+��F�H��S�������lw��lC:[	0�ETZp��kN�Z���S��d����R���OH镰�L�$��!Ĥ���
0<1%��,iK�u�O����'n4��&�O�B�*3Vb��(抰�m��B��z�Y�x��'>���>���(
�+�򙨖+�z�ڿ��3��׿���e�_��\P2��닏�uk�+��6wP�#�3v@s#V2��]���"�%nL��x���T���{0�����р�P�OM�iѣ·��"������x��s�����i\�q�VQ:���&~-��4��7��n��8�r�qk'��\�Sǈm�"������9S[W.����<���x�L���ӭy ,)��hn�u�`H^GR4�ݤ�E��)!���(��9�(�f0�a�[`��a'eH��I*�|����"���/�
e'`�"Ǆg�H:�CFy��İ�a�YEB`���)�5���ڸ�N�Z�����Ʀ��גG�R�$�p1G�Pݬ�9)h�	Z&�&|��� �8f¹�~ x��Hj��:� ��EV4����Hm�*a򢘾�[TF!����´ A�σޮ :N��w;
5�p��ֶ�sF��P_ �'z�2Tȥ�њ��5D�~�ά1�Sc8uz�p@�������^��^.��c�8{j>���2��0�c���������dCc�����$Y�X��d:�'e�t�f���w	��zvs^�I�����U�+7�qp,ґd�$)�q��b0���!zf�fF�Cr
�@��`6�pt����*:Bm�n��G�tEL�L�e��i,�HO��y�?smKK��j��h���x�h��"��bfn��.!��U��χё.x<6�0�2UA`.-��Q�?���S�1�`��޽��Q������D&W����`J)]��h`(�KF`4jE�ArN._���2L/�f`�3 �,�J��L���]�bY��9=mY=7���M�A��%RB��<��Yx�.��_R��VJ�#�	���Œ;;iܺ;��}�,t�u�������+ގ��Cܽ7��è�n��98Ї��Qx�N�R wqy�t&�N�QL��t�t���A��1_̉��0�83ӫX^�E�b���B�d�c2��́rD6�L���@�y�@'��Tt7�����J"�������l*���9D"��Y������gN��
{K��0��5��x�>�.-����(�2|x��et��Co�#�+�A�޽x���$ςE����8nޙ��ZZ��F��05ԁ�>?��F�U���ܻ7-��C_D� 3B����RЙ�n):�L/U���x��gE��:ꭷ�q��M�F|�ɇ04�#��\��%�[�D�h�XD�Aii�J��;wJ�&v���u|�_~,C��#>	�l6J�xyw��ti���VwW��2��P+_[�Z�0�א+�D�kF��)��w>c-��%�vu�tmue���o៿���X� ���|�._�s�}���wqp�B
�Y�l���S�Bo���$��dDSi�W�.� �� �aX�E��.#��)9���V͎u6���z��>�3��V!�2K�q�{�l���E� @���(s"��A�E��p�Iͽ��P&�=�5M`A��2I_l����8�ư���|�-�X(g6XP�jP*��@�I$�6 ��`��`q�P�^K���-�Qz�'�*�ג{�	��\ ���Ӹ���ى2Ǹ���8��������	��,n5e�M��`�i����R����ؒ+�+��O�����8�&etWh���L�O��xB��F����jB����fa�.i[�U Yij�*MG�
M�5#2���@��e�V��tV,V-\>����_����r��h2���e6�ʔ�Y�������fqbc@�$�F�
]�� ��OP��X���g��(Y�ڍ��6A�'�	9W����T�i7��ۿ�������/KA���Ǚx׾���-��o��� ��Z;�Ŋ~Ŕ�cTUd
d�V�^��B)C��:<��#x��K�d3�^^��j���Sҙ�R�+�ś-l�d��΋����k<���R(��^
�^#�d�"T���\n�t�H қi~�I�'�2�!���͹�[�A�hW$B&]�JFi��PR�S۬f١恁�o���z�H�OP�7V'SW�[d;B4�ԑL�p��/�!�X�4��Aъ�ll�ރ�(U�>�¤w����"쒙"Y����h��3w.>���F�Z�X�?L��ia6��#|d��%��.�*.t,��=Z��ʽ�(�)Y���E�QL��9�]��95i�H&��Y9'����F�K2!�?�U���=�>��Hh4X�݇�@i��YH��Іd� m��X�^�CM2hʫ���sL6�ӁP�z4��*z�lD���'�,�E�6�������e��Ƶiܼ3+��p #��ҥ65������NDR��^'��0>Jf��|=@2������.���[�h�{�G��)�ٸX`R�/��f�%D2��~���P�d�w����F��@g���*S�D����]��E��v�A�d/游7`�vU�GN�t��ЋB�mp8\r�&�5�ctr�<�شR�P�+Ι*���ܘ`����E����""��5%�xj�CC=0[U�s��>~��H�d��Չ�����ˢC����ܝ.4l��|���\.�pѯ]����	��066!�Ζ�"x0����Ⱥ����ȕI8]fE����<fVqf	�Z]�{�B��̞��l^�a�	'�idXUUϊ@XЧ3
�K� r��]����i�`5 �bC�Ca��v�N�ɋT�����N/`� �NAp��&�:�K� �?r"��H�X�	V�����uS����s88<���	Y�߇pWH>�j6!_����@�Nz{�`���ŝ;����u@o�#�m��b�<T�bAК�n��U���NL�<�p���&KeB�A��n��9-�ߢ^-"�K���9�����{[��%������c	<
�BB<���������3�X�9=)��T��x��ٙ<�?���A\�pJhO��7�w��7��/n�ǃ��0Ό�=j��	�o��ʏ�*_Doo/{�C�lg�.��q���r�7,�C��+�>�N_��sx��Y�oޘŽ�w���{/�3�G.]@�f���1��_�q�2+Lv��!T���i�
1�.���e'9#k�HN/C]��5X��M�U�ۚ��|ɖ?i�:[����f���Ke���+id�k{�?��琋��</�?��䑼��W��W"���p��E|�K�
c���s����w$!�	�0\M�M
�L�k�W�+��<��fA��D�R�F�<s��Jm�vLMM��#�J�����D�JQ�!R�������չ��y�[ ���ȕ�3��f�2� ��� ?�p	l���w(�p!vZ�N���asB��`scW.+uJRp�4ACR��f�hVS��w���ցB��t�����j��J���˺��%�N��LBbc3��Q�6?�r�\7��G;��4*��@_��ǭ�����T��]�U���P�U���-�?����De�����)�d��4���˯e�����K����R���� N��f�@>
��4n(K�Ǣ���V���T���4p8e�XFc�����u�:N��H��פ$�&J�,�|T5�vBa�I
/��l����H�Ȕ��� �l�LR�Iz8��k�J��=e�:�n�o�.���J�c����Ư��������Rw��b�����7��,_{�y�{]���&��(n5���U�-%5b"�NUN�	O}�I<���Ж��o�A9����qI��1L�� �	9�ѬϽ4���- Sw�d�ʁ�o޻���Pe�Xe<��n�mFǨ蘺ȉB.���װy�.��LFt$��<[�B��9q�2�a$�O�xt0�-H%�0M��C���]*�N��������!�旂���T6���UI�㡘A4�>c#cx��G�����ӷ���X��E�fG�F6�M~f>WF��z�a��ox��H��X�gp�41ͲA�''q �2C�(�"���LN�J�!��dC�PAls��s(���,#�%ٕ;N	�ΛW���N���(r�
��mN� �T��
�_�4`7��S���4N���A�U&&R�(�����TA+k��\_�|��%�z��L�� ��i��b�WV�NdB@�Y�f�uy��H ��ۉ�x��� ��{s������3��f�`���,�-�n�#�`l��9E�4�fH�	��G�PIL\��5�J>�]��֮�z�Lv�yy=Y�dԩ�5�<<�ΐ�m�È�]m��`���dp�bek;�8j:r��2i)d�����i�&�ɏJ9#�6�ǅr����%�-�
�}��$�=tv͸y9(��D����pphn���.�lbieSR�y�vXM���� l��5����?x��$zp��(�V��S���ū���ݽ(�/�8��gƄNA�0G�7n�����PBΝ9��.��~���+r�����ۉ+F���_�X�~,���}<�_F,���l�:	)Ԉ���@� &З��"��Ҽ2�P�s9�VS�j�Q���y�.���qj���S�mC2U��a�f��{ �Y��� .]��h��tQ(Yѓ�V�;II��\ʀ��{�����8����`g�P�=�ہ���T��ISG��[[�B3��̙s�z�������i�ǡ��`v��窮kɀ��H:�� '��~ago��[�C"]7}u?sc��%��٠�l���c�C�	u�^)I1������ya���L�:����d��M�Ш�y�����{R��V�+;b<$����qLM��u�98���f���E΂��h?���/`G�����%ܹ5/r%^��������ԍ3��N!���:dB�p��ĥsga��q���ebv�l�����u3n�\ǝ���Иff���,�2�
qY�8���*&�K
Z��
i7M=;�kZ���6�@"�h��n� Ǝ��Z���]`LZ�J�z%PN�`�Á?���"}����͟��I�s��~�#��W��u����/���������=Ї�|���˿�2����BuZ�by���� x~� O�#ͽ�Yhi�.�0;!�5M�4������#r�B�a��YeM�F��N��-�>�_S��*�o>��|)�̇�$��v��K���!��R��C�dT�13<Ou7��O�3��sf
{$���z�ܯ�6��d�d�Lɖ^�P�}A��av{$�9���D���-v�~��$��ب��OCW&�4����A>�ģ��s���K89܆����9��yhE�BI&����Y�<�wx��!�@�(s��~>-iZ�R$�BB^5u/�"9:��H�(���g�;$M�P����������	��1N�AS~��o���F��C�8��1�^��J*��K�Fy�������&�>6C��2�,^?�VN��a��E��4����
�"�"4����z�2�yʣ-�v֫y�9�t" �K&},��]+d��e+��~��_����3���(�m'=�{��?XX=����X��F�8"oR��>0� ����� a�|���Ȉ��ۭ&I~4jjx��y|�#���\�E�(��&�����;�$���n�FD��w_^ŋo, Y�f��X��&dU�� ���3j�2N���`�S�v��Q���F|sso����4��� �0٨D����Mi��?L�s{<M�K�UU���=�>���E�n�ı�����,ʮ"Z��,.�dJ�p<\�c'�f����������,��O���7�!�.ȡ���F�1el�4F�1r������+���a�@g�y��YdA ��F]�b6�Iu���)3�f'��g���7��77��Q3M�:SUȁ���EU�������*���4O��,Jy�<����SE�^������X��(%��擲�_U?K:8����l���@CmA������D#2�lI���}�j�e9D������A?B�@�\��zG̿zJOFz0:���D'��������`jb��������#�[��F��~R�/�P�0���������[ZC:W���@(��cϢ@4�5�?u͂��5�(�y�o7	���'(]���v"G��ĳbf&��׭�t�|n���]�EW؀���lH��z~a'��l|���yEOZ�瑌cmuQL�^���\���(�3�)����׶$ �{a�c9�?�B�Ӈ�H������G���プAYv+ҙ<��[��S��x�CS����ɕ�Rb��*677����d���XB�����(��q����lL�u"ɘ]ZÃ�ud�e��.��p��Tؿ$��MF����6_>H��*����+�/���z�[&T&������V"&��3�8}jn�Y��QQ;�X[߀V�Eo_;�zC�.QT���=<$!��`���ccr�)}>�ep����	�Պ��.��#IH�R���*n߾�D�.\��+�jv&��oO���]z+�6r�*$_+͵E���T֕w����N�ayL��(=5'/܌9M�1���:[,�:�x��+�ؼ ��*�X_]���"b�Q�^LL���ٳp{�R|��?�M%CVX؉���i�f����x���x����X^����:v���w���3x�ҨHV���p��}lmDe-u��t�,.=4	�C����L�v�2�7��^�( �`���O��æ�ݻ;X��A�S��n��c��/�r�gw�5�`�;��h�da �<9	1�Ƀ��hC�؀�`�É�h�*P���G��y1����1�3�q����.c2�*'�2T3hd������>�IT2G��_�)֖�ȣ������������?����>�0��̳����s��>����?��B��S�j��J6��3S��eo�c��R����Lz.�.Ŀ���Ȱ���?9�	%�V���s��"�ptY@���߷)�R�a5�c��2�R�����r�u
�J���e6�i}��V�"�IT�F��<���0"� �R�b&�[�Uv�M���{�R�E��ꆯ�%�N��\Q
�|�t�0�+%n�<��V;��(*��l����ӿ�!ԫ9�����ch�g��a�[������5%����L	sQ^������M�wZ	���g��f�Ψ�ୂ�U|��P�,�	AS/e�B��)�%���^ht����b��8.A���9=AX�~�N҈%�Ҩ�tu��ſA)�*0�B!i�nm� �w��HM"�Ĥ��f@���I��{q�Ԥ6Ve����f��j��H~n��U��=&��R9�P�I�rU&�����Y\�k0hn�Ac �*�S�]�ƹ��r��U��|?�§�����7)
�o�Y��/�����O�kz?�����F���
n��u�_T���ne����fW���Z&��߇>�8�LN	<�����Ϡ��@����fG>W���FIk�qx����HU��Y\��q@S����'��+Y� �*լ��f��T����m.b��[Hn/���L�$s�T��W���ެZ ���E`ww[:D���'p��9����pc�,!���)�4q��Ź����C;�H7�F�PW�H�fg��˯�ڵ�8؏HX���=!<�����׭RC��i,x��e�V�
    IDAT��/?���{�(�z�,>�E����8��߫"���$���Q�$����ý������$`vP:�`4j��V�H���M���\4¢�EP�Dm]uZ���+�����x�����E��VJ*�L��¹W�P��Y����P��cj�J��`��@��!�y�U�	��X�afq7n�H�����s�3��4�r�
^��[XXބ�bB�HΜ��㐢�>���Cl�n��qx���^�)�)��� �����S�F�BQk��sB��G]>5��X���!/ɪ�4d��7R�Ҁ��I.Όb�7 ��^�;{��;D"���e��̰L"#����n/���ɗ;NJ�����=�ND�.��v��H�a��?'�I!����ab|c���!W �Lo`~i�2��̂h���A��@6���̴��z���8���8��[�������\8���&�̨�d�u;;{(��2ε8���U��鱾z���M	�
�����Z��>w}���IllGp������k	�=J�t,�h�ePUM��8!(�w�(2��GF�p 8@ǿ�֫VRL�T�<F�:&~R�id��6��+S�����/6��ְ����*��y^��{��)�t�n��$Y��щ���N�`����hC8��Æ�n7�b����XY]����@�c����T6����n߾���=\�|�>�� I7����^dm��C�TCC��$�i�;6A-S��&~�heh2��d.5gƢcẠ&�����-f3�y0Ȥ���߁s�$�����ۍJ�p���R�6���c��B�ZB^�L�����R�̈�do�}����tįE@������I����&�Y���'p�t�\�[���V�ץ�nz$�ht�&���7��w����'��:fs1x\��StM6�ϯaog��cc��+b0�qp��o�ca�Z��	SM��-u�Q�n<��Vs$��̂�F�:~)M�V��]����Jb�.�1��YH�ٜ�X�6K�{�!�vNC�l��_��3HF�eB����wv��~�����3��~���7��ن_��3�·����?�%P7�l�i�.v����yI�g��N:'�ܧ4u�z�[����-��$J�̜�5�(ܣsY&�s-��in�؟��q8��Pm�!�d���M#��Z�V�S�Jp�FU�ԡ���9`�Mˬ��r�3P�}L#k]ܫ���Js�RX��#�q*rBɦ&�5*1���{`��vd+5ĳyjA9T�	����j�p��Rd�1���q�!��-��g?�I��ʋ?��?}ϟ�Ǟ�(6vvv���"�N����}�ȃ$�ѐ4m�����
}�-5-�4�̏�D���(�%� 5�2q���>��<T�at8T�*e��1��a� ��9X~t��$G v�b�a���g����C{���FƑJ�1==��u�*��G.�~�I/������٠�^G�kJ{�;���"�����ҜN�{��z�m��d�oIr7�TM��B��ϔV�
5��͢�ׅ���Ieh������g��?��խ_��໋�������ݭ��;=�'�|���:̨V���Ұ�pYU#�9�Q|�pg~�pVn�4�9�p��0��a8\حF��D�c�����AN�e���/��7��y��z���Ȗ?�5	bEH��o�C��P�1��#����*j�v�ag�6��BS�èeǊc>t���{�8e<&������l.v��~����'�4#.Jϙ-Fx\n�ص���Hw%#ЪE��21f�<`�S?733#ƥ��ff�E���މ��!؝6��A���I�P�.�����������|0y:��1����Ei��e:@������"7���*B��a��$�� }&�GY	U"��]	{Q����"�O�.��X(�_5#���,�^y�Wp��O"�m`/G���f
�lX�Q��C/AS|(T
nx���0Xc1 LA��@��r�:�ev�X݊��[�E��v;18Ѕ��0�:ݢ�7j���ӗ��<��s�w��.����܁�q;�Ql��gN�HA��W`��͕�LUa��eщD�{����\��X<���-,�1�"�+]+;2��	AC�������>դ ��G_W���"�����1)�5��ex]^<�Ky�f�C>���-0��;{G�d�^��qV].ޅJ^̪��	v@�b𤶳��v��P���"�a�|m+���M�s�<h��Po'.�GW���1v6�d���p{p��ȳ�����nJ�����p���:�)�!0h� _RYLY�6���P�9OgF�0�?{���.\<�s�{��T�cg?.~���"�\~NҘ�I�5ʪ˦���&� <�j��-�N7'kʠ�>� f�����:D����4r�����)��N��e	&K��]=�b�v�;^�u�/�.� ��%��kH$Ӣ���mw�����jT�8���
v��Y150��Pn������g����t2���6�l�����N��W�p�k0�\�5�%�\�T�5)l�T�9��@�:J��a24K! �|��`:+R��n��dB����8�b��P��0��ŹUI�&G��+�$uYc`�gE���<�)Յz�p:m�ܟY��7��U��cw[0<�g�����]�F� ���>\�r}.DYܙ���{���ȧS�h��}ｌ�	&��}��[XX� ��HP�*))��b��k+�����cd$$	�����O�bk7)�N%˚�j��Mj*��+F|�IjY�a�D�J�Sv�i�U�3R�R�IxFUo"�Pa1�t�9iU�<NX�)�5k�RY
2��2G;������������瘹uC�O�������cW����}��⏐L��ʣ��������_��9>+F�IR�'@C�C5��$5D�ǉ�'U�k9����I�⤄8L3+
I6W�L"���)��O�D�/������$�S�9��3h�y����0�_�����"%�(@	'�Ve>����J	�J�6�h`�W�
�I��4dH�1@gq@kr ����2b��3C�J�
n�.��6h-d��iDg!�B*[P
"P�;�:����,ʙ$���Fyt!4�����i<��e,.M�o��/��~��r�X[[�����G�[lu�e��>�)�uN�T\H��K�g�ł�I�jQ�Į.��J�V7�ʐ"M��.V���5����E��T̢��uz)8�5�\�:u�h
�h
�LA` lx�ؓ���X$m���� 	f��Jfd�?� �B\#��<JH�}(;eqAA͠����lh�0�X(��.�	���l�T
�<�4��~�$USh��h����f�ň*���A��"�J*V:Q9{z໿���/��_�����������k7�w>����7�{� �ۗ�d��F���Z���K�����
���V%A�ZA-�����1�O����z�|pY�0	b����Bp����*RU7t�L�-ՙ�V�pCfQP��T"�<f&��*���"[�]��Zb(��#V����V�$���F9L�R�a�������)z�=�}�{/�m.$�	�cW:¼��!O���Ȋ��th��e��+����5;x�q�dL�[oq2p$��t<�ӧ�
?z|(�=�f�7�dC�k��O��|_��+��t�- �����ŪB�4Fm��E��9�P�n+tf� ���W��Ƒ��Gvo��`,3�QˋBHRJ�#%sWכE�*��B�
��"�'M�hDI0(�`
���'����{�v����׶��(AaA�ng!�s��	>�W��lI������1:�%�DL���k��D�x�v����b/�:����
v����-��o������?zmmGR��:��ZD(CD�;;�`��rVyD6��J��-����m9�w�����/_�<�
|��N� `S2>j51�����>;e�,~�0iع�a��]����I1]E)�8���Vgg��z�A��A
���=�����B4V)]-N7G�f	¡.��9n�,���`h�W������Ww�eP�Q-��t�ҙq	m�%��N���R������E*[�YܹsK����g'a��Q"ݨ�����]�d�0��ij��p�2v�րD<��_����}<���q�ҘPe��h K�������m.���#%yɨ�KV�E���<D'���@ ��:�{�U=U7���w0�
UȂ@��}�C��@{���>tm^+��,*�(�=����]	yc�\w�ڼvx\1�%3|��?�<N\i�%�& {<nDq��[Hg2���v1C���u��+eb�Rv�I�gC+�L��R��AIc@�N��^:��r�}��Rr\TSC��[�!Upl/�f�|D�m5I ���B�ݝ835��6*U�sK2���L���Hˋ[��
F���)\�8�j1#��a:ID
���#�oB*�{Bpz��;(�7�aznV�GI�.��:0�B�\���o`anW.���+��o3`�(�������Gk���N<r�,F�0�E�P��ۋ�7��BQ�ݭ�15��:��;E���:����L�=���g�S����.^��=��`q��	C�Y��j2j6���PEСt�\U�mJ/�V֜Έ_C���K��\?[�bYc�{i�]t*���D�QD61������l����o�87-�7�Â������<+SȽ�m!F�u�KQ�ͯ=�o~�9F�H^
'g(���`��Ѧ��(�c��E�j#�R9��(W�"/b�D��Liw�#��mv��֩R��\:�t.+ZN�x��l)�E��ei25s�ҳ�6fi��/��v�����Af5�OI:bfK*���~[0,^��I�LR&l,4\�v�O�C[�����R09\�{�(q
]*Jދ�₁���Bz85�:Ӝ\�w����;��T�T M�Fh��orzb6k�g>�g��8L&�������^�gϞ����oݺ���m��FY����3OC�xj5)�ш���b�Tr
Y�����h��	`���*���M�5�o*�÷�h�b��},6;>��O����������q�<�@Y�X�Iם�kz&ut����w �T[�*8M�0U(S6$T+�\d���U�u$�Uk�˂���JQ�/Q�֔?6����ڬf���bq� B�
sQ�]0�R&�,�����K���5+�����]�xz�_��G������_�	����o���?|镟�nW�;�?��.���umE���F-IBF���Auf!�?�ۿ�ݹ�zrq#�VϪ�\������)�>QBE�.3lF�L��&��r*��f��_\ז����5{D��a�1��x�[�)j�U��Єh
Ѣ�����\d�3o�݀�܀��A%�D�z6���6㸹�R'(�+#�ʕ�Ǉ���?rUzG�QI�<8�9����s;]rCw��ho6x���C/1���[���S�&1f~���!��p�^O�H?�#����[�R����;���}F�Ͻ��~� ��:��6h�6a�k�F��HI�	J�y%���*�%ͯ��8^[G��R
Z#�P/*S�,zvKh|e�TbJ�?r@�y7����3��'�q�-�`�9����u\���LǱyp �_\�X0�`�j���jM��En��m���h,�mi�TL�����Sc��d��ູ�����*�����!�`h�v��\��{�g;��6���q���A/R�V7�<��L2'�d�M�����R�<f斱��-�`��W��I� ��"��B�o:]ƭ;��ߏK�/M�j�T�7r�d����b�I�ª�Iijt�~�,<�᰻ϰ���}��Č���@�H����E��$���삄Z1���jW��#��=�2E�X���:��lf=�V:;���a4YqtR���l��\��&�i�c���� 5�Q��:,67�&;���O?��҂L�Μm�ӤG�@a5{pp�5�<l��e��m�X�H�H�r⃠��ܙ�x���ʛ�&Wjh����[�V��`w�E�٨En�1�݁n&?[,Xߎ����eN!y�� `WQi�Q��f�(hQw\H�M��y� x�b�!��);��+{2Y����v��S���;rȠƛ�~��F� ����BowX%�k��=LOO�362���>�,fdry9<��!��bA&���0����H�[�����&re�j����H��>I9on�Lu���:��	�b�����W>����}��.�r�����`t�S�2rt,����Q�K�����	��\N���K��j�?�0���6��pȮ�Ղg�q���D�u}�oϊƟ��6�������ۘ�]��_��3�p8���?ĵ�K8��?)�4ϝ��hlNr�
�Ϭ���M�z1$��g47� ���1:��ޅ����It�t��ˉ��!Y%5���2U��|r+�6E��Z��$1�A�D3���;�U��L��v+(���Jk/��$�whI�Z�M�`�Ȃ�P���|<�Í%�|���p������/cei�*Se�R|���᳟�ut}�\�>���Ǘ���x�/�R��fq��')P/t^/���@�PC���-�ǒ�c%���B))��	�|N�T�ʪ9�?����B��N�]���ڞǱ�����=�$��e��7[��{��؆�뤃��TB*)u͚� 6�ZqU�zS�i��}�tz=�̽g���y%x���9u�4�F"��L�b�HeJ��%Y�Z�g����=3�x�g=���Y{�Y^[�d+Ӗ�I"���9�����+�{�[Mj���>2@�@}�y��>7(À��ް�����"���>�Cw�����]�[K�����0B�n9;qh����I_�t�d
ET�I��H�-▜i�%��Ev�Pg��l:�ٙ=���2�n�~�q|�����������}�oq��x�<��#�+s ��_��=�����j�C��hD[[)��c�&d��JFw�f@��8�D`m===j�ٔ�k�r@�Q��h(�xW��n'������!���ɟ����u8�����0T4�y8]ģݰ���3��@9c �����܋�����&Zn6Q�57 ҽXw��M*�1���S����a/�ͳ�m����Y �T�p:���E�� �����B&����6k����������~����+����W��/��dOO_���1���,�b$����|r����0����~~���~�c���5K%�i�����G0P��{,!���ڍ}f�aӆ��?�ƏN�"ߌ���Q�rY��@���c�ȁ��a�����$������[WP��
4�p{���Tء-+����� P����_"&b����|���7ɼr�._�(�y�:tHɡ\�QXu��u���!�s�^��'Q��H��)���b7���oL����gPT�ŅU���/�^�=]�����V1q��]HW�����8qa�fMG@I�\w�A�J�~��G�.ā��5�F��4�������^��*��*)���+�Pg,D�p7�Bt�C�Tu(�����j���u�����|��M�n�p{{.˥�����:}Лj�Llz�(��^��%	(�(��ɉQ�19:�e
-��L+lf�~E.��IG��e�(�S�X_I!����F,Ew��K���i��XҰB~�މЄ��)���e����X\�Do��hD��U�� ]�� ��
�g���.�Q�
�d��9�����ԋFE�̲5�%1�ׅɽcHp -�Q(��l[Jt����ښ�Kr|)���o<A<bCn���[�<u��|�iS��ͬ?��� ���� =�!�u~vV+eRz��r�@4֭��ͭ��؋�I��5�������p�A���~�h;76����8{���$����=Qwd��\��v�g����t(F�J!�����P��ԥ��    IDAT�".\��F�mO�!��R�p��N��x/��"�P4��߇6]��y�%����>�7�p�z�������n�Q�����@B�:��]��5_���	h=H7����x���0���"�t����,�]����I�=	�\���hWZ�N���������76>���<������`6�W�_�߿o����21�M���\����T^�\���5�?(�{img/^�Z*W�[�R6��BI��Dm
g$}��6$��m������-�ncz�B8~�(zb����`�h0ҳ����˗n ��*(��;����VtI�F�"ޟ�N^E�X��@�^��@O<~Ɔz�.u��.�XB6[U�Z<�+XODT����q����u���.�l"�S��r�V�{Y��ab�OM'�6צq���U�PW'�����㇆p`l6�O�R-�z00H�P���M�=?�KW�Q���%�E�l���:�6�bQ��P�,��~mI'��kͷJ������4���D)���	�R�=���4[o��A��C&���D��k@ju��ۿƭ��$���@����>����S�
f
5��ӧ_�_��gq��s�g�j��?�#[�9@51���ӯ^�F�Y0nx=!8�zx=k�eS(��p;�yD>�D)G�a�M9�0|��/�xw�xH��NjG��V��p�u"C<�M�ep 0�mY�*K��5Qg�N3��;TY��KW��q
Zmpz,�<�����p�-!�K���M�+���Ľ>���I�g�VS�ź�Ʊ�/!O��liR/�_(jʦ�4�-�u�v��g��:�*�Z�
gQ���N:$ϧ�߉�H��;�����u�z��n��FrE� 0�.��]2q��?Ӱ�ׇ[ѣ�F(̾G���:��c�<��ZjB�s���N�YI���ӫ�t��[itw�*M�ߛ!^��G���-
-���/��7�'Aq�Ep��>����S2��I��h@�ٱ�5��"����6�/���rڊ��6��xݰ3 ��b���\����׭j���<lt2�h�������j7�-�?�R�t�+���^D�T�%��-"�8�����~�����#����ۉ��w_�ݓg�}4�ɹ����3��r��j�;����so}�ņ�s( ���ƈ��(A>�����"�nk����X n� ��SV\Tx'I��5���
���� Z��d1�wqXmco]����
[ȯ�!�x($a�Kh�v��n�艛޴�p;=j��V�<ٿ��;��w>�ׅK������Z��cPR�|x#�^���������؁��~�����K�p Nוjx�W�rF�	��8�Ο��WO����Ao�~7: /���E\�v��O��}蛸���Ó7��mC�]B�~�Ssj���"y��j� �c)9ֈ�-�63�,. u�l�lV����a���S\��	���|���6�<�_��]�6P����y�)<��7!g�!�͊�D�r��/�B���ؒrD.)� ��Jt'��g�I�#��g���vV����ml�A@M�{��04@���
A��8��kH��R��\6�Ю�+)Ģ]x�{e��r�ĉ$�u���8}YN�����\w�=6�2�P�L�е���L��Z��m��l�X<���@���R���n����`&�	�(W�*�m!�����u�9m����QD�^=N�5�SM���a#��p<w���,�FI����z�܏ѱnafܪ���q��YT�y����	!J&(Ё��y!���iTh+�h*h�.8{G���A��Ѵv�D�I�KXXY�{�ky��c�^�R�v&�����ߞ��h˥4�JQ��{��&���ifLcn�&�8�#�� ��(��6��/\��&R��&�~����]�`l8:��X ^���ڦ(k�&7mD�88��@"��ݦ��
7�:�E�C�({���#�t�J�����R����좾�'�]wLbl�K�[��qkx����57��sh�t|o�b��ƍ��?����`/|�ׅJM6��bYu��rR�(��V���N�+�8sᒆg��#kD�	��^7�����9���Ǡ�M8�}�( �C�G^v�HP(�����B�s��eKG��h��aC<����7�Z9'�ǥ�^>u��,Bј�Rz{|x��{d{��2�n3�I���&pp�}GН��h�G����~�����8q��R55�>r��4+�ƾ=���f��@6_�����+�p��RQ�ۣ�1<tl{GGD�=w~�n�"����qƵ9d��/�����Q�Y�CWo�¦2�i]{�]�:r[G�]&g"���*"��d�ßلh�����lmwàJL-��͹뺢���E�JE؈�g����~�7V��/�=��\T�
C��N�t5�7?������p�t��E���N�:%k�;����<���142 ���8�?���*�Z8և��q���{��Z���2�����H�,"u{�lA9�x�ۅp,����OC�D4���i�1�v�q��9log:�u�Ă@��l���['|S��5���1PM&��^����SO=���_�<i�D�S���[��d�'��"��I�TZH���hkR�<��3y��I0���d_.MEΖ�\Hsd6C��A��C��f�k�Wݸ�h�_{�웟�G?�~�<_�.�/��g�x��������S�>���
��2��5�Ͱǃ�VRtY�����l�	<��F#бk&�N��i�܀�Ռ������+{ፔ(�|��x�;ގ������(�����_����m��A�҄V��-���]0i��9U=j��J���zE�0Jcv0@���4��yP��
��N0�du�ef�D6��>�'�����A��:�c2���Z>B�(�A�h���L!�\m$���?��w����ѷ�z�����տ:���ݟ��������~_0���^��P�Յ��ho�y�3x�[ߊ��<ʥF{�34�[b~��A���YY@F���"���6��j�M�n46rm|�{W��Ssȷ�+b<��v8I͇�^v!GN���R�b���毢���yX�,*�-�]o:/��^x=Ax��b3�z��F������W��.������ܹӸ>u�}�Eww�^ ���B�7����`�_�V�D�U�hH������իZ�ix�<��x7���pkj���?��Y5j��l�(�V�ڠ���=�$���u�����ZB�ݥ<��(T��:�$�2�:�����gs�wB1����-dgo�4��'h#�iӋP�5�����ɼ4S�[��p��K��Z�jjM����	<��gPt:���%j���Bn�\��\�́&��d�H�Մ�n���X+��;��{F����P��v*-n;�L���\�� �ph�]�t����+��p�ޯ�(!��]kqa�J[[fM0/� 	��:y���XD�����h7Q,1�����&p�=��XH��{����I��N~���r���N�6E�iS̀02���016��_"��o&Ӣ���Cg��^L�	]��ɛB���������v�K���*�\���r~ G�2��E��Kl��Q��\A���P\K�\݆��\�2�d�M�.?��
�a�L���䰐5�p!�����<���P,�g���{]	�~Ձ|���[K8u���Q(�ĩ����kҨ������w߁@4�r��d&���.�Q���D�;(�Â�$/,mjېɖ��e���p/&�a��K�Ϭ��fM�0��6�
��"Q�<�MLGk+WsИ3��sT��)z�|x��1�X�*ĭT�a�����2f����w�ȁq�����VW�nh����`?�;&��k��k׮��;44�=�#���_"E͉��$�g�4X����O���E�C���\�����*����,��x=��l���a���(A�]-E�&��&�Z��RgF�grb}�~���\˫�������sX^I*o��s��6-�����Ǿ�.�v�)!R���s7q��e�*5x��(9ǎ����	Y^�v���D&߀�t"r�ر}���xS��6�?�M���2^�x�iz��Ն�����D?17��6SILݜ�����̰�zƼ��}�=pH|����8��}�^���~PGK��ӧ/�,Lgk�хb]�����o�>L:�H����5�t��u6D�e��GOY�h[�7�͗��\ǎS����ȟ��}�@�Mn��Gi'���^|�����<���/b��%8��/�@_[����!��η�矇?D;�Y�ɟ�	~�������?�>��_���Q��n�Z�����g�.�A��o\9�pH��bn����]j�m��`�5�T,�dO��:�Gy;I����P�?�0ڰv{s��k�JPH�&�,�x�S�L�A�����Q�t�����=�U�E�Y�a��c���G�'#�/_�j��m��!��.4�����t#۰�n��nwJT�PZ�6ɴ���G�ڒ�5tol�2�<j|�D�#틉��D���t�6�Q��7=�$>�������ʑK�ۋK���?���T?X�
�|����@�S��}�����\��w��x4���th2!��\��	��>��-���\��Z{�!��B.'-��������'?�w?�<X�����������7EO�f��zZ�2�M��S:!�d3�yM��h�2�/��75[.[�R᠖�XLS�
 ԕ@��B��_�h�n Q�>ޓJ.�6�Zj��/t,�5P��-3��3�nn\<H���khW����﻿�k��O��{���&��������7������@0��L$�?��֜��pW��g��'��۟|�z�s�_\���&�Gp��a�u��Z;#���z��XX\Ǟ=c���?���(�U�w]�RT��@��.e�����ʋY~�mx�6��<R~oa��e���^����V9P��K*Y�[y
����^*��Z��h?���7�]Ͽ{���t��[��IhP�8��2׋\I���,��~m@�"�jŗ��DpY r��Iѫ�hc`hccc��@ţ	�ܚ����7���¼�
l@�^�������4��w?|/�V*�·N��g�a����MN���E�T�aw����đʲ����ԗ��6���;s0��!����1��ա!���S��2�����������X�������oG+��JjC�aD��
x��o��ͯ��dK��v��.8h2�Hģrja�o�Q�����P�\���RPdY������~L��cRu�v��Ҿ�nT�%%�nl$e�7<8"�(����ؠ�)lm�!vhg"l��r%��D��H ��N�̙��Je	3�,&t����äu�N��6��Riz���CW<��Z�Q,ױ��.�I����p7��5a=�X������ȭGE:B�7 t}'�|�".\�!k־ބ��D����f�3���P.�������˘����Ӌ��=7��d�����w�]G'	�P��D�)�m��1���i-80��ѻ@vO>[�փn_3k8u�2R&�a&~R�W���n���{�����
6w�q��i�����O`�Đ�*��PJ&�
e�������]�����@�V�m|�(�73�xe�Ԏjt!/U�v6]~C�ik � K.2��N/�K��6�{BxӓiPͥ�u��Mk�n-�)C����"%l@��?e�5��|^sn�Ƨփ����k�%�<t��z��c�kۆZӆ��g�깋������탃	Nw;������]���ƫ�a5Y�7�v�RW�E�|)6�y��)�d6`�-D��%&Ո��ha�� &'��u��3��&c ���v3s���Y֦�nN2ܾ�t��<��1���fn��{y��2^=Y��dDp`��;*�Kn�+��}4��s ��7V{z��V��}�(?�����X�d _\�U.���Pw݋����S]o)���kHgKJ&hsםq�~�cy9���^���SBF�x�A<����������n�7��G�f6P�z	��_6������m�� /�x3s˰��p�ʭ'���-V�"�1�P:5�u~)�6μ�fKN
z�b~��B��M���|�]<�/��H�^��IAk)����P��:�_��G��U�ş�ٟ��?�#!|��ǯ~���~��k�26�r���	/~�%Tm����vp�J����KX-��$����P�g���D���l�#��H�v�{��rH��n����0uc��9�&QS�|n
����b�/�лH����(<�����٨�I�^���>�F��^n��dm���k�1���b���
���|�י�K�%iA6�M5��;B�I�蔛S����Ԩ��a(�5�<S��|k��crRx�r`A9�GhC��c� �w�-�Z��~�3�5�I�H%�3���T��D��h�X$�I{�.^�$@����PD�����M��O���_��t#�B�p���{��f�.�S�}7������m�|b�.��vL/��_�&~��SXZ�D�}˭?�	k��Zٸ0��h�`��M�=.�!�w�V��#
�V����:+D�����9Q�h=����8�N�ϫr�l���%��u�y�#���C5��)�7�46�Q¤3W�p�K�{z��[{��|��~94�|}�������ϗ�_���s���Ð�A�B9��c-�ް�>� ~��?�W�^����/�;2��{�|�7�����O����>�����������E���� ��5|���8yqC���=�i�t 
}5�ٍs�,N�9�=��(��}��먬ހ��Gu�▬_[�찹�j@�~��U
"����{�������O`gg?��06>���Gt6n�|N8-��3������Ŀ+��^�^ �TQ���lY8%����!�����ҩ4���q��9|���b.J���O�'�A�$�Q�\���N�s�x	k�.�{���օ7��N�p�!:T�+�9��:��!x�v�N/`��Z+K@qG�͢����5�֘�M9-[9�Q�-� �/�u$OOA3t$!oN�̎�!ҷ�����|V<�ō5����+\RČ�`�1a �ܸ!��(�#�1;-��=T���
��F�������<D1�~P��`h�mn(l�l�ȑ���R��O�6�� J��g�nd�FjQ�Z͎<�|���l�K�*z���g|X�f~n�+�2�pr �������^bA�1ͻ�&�⽠�'���~kb}3%�W�}]���&%&�!pq뎭�,�;;�Ts(FcHm�p��nͮ�VnH((B_�ī�A��)�u:k���@*����T2'�aҭ�m��j������8��<�yn��ҷf�1?�l�e{�q�Gd2���B�L{6kIܘ_B�L�W<����k�qdr?x�.���L�.gs�t�2�o,���w�}�N� A��I�W߬��'��沐)��āz����&�N�B�ڔ�;�	��ٴ�������19`;i���6Y�\�Ku�����D̃g�z�J��D�k�SXg@��2�9���`=�߅��9����q
�(kv7�����Ü��H8,������Lm�_J������_D>W���E7�٤\u�q��~�\7D�:{�f���D�X�p'���*�k��.��	�i8���9!{F�!��L'ക��9��r�)s�BJG�L�J�\I��멌�ݑ�c8zpng�4;f���p���^���������q��*^���r��e�h��`�������`����N.�l.�ͭ"V6Iwh#��"�����0��1�B��������qk�$l�`dϸ�����P��\�0���f��=��]xӳ�Kߔ��P�83�����dJ�,�v}ttPg����> [�Sy|�;�E:O�"�' ԕT<T��N���_�!|�#�7���t��U�P+6�-_�9[u���H_�:?�.�P    IDAT�~�#�76ej�ڴQ�U���ˢ;�#�<�g��D��_��N��7��c�>�}�=��Σ��R$ˀ��|�+���� W�����"9�y�lΫ%X�"��n����@,��XK�Bf֐��?�-1�E��?��t)}�v�?��+�|���!|���[&g��iOO=�1L�&ȗLn��3N�&߽ 7�?{�(b���a��^�{�|�ZI&����5,�na5U��V�%�[z��E`s�d+J��~���-�<�e��U)�Z,�U��Pŀl���{�8��'PoYE%���k�{�������@?��cʃz�嗱���A������ ����+!��\٫���3�"��C�B�����ζ�����{ �9�ŵ9d��s�m����0�N�����{	�T����Q��M�������~.��Z�K�� ��'~_�v�rڌ����M� '��~��sΨ�`��1����w%��Q�9˞�Xg����v����&��,�쌈��hol���S�e��q��l�A���;4�����ǟ8���Oz�+�Ք��~��O?��?z�ܕ\ސ�VZ�@�~0�]����COЋ���>�� *@տ�J���o}��x�0�������A_���p��p��x��''�w| --Q������' �/n��������(��
6�Ä�-�_�QQ�Z*b�L
��%dWn������7����{M7�+�B@�@�Y�K=D_c�x��o��� nޜ�ɓ/��s�G�r�of�r��-��CDkWX���O���k�1�#��ѿ�_��X?_�~�J��J�"�J�TË/��s�"_��f���O��h�9'�����?��|��QĆ���l"_k��l�ؐ�J�9�"����F��s+ظ1���2��-�*+��V��N�!g�#t�Φ�H%1��i�q���y�f�4}7���A�P w��a<���camղ��w�]hR��N�b���t jp�3��۩5;?!��Y�YX+�l�x��/�W �Qiuh����9)��=�Ji�AW�0���G��N�99����۝ύ��#6�M��ɳ�|n���ķ��Owcmø�8HW�n�m/y�y�$���T�X��m�����T�O�K_�RB|n;"A����GW��Z`}3�`�I�Do�n�w�PfwL��{���A�E8O�9mE�����N��n�l��8��*s�k7@,va�hFG�b�U�-�a3�#q&��:��#�\,�P��!���,R�Z��PKK�fn{�\ݱ &�C�p/�^���u����tQ�؃���`�ǏZHn$�2��	:���ΡTm!Shcfvs�B�v��T���f�%����5��g���/��yy�7Pi	���7܏��4f "^���6ֶ0���,��x��.�w�9a�B\���Ϲ\�$��cBї�VD%��E_O����ו�5�6s+��O�U��'t�Ir��8zd{����iy���
N�� ���I��W������U����ԁ�Y�W�Dw��Z\`�/�Ѿ(|�|�:~���z�&��e�ݩՑک��Ԝt&L�C���@r �-be}S�}���XDMb�X���4�M-cn!�'�:T-��t�1����H\I$�@�ʤ94P(���,c3��Q.�16ڇ����� ����k?��|Y����<^�~�����H%�8�A{fA�Ñ�{��wb�/�v��3l�%��L)l%71�w ��A$����b6]h�C+vB[mz������������^�~q P#$Ӹ�N�"U��tQa��6\6x)O��U�A�e���V��$%�D�}��5����б����8{�6Rk�;m:S�{�q����'h�������X�)#W���ۣz�-@){��������E^x������ɟ�~=;pW�y=礪�]N�/�!�������'����z�!b�������8�������	�	�\gϞũ������-���	��|�'q �=����VV��h8B���f�qaj	s�i���Pk�`�D��Ѧp��[u9�1혯+���ʨ�*�*��l�tg�Mܜ��$�M1�N���`�z�(=[,D"���BKE��V�Q�0ŭ��	g�Z��Β�yRd:[�g����3̲�\)/�^_o�1���q7�(^�p8�^h��TAn��K�����{�g���<nL�Ȍc+�G����P H@0uY�fLf�AӃ]g8�ln8@���;$X"�إW�5��Q��>?�pm�Dj+J}���Ѱ��.�(X�"���V:g�t� (�Nֈ慓�W'��t36Ԭ�Ԩ��@��Z~�v߱����������_����n���/|�o-��c��d`��/��Zi�Ǉ�Y�#��ޣ��wcs��p���#n��Μ�o����X�����z�.����<��#����p����i� �ZХd_��Y���*��n8�	�0��B����b� 	&ZLgm���+�H�L���r+l��m��2��Ku2vs��f1?�ч�Ǒ�	8�L����'���k�q��K����x"/&Zh��vP\���*��(�]z������HS_���T��y�'�I5���I��H��f��r�h<y�Q\�>����{�ɦ�q���p� �==�)�-�_�G���M�M<��}�"�/#S��4W��K�G��`$�&���/>��W7�5;���2��-�m�Z���&���6=��QR�)�����2�0q]�F���rb0�	�Pg�ឧÓ�y;	��꒸�D�����kȤ���7 �NY�����e&]r�jԘ�Lv���:$���*�3��5�mU��&Փ��27Pe�!��i�h�}�+�+B����f����B�m��h��fɤ7�Yc�E�^C�0(L�"B���{��w2��K*�����s�"b��˴a�
�;�؝�)>�a]�f�J����I�Z*k������N�|m��R�����l^x�bQ���N_k�ܓ2���%�{/+�O�t�X[W"�%���VY��@~���ִUQH�eC$D�}��Hܶ(`��@��NrD�����?��3���>��w#�P.`c}���L^V�]]a�yd��p���mm�=	��.�U���!��"��bqy�TҸ�9��QP��]~��zw S�C��C�`[ݴʅJ�z.w����c���u%_�b�v�k�_e-`C��_"��`o�6W<p�g�`�;@ʗ������"������ � ��RS�76��-�<������{�g�^0ɕ����^�����L��L�zG�ʍ�|� m:�d�!1���u�h%���WNS�X���k����-T+�a�h��F�	:_z�R��05���W��;�G|~��B0��V����Ts���(�������XZނ�lؙ��B$�ơ�Q%io%ױ���p,��#����2�V2��Ӯbh0��;�����Ŭ���V)�-V��GW'�~+�*��(�׷e��͕�pǢA��q��^nx膢���d��P*d�z�?��&7Wlcfq	/�zk�����YM^$nI��A�U+L���^@�䡓�{�瘎F��t�0��(�שp��D��[W�\Y@3�S" ���ZNju{meh}#[IwЍ�l�>��;�	���[�/�L��KI̯�1�̠��A�%�	�c�!�Q�P,���~7Z]
S������.T[����%`ǆSvʤ���X[��O^:���$R[e%�a�888�'�x��{16ҫ��g7��O��������kS=�ΒU�-��t����)���b1��w�_Amd@\���W�^���6R��V N?7~��qC@�n�^4�#��X.)GÀ�&Ԋ��ͧ��x���W ��B�\@�L�h�AQ4s�8��>F�s�r�KL屔�:�Xw	n�� ݔ���q���S_@=j$y��O���h��۲�m�ͽ�����{�s�����uN.��,����$���A�Dp�l	���8f��+�~��-cC�m���͊��#~?n�M�Bj?�՘���b+�G���9�"���S�РYs����F)���Ђ_�
Y;�?6Nf`� ��ِ���/��6-�
ET2��C���o|�O�_���O_��W���5Xo׻��g�K�#U	:)<��S+�=$�E�O��L|:���O�~���r�ȇ>�'yS�oaui�Lbt0{�U�D;�h;�Yv���/�<~zzt���2�l@-�%�DN����*��א���Vf	�m�MXm���̖��' G#>� ��x�s����8vҫ�3>"����D��M]�׾�Uy�9���;1�a��������ߟ(FMr'��}�eH�c�U*�c����N�}}��Ў�bjH-��7�
�a�����(,�c
���pvs6���/?�o�'�5B�s�m;�ng�HWj���E[�5�ǡu'����J��mV�к��Zf6aw��p�Ԩ��Lb&m�F˳zYu�8u0�e��v��@ECA0m4�.�=���7��?�fЇ��E�km]gڟq+�3D�h1���A�P� �P���
��z5i 5�4�D�,"W�7u�(oVԼl'R�;ऋQ3��L�r�0vkL�&�����!�=!!��@���^�;L��u��7�PI��������Xx�/�ntDO���x������Y`��	#� [6knԊt/�y^t<�Ӽfk�B��b��Yr��,,�m-x�Ɖ�F��dRAd3h�/�b��1;E]����I)����
lV���j�x ���j�!���7:�4��*��pR�h)�k���.^�L��h��9��rsXmT�`F�hT((��I������R~��	$m�jHe��U���o��g�a"����^�,��?@���il`�3gǕ'[$Ռs�]�t�^�5�M��t	�2��|��۸uh��q�Н�I���8^�
��
E,.�J�GKaZ?�U�@!���t���9��g��0R�:����׭!����R	3���d��8�#��46����wŨS�� ��z��f�)�}4�qYmD��7.�N4h l�j��d���^9berUl�1���7gQ�T0�Ӆ�xD�!��EC�̌�G5�)�Rm`}-�3� �� ��{�G����@G3�!��X\Z���w�aye7o-K�K�[6<3Ba�R��"��J�&��Z_�6`��c�#�S��joI�ᯧ�U����	�Æ�ϩ�� 7w1�D�1Zs��/���o~�P���,.ߘ���m��L5i��wM�(Չ7��-{�1)�ry3����x=�X���T����DnZ�
An��X�v	s���/NnS�dicy�Y�Y��J7`sS�܂3��k��12:��DP�(u�z=���w�+���:���u�`�I�mV��0��`�w��z6��!��DTr�piyl��E�k�PN�Oבc��^>qFt=f�x`�!2}��A|���3oz� �qF�ŕ-����>�������@( F`��Rt�����YR������?D_����n��秮azn�\[��nf,9�ږ)j�Q���&��5��� ��9�4�S�M�#Kpi��S�)q��B�ZJ��'�8c*ěgX�[���5
�,��JTB�͎���Iu�؋s3���@q�<P���6z@1wx��}���P:�W��������69�8q��/`C�n#������G�7�u{F��j�ag�Hg
�����c�����6C�J%̜7�c��GgY�X����v���r���I&��E��Yd��h�+^v�5��$UAz�I{�7��a�w�������+���/|��G-����W��_M�ι��������~�W�w��n�o�^�ỳʜ%�;�x���]^v��t��o��G�_������~O=�4nL�b��6NNb�;[���@��U��߹���ZD��M�V�+���_n���e��ن�U����M�G+�4v�ZR��@&I�;r��FF�����h?y�>L�F��#[C��BA�|��������:no�i���C18:�r�,J׊���6��BO�KBTL�4��|�on`ff���G#r�����Ӳ�V�b>؁W�| �+'\4�,.n�o?�u|�K�Az�Gl��߈�G�V��T���ݍ��|`U
�k�E䆺6���D���$��MԶn��(���3���ǀ�z����(p�Yxz:I	�ߓNmrR���łU�6`�r�q��O�M�{���Kj���*$�ݮ��:t8���jX�x�4J~
�ZfJo�a�:a��zE���T�wRW):֦�n8���w 
�$&b��v��Y*�B�<Gn�ZlX��_ϯ1V��Y� �˦IJT�,�\%����n�D���i�P��q�s�p�<�mt�J��˫À�{�R�B��1"͖�x�~"k~Q��BA��D�ZE��EU���ϯ?�AhDZ,�lɝwj-��dLׇ��||�E찷̪���(7Eh�ժ6JmiF*rKQ��2�U�&Y|�����d3p���U�X�א����9�M蹩7�`��磍6�U�Ɖɢ
b���B�I+MRY�;F�BX[Ru2.#v}f�C3�Q�F6\^xv�5�+n	��:A�tk7��V��&��IT,Qd���EUj�$(G#���k[���g2�|�����E�g���68�"��=B���m�'��"ڤ�x��0Pò�X*#S�+���ݯx�����g���>_r�0����lH���)��C� 72lH����E_ODw���9%�,�+�ftd�bA�ӵ�4�r�g�Ъ6v��w:���qە	����i�8ئ6�)�{�G��`����{G0������Ï�+N��˳�zm�2�E]�=��0�߭3�i��'��z��L+�:�-c'K�Y~L�|��1u�T���,lm�ò�q��9=�Px�.�B��ظ�?���+k�q��y�n�����%��ѥ��m�I�@��n�#�Ƥ��>t�a:b��|�)&	�`��
8�5�x��Ν�;��Ӏ��7�1�m��`  ����S��q�ȱ�8txJ�4�\:���)T
ED���=�,\�\]X����W/WЮVp�1��a�`�LsE�^���U�M}n���qQg]f�m8���VB<]�fn-�qS�N
A$����}�}����0عn++I���~���3��,SK��r�Y��J��ݥA���
��Ό%�ު#�#�7�`�S�p��"6�*h�T9����J�(�kT`�Ƴ��@@���&6��"\kw[�K��x��1�e.�Z� z7��|F��`4�Dw���*�T8�*W�j-Ke�:f[��,tB֜���'f�o��tHst�	x1\Qr+�\���_˚Đ9�6�����i��H�����nMϨO(�j:�<W�uB�.�N�S[{��U�F[���Z���?\.c-4k��94���n4}n�A�xF�W��@A�E�#Чs#���B՝�(��A��5���P�v�&)I��<�t�&��I�|��W�#���/e�'.�|�o����|�g<L��p���8����jՄ�G���n�B�mo;_�7���?�c����C��qu���i$p�V�*��:���\������������R#���:Ƥ`6z��rp�ۤB��]Ϣ�8�����,�4PM�Ɣe��J��zʂ/�������h&XN�+@"���ذ�9ZԘ��B�V��3����-{������w��p�\&��Ԗ�2�A��.ٌ���t��/vv~���oZ�q���׃�?���, B�Y(,�q�^G,�%���SW���w��]�71�����0z�>4=>��
�9ikW����r�hK(JS"���ml/o������;��rp8���e�UF��`%6Z�]�+1�D��v�In��ņ���@�oN�    IDATR�u\�����O����U��V�^��X�a�6C��΀ m��5:v��\c���47h�b
��vJ�m��,�?iPoٴyb�Cx��q͆��(A6�w]�,�a�,0��D:X4i5� �&'jU����f��@���RY�H�O��]h6�,~-	vW��E�r�,Sϻ�&�M��	�H�`�%�+�6�w�:Xi�tآUi�	.�W�|�=����A�)Ho6��v������q��z�Ɔ���_�o3)Sl}y��_�kb��af�6��č2�hK4�b�(zj� ��ф4p���U� ��\�;N�����ψ~�lN��+�h�b[K���7��9�0>��$��g6E�I�5��y�8-�I�$����8#��jD���2[Z���9��1��ְ#_����`�*]��6�k~��j�"��y����J���߯AA�.^�z�r�FQ�:��k[B~���/��CJ�.��&�6��6\�rx�@/ݐ�@��L�(��,j`0��Kg�B'�f�Ϻ�h��,"n��+W�re�}�AN�0W��2G���I�i�Yu�ٲc��F	M[	� i	�*^W�[��H��ȃ�r��kܠJ٬��^ZT�]B\�Ɔ�����i�}f��*e��Dġ�TEh�=�FW�p@�n�]���3�Ц6H���a�͵����ŜU*EZϖ06�/KUr���5_*cyeM��`0�B����-QR}�(jM��tt9"4BJ�?��[t|k�Ɓ��4�Kb�=B"S?w������^�J��x �w!����ԙ�@>/�e��h���.p�X��y��Y��|	tE��±{���� f����+/!���&�{	������p�GaE�J_�Vr�Cɀў�����u�^-��M	�%�,�I{G�x���n��G�lD�NRR"qm����(t�����E+8��4Eܿ���xX�#�(u��yQ����e���Е� !�;�@w"����d��>o��eYX.�Q��r���2.^���z嚅Z�^�BżhUT���0�̨)����;�x��kYq��ɦwMzM��Z	�JNR>I����ހɭ��p�Qk��=_(�J��f�<9 Q3�k�� YI��@�10YC�� �`.Z咝`��8|�Yb�	�n�
#t!�Q+���>,����ի�5=��	5n�&ưg�z�����2����|�-��Ѩ�����9�,�bs#���pL�'�I!�K�������I!��+}K��\�Z�rkM+�LN4qY�����@�{���I}g�䃽2|���r���C���'?�§?�˲!���_��/��_ͯ�?�?8lѕ���۱/�zȡ�+���cx��C��B�[Z���*��l�~z�,��?�S��?��O��c���)�5;t�]A��"4;�O�����VK�KgVQi�����s%�̓�֌D�y�y��'GGyե)l/]E)���@cۼ`z�8���n���HK����(�M��݇���#�:�m�%똎�sy�ng��J [�cemU4��|@Hav+�l6��%c,���(F��L�YJ�_1��٣Mە���r8�������G��*d%�Nb;��\� �Q(����:C�pq���?­���6Z�.Dz&1|�.��F���A�I'��u;�,n�ӹ��i�Ë+(������vnNg��[;�&�R�J����+�5��e'�������@@��r:�4�_��Yi��v��7�Q��ߍ�n$���(��Η�����w�9;�������p��i�,6�l�L,<z����T��9lwH�����P�<'0��;�|��L�RV�����F�5n*�>��#��a�T"ϝ�ݳ�Z�mZP� 0a)v��4��#����y����s��i
���KFg��aT������)%�2���69��Lm�W��;3��C���c܍Z���^��\�:\(�gl�+Q��ܶ���v��0�9D�% o�X��ckɖ�{.r�98)U8r�^�wD�uNK�q	��y�F�+or0�t""����Cz�^��8n$v7�&
Ղ]�L9�^8�GVj@sD"9ᯅ������n�L�5�	>����Qd�U}�X�h�D�Q���jǃ�8z�i����i�E����Aت1���F����6�L(U�h�׀8�k�v�DU"tD��.�Lf������!��T�����i.h��-�L���b#O��ZGp'���B��wJ�rMJ����RQXg#��;ͦ�N�\A����I^�C�W|>�D��"l�ꨁH?��冻懣�N�[�
�<l�<��d��MA���5]A�Z�;��p�PPXS�i	@"�c|���G�+17�(s�9:�>�cQXn�l�BNg�*��|n���Fw�����~:ƴ�(3���.�W�	n�8�r ��tP�YRs��W�oz� }/��~ؤ����`��j0�`&]�Z�Ӌ��d,�Mo�g��)�&����]�E�݆|����u!l51w�4��x	(� Q["���$���fsh�"táMu�X��½���K?Ņ�'P�fD��6���#�w=�f�>���ܼ�����(�6`k�4��}��v�zI!�����t2t
6T:��1Cg�H�����a�<�[Z����7�E���+�r��tI"@H�>��~�Em���VC������E�s��7���t?��X��;�v=����CQ�\\�Y���%$Se�Y\���H�0�A:�`eB�����hvx��~����ؖ�٨���F����'�}n����;�2;Y��e=[Dwӛ�ً%Rx���
[噳���-�V-,ҬS�8MQ3@ ����%7�d��`�N��|�]G"��A��:�[:@s�z%+�w�O�晠IoL`h�^�&f�N0��?��giӀ?lU��Nnca~Y���7�07=��[2�������`�Chv��̷H;�@��%�������ZC��� ���L�xS�����Td�m�8��̽g���y%xnΡo�΍ht@H0���D���9G�ؖgj�ry\�k��;ikf]����lY�i�G�hF�#� � rjt�����9�m��;��V�j6�����{��9�	�2j�d��[<�k_���<rl�b�f��>��)C��3��|�������ڱp$*����J+�K��ܔP�gob������qݾ}x�ݷ���/`[G7|�!̬n�����j���o���	�?�r���{���+��c�&jؽ�՚�8�X�l��ϝ��-����2H,dNX$�+�� ό���ud�Ϣ�:�Rq�n��q#*���6�p����O�����"8�o��~�����X�����1]H��{�SW���+.u<�5=�龲��.4�e'��Uc��Ӈ���h����i\�tQZ��;��*t��9�Ri�~�x�z�߉���}�ML�N"S̊c�k�^<�������W��o�E��ĥ�KX�,!�1�����ߵ�k�(�ߪx=�q�[����@HՈ�>�l`sa��e���&,����$,��UψSh�R>��J��`���=6���@r��rya�WW�}x�{�|�����X�o��&��(7�&Y�֌�X4��Z	"")A#_K�9Ц�0�Bn��)�6Qxn׽�W��xb1H�2qyh�M1�l�m�m�cG�Ĥ$��
U��;�∖�S����l,�b�V5�r�)��x(�v���f��87>6tq�:+�*pX���0�rG�|E;�����؜J��J�H�66�!�ֆ�x�bE�8���Q�16.��5ΐlp�FWA6�U���S�*Ő&�Z��ɻ�5�V��4���I&�B�⪐k�l��+��C���cA1_����k
����Lq�]�ʰ"���9��ōfQZe��|�|��4�D�����M�fe��{b���#�J��)p����4��9-�$�<� �r���Q4Ά�19��,���GĶA��F�<p�^,,�h�(��E��P���C�p$9�ֺq�b�J��/
�Y#D�X��.D�����x��a�q*Ģ��$w�礞�^m��5o�ې�GGV���kMp��L"nP��\]iz�~�F��Ԙ[�=��$o�M�"�(UI[(	$��E$��[�X�z�� m�-��)C�fe6b>�*����bC��Z��dl.7Cԣ ܸR��v
U�VXS�h�\B8ȵP�0�^�l���2���,=�� ʍ�l8e].	�6�pX�
	��z�t:��FgG��0&���_M����F�*�IM��z��*~;<ހ��,n�a���L��Y9l��ɹ��do�Ci-���rq�ܱZ��,,	>8��ٴԄ�G�V̜=�so��3z=.(t?�>b�WDL+�ȷTaWnM��7�~3��u�&/<�4N���N'�.�4Y�D
��N�v��=p�V�	�ؒ�@1{���ӂ�� ��|��SSF͍&t|f��Z�j���	(�<Mg����z�݃ٹ%����H&�؈�P*Uu-���L�m�N�āa��t
����X,Bw��=B>�@�R�Bf5J�bIgd0���:gE�w���cf~//bc#�l�*Z9�Y�jY�4e;j �9w��Z�
�d����9H@��ԞM�Z��C[ďѱ��M��Lk/��������6�cjf���&&�g�ɒ�Xo9/2T�L&��56�_��W��̳�˅�R��^>WMRB)Z6��,���d�hbN=��.�kX{�ո�]+�j��3�GGċ{'p���@��V�F�<#���J�+�{���4i���ڒ6��E� 9�U�\�1?������.NN���,6�>fw�B4��5�Ȭ5����.2ش1��P���&u>�4=�0Sy�8�u:�4KU4
%4s��ݟ��G����؎_��౧������m��.�>ah`���~j�A7vl���?�i\� ^{���駰w|_x�a�2�?�'J��׿����;o��b�����h�Ӎ݆�HHT�L��?�\݊�XO<}�^��;HF�#��t�����薽#/r%������PM���؄�����������(���r��d������=������0����)�C{[H���U<��c�x��P
���߽{�8��I~�f��"�Fy��v�ѩS����7h�Z����ܜFY�J�H�=X^\ҟ|�i��Y�؆��#����ϡ���fkǹ�s�xm.?zv�7ڇ�L�rN��(�mDG�L���9MՍU$f�Q�������4ʅu�����N:y�:R0�@���� V�[�9S�*���jy�ڔ<�q�I�R`��q��q�s�F���R|C��b��Vr&y���G�j?��`>����2%Z_�yP�}(��ߋ�<�iڬ=�Rc`UE�9}3����|K�*.x�Q��Q#�d�#�K��X2%+�d<�P�]E.�k��#�ފ�'%��� ��(?���H7�V�P�r���$��`'���M�/�/h8���P�,c�A�
��������"�����..5,&�r,
�],�(Tr*VH'	�]��������7V"�~�ȖST�%Q�Xܚ ��k��e�3�!ڣal��s�r�^w�R�v�܊��ʏ�ut��p"`�0��x�k��B&a�<l�d�H[3�,nYl��Lyp��X����'w�º��i��r̨J����4�+���2A��fW3�恮1�=mҌ�#���&��e@�y0R��p��_�$�^Ŗ����;b)�9a*j��� IcT�G�:*��������}U���>:�.cqע�m!�,@DH��;'U�ㄏ=\�YdQ�BC�|D��1H!jň�I�W�u�b���L��G�6��!ѕ��"e�k(i�K�]3�i�v��&ʜ*I�c��a��M6�'��ze�*h�L/���<5�p`�)bn:������E��k䔏�:<n�����FE͏�eqM��L�d�T@�φ�)%:�Ҩ� �����P�Q�c����rW+����*��Zʩ�IX5CN�x��vƿs�m�'K�?Y�3�ȼFi>���M�5i�e=�D��|�k�� ![!;0O��o �"BL>o�RpmQ[W�3&�9-���V|��|t�8���ہﾃ>�}d67�a*2D�!h�p��sp�)L^��ܵY�������V�P�~�aY��
�0��6F'��5�ϫYf3�t``��^�8�1��䏰��p9bX^K�g8�n	Lh��XkѬ�4��0atw�~��;5eތ�h�N�	���(�����/:���v1����_~�s ܨVL#+�H�V�l�9yf�X�*T�B�n��xր��b	��٬��#=x�+�G�p?�]<��{NڜA����;�هB[8��W��g�W8}�*��"�U� �L�āM{�&�����>�(B�6����x���155�}?m�Y�S�S�Ŧ������%���OE�]*��z�&NSz�E�pG����n��b`[7�C�,گL���27 � \��|�l��.?4����0&$�
�r��ӀK4G�Rm`ys�O|�+�K�03�kKkȗ������4�嵧s^!��l�j����,V+�1�MUz�޴�u隩�^>Ӆ
�X��{�>��_������� ��_{w�{?|��g׎qt��p��G�o�^��ʋ���{FC^��㋟�4��F���8�����7�,��'ψ}`�u��^8wQ��ޞ.�`Y��8uS�A��ՎLŊ�xO��$�?�
�g��͢��1���<9sx�ؚ��瑘:�Bl(��RO�Z��Ƅb�<�~X\�C���r�p٫���αA�㺃�ePF�T`#��?�����{߾}�.���Q�0y�gϞ��Ғ6鲜Nr:8����هP$��9���BcFFw�KNf�����8�<*y�����:�l�( J:5����$�;�P��p��<Ws�em�y ��A,r,Zm��Λ
v�-Ah�T���������֮^�a��c(���(�`�V����I�N�
2eS@>#|���������ٝ~��!X�D.j�:�8x�m���kB���4�2��q��P�8�_q��%^&��mQQ�lE/b��aB6.�Z����@�\�B^�;-ȉ����e�����.�A0d2�R1���H�_�#����Z�����s��P@��)�M<�$���\G�W�q	a�&LC���\)���(�Vvr���Q�d���G�qw�4��2��rLlv;e1�@&�6�܊HE����t7	n~|�`����;
`Ea���׉h��ɏ`X["�A6[�0�V��T��dS E�B��2�]�-�)`�i�>4ԃ�C��<u�����²��t�ry|:89Q�iLd<���9���œ���Z2͇����%rdj	�~�"B��ovg
)��zո��2z�I&N�Bj��l��~��tR�i�(�g�JjK��x��d1O�}u{�f�r�L�8�Y�h�D�`Y#��7�����D~m�3��SP�,�=�'���|���r���}��$]�UQNjV��)Sj�F��@�&=�6�6�(�I�r��r	e$��|�E"�L/ͫ�&���8Q�V�kgS��+*��Y(�n�F�E��Ċ��'��n�G�l�PG�()��hI��բM��.I�cXe�4�ݪe�`���,��`qu����Ph�#oQ
8=�c�K�X3m
["A,�f��:pϒ�d�p�4P�Z-K�
sY�f	�BM:t�Ot��{p�|��j.�)�-^Sԓ�%��J:8�!��HnO�G�Zw�iq��&����7#6�N���h�� �쁎m6��Q��x�Q��g>���o�A&z�oi8wO��TP#a�#��y�KY9�:�����{�B|}����~|J����û�`��7����s���g�ѬҶ�
G�.�WgЇ�#B��y�%�ϑ>E��k��A��AM�y��Fw!�މ�'N����rP8��Q��-/��o�I#2��A��A���ۇ�t�*d���l�U�X�    IDAT,5�SIsY��qO/�n*����ݳg.L�?|��^QC�Y�;��6W�o��������E��tr$2�j�Yd3Y�bG6We
��G���������܋/�{�{�1�
ػ��x�_GOw7.����w��#S&0T�3�i4����sa���*��������܅�x��������@'-<��8Q��?�گ90�A��MN�\�v�ȦXg0�)���'?��v+U��1����h,"�H!�+ɱ*���⒞��f�U'p
PB1o���'댎�vtwv�>�-2�]���
ɡ<_a.K+�q|t�2^z�L.��Ɲ�3u_
��<��ې{"�	�E5�;^k�EF��}�M4I�e�U�j�\/T���*����'��_��_�������ɹ�O��;�wl>u�}���?��x��p����}{��/<"�������\�����pߐ
�t����qJ:?��`&��١|#.���݁<�N�+I੿��~����G�D!R�����EE�i~�MAze��KȬ]E#?T��5
,M���5���0Fv����\�Z��طs�=]ؽs\�"�T��Sb�������D7��k�҉[���]�ũ -@ҿdB0�1���9=�>,^*�I��^�F,�D*�l&���^l�1�H(,i �r���Kk���.b��t'O]��F�C{P,�p��<fW2��#��G�;f7��R��-´F�҃P��F��k����֮^�3����C���r�!OI��F��Jcg�D��k�<�������"���ARH=� ^;:;��ϗ���q��[q�C��tc��2ż���t 6�QW�[��G�A������I3�_����J�߬!�K�Ҩ�A��u{��ak&~|;�f���4�GV�b��,Z%�S�K�|~�#�}8r�������b��E�%S�EK��Έ���"�U�c�����/T����K�&��� o��Q�&G�>�[�0d��������/�Qk�����/d5! M��hY���Ul�'��gu�8���3�J"g<dt�K���s[����v(�F�6�D��ȥ8jO�w�`\�(R����j<H�"�k�
�	`t;��{�t]����A�)�dpi1�^mp�_����+�Ӌ\�����@���ϠɊ�'oW��ƝJ(m�y�$�E1$�Ă��IS�RAN<�2���̉(����O�2-~*�<�#ѩ�1�/�Q��[bv>�*VC�QB��E�YR o:q��gC��
� ���
�f��3C�D�nO@��5�ԏ�X��DץF����ynMH��u�ف�5lN�b�����'B�*d�K�E>;�p���� �+R�v ����W�;(�e��3�7��-� �,������?߈�M!J���V�9���C��]j���;YgM��}S�,�8�<`%k2	�
�.���S2��e���k~��
�z!'_�#���6�M&��״��ϡJ�"��e�؝��������Ӏ[�Ϫ�J��u��m,b�I�]ᤌ,�Rh�`�B4fY wcN@T�4��܈�4q/�d��1?S�S�2	�a��J��5t<��-���q3!�Ur���\���:��]���i5V	�h���7�+_�2�G�ceisS׌�����`P^韛�V�XMbuae
�9ղ4�'��iG4�Go7�Z�o��*56n�[q6FL�us�hw�ޏ��D8Ԏ��/����'��A���f3(Pצ�+r�yQ���³��d>{����nVq*����%#��4�NƑJ%Dg�n���B��nGov�:���cx��	���8w���ܚi�7�#Q�Y��X�S���y>�_�9I���;A	j[��������O�{������.�	LMNcdhXxc���o~�w��Եu��w�/��:��!�������r����'���o��o⡇��:yu
�?�~��O�����
H�B`� ���F�N��STA����,��vR1����dp��~�s�����(�~����9	�I���
X]����<�ԸٜbeLO^C.�F�M<����z��M�������3'���]���AWO�r-BA꼀ٕ>8}Sk�<����F����=�C�S�ZD��7�B�N_@��|��L����=i����tG���R�l�r��?��~��?�2!��k�|���bjv���X?�����n�.������go�_Ѕ���?|���/邞8u���p��>i�.M"y�b�.i~f�͘
ː?�p8d6-�Uvَl���������<�M��L9���%Z�o6^Z�XRIc}�
+�Ȯ^E37g��FAM��Lv�6!o��{btl�l4S�l��w���;��o�W\/>�D|��?�>�~�i9r���g���@�N4F�YP��v,/t� >�<��������6�ql�cr:��6��]����)T2�ʢ�)�k��:X�����ꡠ�lza�ki�<LA,���E�/g�
�cp�u�l��z6�a�	��L��kޤ��Ө�+Ed7W����%���E!��F~h�d���EQ=�q[$R xh�3��J2��A���B�@;F�Ɛ�䱞�a�����A3��Z*�D~��F�Ƶ�F�vډѓ�v�䐷�:���3�����eiV�� ����ۺ����!�R��,,�����A��J;.��K��3E��*����6��8�Ѻ����!䜼X��!ξ\T�e�P��_[���S�[\� nK��Q*�lDT�ܒ�R� 赡+�C{ă��z���\F��$eڠ��:��2Ւ��j�&���D"��K
H�k����ʱ�#z!z�(R�J��kBkX8��k"g��p5�ť�������t�(��FG�'9ldrB~��r��uF�ķe��煿���� �pHD�5:���nHd��)���"���O��1t�X.�������p3�5���?Z�Y����iW��"W�b!/jC������!C����˽"
a-�@&[��a�r������	6�>$_ȠXN����}�ެp$otQ�r���;Ȥ[����I����fF��1��^"]����_HgQ(WP����>u{���c��|��(�OL����{�L����7�SK4ɕ�+Y�=FwG��K^N�H�Z^[��i+����PD:������A~���ɥƇ���%�'b�f��i*[HG1�����.� :�P<�&K���<�j$)$�)��h{��f��͍c|�m`J����uN��K���@�m����#]��߱�bR-'	nPc�Y�����!�T6�������+�GZO�����u��l��� 0�e,�I�C��sM���j�WT^G8���w��+�Q��������%ңx�
�
t��Q�����}A7f�|����$cJyeQbͦ&7�~N�(R���^_�^���~|���d�i�4�;��L���.�����<��	BU�O�P�q�[�-FI�ΥSp;���B��C&|�*�6��"J� ?�5dN�R���\^ �e��rhp�g�H�Rǵ��h�$,�ޑ�$�ͥ[�1����?f�  �M�����at��#�Ƶ�9,���G=���"ړ�����${6�f�e�S(��|J�ti�hSD��H�L��p�O�������c7�ǵ�%<�����[��ge�Ix�.|��_���܇d&�������g^@�lR6y/y��Z���Ƿ��-џ	�||�,^y�U���I���!Q�j�E1��f>Ӗ�֩�����(��pYq�-7��i�ph�4� �-Q��q��5����X�'�c�Oj�������Sѥ��#HG��O�*0�!
?oq�@�T(�؎q�ݿ;�G1�}7=��H
�&2�r�������ƻ'O����*���)A$�:����"��.��!��� h: �%�a���<m5�\�r�M���7������4��[������x�}w�k��#_��.V�3x�W1�4-�W.��!\���0~��q��g�"ab|��
��4�n��vb���,gg�C�ɀ�Ć�M��/�t��?x��dӨ�o��0�	#Í}6��6�f5����HΞGi�*P\j	Xjy�)�O�������oCãh��l��Ã���q��>Y�Tk<�{�<�ԓB�����q�]w��r��L�yZ��`'֊���%x�.���s�qmzR8�|@��6D;��nS�J��M���s��?�LGL���F����f��N���2���t�D�wD�!{0�z��J!�P9�a�H���ZB9�Bfi��e��)s� ��̎n�93wD���;��&�ո��Ł��<���&yJ���m�3��I�!8��{Py�J�t��DZA�؈N

9�F���ل�m�.l�}�7��r���:��c�PƷ�IQ.V�2ʦ���M[�g�i�B"ml��>أP��p�U6��ӂ�`9m�|��� ���0��뛅7��d�f��"�T�%�`��� �a\��dS9�������ͥƆ�fY�Y��{hy5l��5��5T��Mߘ3�H��Gg09��J���M�dl
��ӕ��kC���'�O�^�PF�֜��t���̦7�#�l��I̮��H���TJD��L�Ѩ�f,��EoWD�!����D@[�߬�ǑLet��E�n��ZL6��B����+W�v�W§�����o��(I��l5��2Fj��,w�:R�M���ub�	l��Ŋ�I.�D�L�Ħ�T�XX�D*A]	���>ن�!|�
�.���>��x��w�4V}�r�jV���h�&-����?�=+_�N�k
@K�p ۶��V�������d���̆�� ����O��F-��L�j����סtꚖ��tqJ![D�J0�=���c�{��}�=���'�X���
��һ��bc0���k3��}w8iqj�Nx� ����Ζ�g��n�Y�ժ��c��ƛ�S#��<z�;�w�n=��Gs/����{����̼x�ܛ��z!�O�A����l�+���bp��a �/�����fF��&�MR�H�2Ϲv�G�4��X4�V�<�R9�Ξ(���������z�-M��`T�ܴ#���3��nNh�c`#�h��2O0t'�$�VV+�2�v��RCZ��9�{�,�9h�*r(<1�iB!_��Q�ytx�� 6so=�4���}�36&+q^�D2�D6�d6�*�*�>�)P[��rA`���6�|�Ql@��]o�3��8wu
3KKX؈�V���р�#������C�y�pl���t3A��I��Y �ꑠ�t͖iVԿp
K=�^���5�Ɛ���v���i�F��JǴ֕�S΋ۿE��}3��Zg�W�1t�2璦.������{õF�	;R�A~�ڢ�ɜ�֪py��E&��TI{�CN�YDk�4��|�_���o(/cfn�����*�ں	P�'���ǿ��7�������?E1�9�]��S'��Rf��z�ȗƃ~J�6A�w�y�s3s�H��2i�T�&�7 ��WL��s����ͦ6��Xp�7���,����FM\S��YXF�a���><s�t�\�1
	���2���C�熇��\�xj)81cC���VJ�y�r4'ڦ�ɍ��g\�<��<v��s����=�Z�:p��)���W��VKe03;�B�, ����֜.x��#�<�q6�e6V�����ojʨ�!�q�S�����/��П�����>��o��o���g��GF����t(�7�w��ӅJx�������*�m���B*я�����~�$q��BXN/�V�כx��8~bu{|�m�e�jl���Dpt?�y(�*!�6��+��9�@2�٪�!P����^Hm�������(�"!;��f|���X�,�f]H���s�=��>������4&&&4�f�QM���-v{%���mzn��˺�]]�'cXY_�Ȕ{:G�p�@P�%rω�p��7��#��Ҧ288���D����`��q��5|t�
�WR��ic�7ڏ`�v$�Q��X3#�V�޲�d�B�b�BRL�\�A��5X�)4�����b185�iN�H$u ���䴽D���FOW�l8��
��v�>p7�-Q19�B�[�{E}�p#e��5u�-����{j���}����>�Hw� ��Awԋ�C���+��Z�"�-a~)�W�ˣA��,K��;(Yt�Q���(>�E:�0������Jj�Q(�j��3�.�Y��� �F(�/��o}�S����J����w�)lK�+{�q�]�HfrL"�����@&WF"�G�^C��!dVtE����b�k��]ũ��X������
H�F�o$��`o�Ý��A�i���|�|	M�hAghl y躉�Y��X	g�\��ʚ���GA����VB$�Ǝ�^�w" �C>�ս�F;��z�L�d��g��^N�X8�����|i����?��܊��.�_#Yyfۍ��P�-�9�`��D��a�d���&
٤���Fp�!�F����H}r;��;���^~���N�ås��������`�a�M6m���ׂ�;�q`�x<f9_��D�d�p=�~��3/#�䨼��GE�Â��^��9��n6i���07��ɹ⩢\`(����-{Bf9��o��㶠��c��6�
�����S��]A*�Ք��%����mlC1GCj��'݌NlQ8h�KD� R��6S�]XD2�E�\����<�gx<a8��36ׄ��l�1��eP�
R��D/�]�14 zD(�W�5*��Y��C���FK+�XYO�Mf�����$�q��}�/� �)94.YF�Λ�OQ�5NY����e�beQ�������|6�tbU�]�!��vhm��#�@,�����
N��67Ә�O�nʙ�nC�#���0��U�;\��H[ u������6~ �f�����D|#�x��	�^9�\�9���1s�}\y�5L����n�ݪI6i~�L
�l�TR�����_�LOg3X[_Q���m��;OR-�b1,s�V.#U(�zA?�R�,�h�lX<���s�!���|�hXI���CrVZv�O29��a��d+hR|}6N���T���DZi2,�9�k�rp�=Ғ9)���a�l[��n�8Q+�Sc,�Z�@|M| 辣` ��
U�.�*�Ղ�2֔�J��Ki�<��ሦ\l��q�I0cea��/�{���g����Y�W�.�?z	��>��T�k8v�]������ݓ?��x�mĖ��ޒWȓ�UCg>q��
n�e�ۍ�W'��K/���?D2������ݑ�sch�N�䖳�F,<W�����1�}׭8�{����*�����S�29����l�B��4��y��64 '3�iD�>�N5��s�!$�"����y.HA*$R�	B+���@)�Mt����#�3�7��#;�F��O/�puj���6�y�$66�� ��{� :-�I��X�4�0�٢����i��
��j�ݲ���ˏ��W��.��x��o�l��?y����{ꩿ�H�n���{�����3Vݖh�F~t�ld�s]��������[!��r���d�YoW=�n��F�wwh�Ǯ�/�Y�����vc9��x�)m����0���ǩ��R�\�*���&O����j�D�[[6Ov�OBW�d92ف������S�ނ�n�Ai���XX��w��x���dz��w�U�A,�����'���O�D�@�˫��������qÍ������5iH��%��[�ƴe/W�0���l:/����\ n�D$�"���F�̔��'05��d��� ވ��Ӌ�<��@����nm��m�R@|v��/ �H �/��iЫ��Y:J(��x	K�k���Q�Tatkp�`��T��ay�W�6�?v3n|��v�o,k�D��.N �#��+q���VS#b���5VXj�V~J�L=x��    IDAT�F��w3��۷��ÚJ6W���&>:}����PR:soW}�m��Vz��S#"9tC*PH��G��!��HA>+�H$���(z�"���J��$l����ά��W��F��`t �_�.YvG�Rmnv����}��R�Kk%֨��!�	�(�v�B�RF$l��۱o|ȰKn$��Ss�:����8<
���:��`�H/�yL!�*ԑ*�P��R�F�d�B��0������z:����X�eష)h���:Ρ�+�B{���ٳ�cC�����@KM�ኳYX�X�4�a>X���X/L�8&��t{�0T�����@G�V �PFw����r��T.��D��C�سk� ��8�l�i#ɉ�>��sPx�����9��8�Ņ�%+\� �mm*��0d{�c����ؽc m>�4\+jd�m��M-�)��3i4�^:13����U	�����$�iS3��8"a��	�J���L�o O��ƟA�#8�#V��V5iE:�~�����3�@��`f:���U�?)��v�F�p��>�8�O7�O��Y>�jdN���&��<��`Qǐ%��XR�/��x
��r>/n5-�5�i|��7�(��Po��`h[��(�g�W�젡�7ܗ��*|�嚳/`~i�+XZ�T�G�
�E;1gi&%��K��kĐ�n9��Nѯ�����J�J[�g�PBwg;Ƿ+�gD���94j��HY�4��D"�SggpmjIϬ����.�&uH4o���27��CC��E��\���K��8��E��XX��ZC�ŒbG��+oæɵ�RG�^2����k�Us��G>���w���e
j�i7J�)!���:����c��5))���xO�|۬�n�O��Ӵ;QmZ�-�����x��/;K��R�f��d��kѸ�W|g��[�5����8<;H'�Q*"�J��d���4�V�h$�tg�,+y�9�M���ێbd��T�#���Im�r�K�E 5ԣ��-�q�tH�B�̜�w4&��A���@+��M\���ȰQH�Ӊ|�"[�k���j��><��~���w�8^}�E�,^S&Ӿ[n��o��]p�������3�1�����ؽ�����~��Oj��6�n���
�>�Ʒ������`׮	�it�y���x��gq��G�	r?���P�-j]��l�Z��%QV�"���=�Cw��3$�bz�2~��ϰ����D��6�f�`�-J��UÃ}��hG���c��4��}N�؄s�xܤ�D�,����2����5McSϠ2Z�WJ�*8Ь������#8v�n��&t�w���V��;�ěo��ǧ�#�Y@����.�'�Ȗh��S�)T&���V5�b�!(�P/2���Z.Q���CO|�k��{�0�={|��<��o���G��ݏ���	���i�w���(vn�X�ş~�?����������A3��51�ߋ�����92iT��Iڐj�t/�6�E��W����+�e�p��DQ"�A�#��EH]N�uؚ%�g������PZ�)X[��������w����E	{�g�0��p��
?�b9^][]�_��_��?�7܀щZhD/���ܴrH������\����uو�sy-�cw܆D"&A������ |� �$V�64rB^)#c0�+����w�����`6D�PE�f�z<���1��k���P����=E�T5q���C+>
��k��^~��z��i�^<�f.Ҳ��9i�æ�Qc�Ƒ)�kt�u�z$ʥ�o�"�as�e'��)�����>�����'�w�0�N{LS��C�T��tYxj}���Y��ㆀ"⭆���n���e���ƀf	�Q/���ػk}�a��t�������~��6s��11��j c����/4��b�@��`�d���{�w����r��ZelO�B7Z��6��������d3�u�㧯�ęS���Ѱ�P�1v���)�-E�tc�� �AjS�8ـ��}'N����3H$J�l��Q
��Ò�}�Cp٭Hnn�5��e||qsk99>P�M���G_��va�H���ЧLق\�<����Q.�v;�sZ4ዴG��Ӆx���/Lbzq��^O �ZI�ug�O���n�Y�yϗ���X�4��V��4E��-q���M��/#_$u�g��V�ֺ��*0�)�b�t����F���ń2	l��>W���ct�;Ǉ1� jri!�Sk�Â{�qY3�sU�ry+��ep��$�;}���xPj9u8�N����6�v!����M�:)N�F!�Z�l�jHgJp��X�e��M�.�I�ka ґC�p`�6Ж�B[���U\���ܥYĒ9��t}I��s��$���h�����.tw���vY�3Q) W'1=��X"gP�FE�{�{��T��kDd�f=�I��L+�$�I��l�t�"�a���&.L�c�\�<iv�Dձ���@*�S5:�2zB�݁p���955���Q�E1?��l����.��t)�$м��Ç�Ƶ�x�a��>�N՘� ¥�*�D���ЄL�`�N��I�att�aJ�I�&�[�
�����Of#��8�H�H�{�#��h ��_�l�t�6��g�+U7S���������P\\k_�(��,�
K@�Q�gi�ubQM���2p���^3TR��J�F��"�3�q��~�Kc����U�=��,R#t�z��m��p{�p��B*�x��6T���p���{�����pz<���aw��0��'���&gP-����!�4�{&{��譄u�ʤ�㚑��p�a���E[5+&O�{
��h�(~��X���h&��S�MD��O���c�qY��A����R*�%l�0-}5�$p�`���"�u7'�l�9(X[p�����IlX�M�F�&;��ٜX����o��/����ѱm ��ˏ��{�mX]^��?��_~��\���������ؽ�:||v��c��
%�r�P-ep�Λ��~�[23y�����s/ ��A.��#���w߁�>�����_6�;���+�aan	�no@���VNIrw4�rԡŨÊ�^����r="!��^>��^y	�\�Zl�`��rJ#hJ��]�j��v{m/���Ōhsl��v���E�7?�.sm"6��e5����q7ds\�xs�K��d���ie���cc��֣x��{18ԧ{W)Wq��4~���|~���{qqvk�J<�9K���aU(�?� :�!��^d3PD-�,���#���/~���7������Ϟ�����}����W�d���m���hқ�)m�[���k����N��#��Sx�ݏ�+��d���v&箧��{�>�3!G�r!��ϭDN����D�T����z��\/�v�+%xC]�s�g�K/�fM�Mh�W�:�QF[���&���;���fa�V�ޛrB��S����(�"Q!)��z�!�꣏`�D?Ƭ[c���E<���p��8�cccz�Ñ6���B�Q������4V�V����10Ǒ�ƑKtte�JՒ��N�%7��Ga����qj���,������Do���B()D����z�?�V�(�� W����텷�ug@(�l
��FQ)tV�4ds�>u�˗Dfkҝ'�&�yX�UY�jR`"bM���&��-JST���vо�#%Z��uȢ�g(�#�݅��%�+��Ϲ��r�lu�|���CdGX5v��B"ԫƇ�E��u$�k�{��� �a'F��`�?��ύ,Gtu�&���!6��% ���!.��h?z;B���So
�[�L*񒖥�T�Ix��Ƶ���0 o܁�?4��G� [���UP��x�ͬ����G*�"�Z/��ӈl8�k�����0K�O'g���{�13G����7�6&_���Lal{'n8�}��XY�ǵ'���¹�eX�~x�4d�����n�th'z�L�m��!Q��z�ҵY,��JL�ඔ16L�_��E\~:�Tq��%\���B�h�_��{�w�F{�&{���Z�l������xV����������>���G#���e��5#ԓ���P9�8Vx�L�cWWqfmT�9%Y�ڻ#C�URB�-MN��X_M����=��49�/�-��c~ur/��B�-�V�MC ��´U;�n�PW��t8ԫp#�*$���ėד)Q�(<�%��_X�f<m&d�M8,�56�lp��	rk�9+.M-�����k�+�v��v�4�����ng���D�M��\�.����"R�Q3dA�oí7�8�F/~�.;5PK�"[�m*�?�((en�[��RU��{������Z�R"�|Á�ë��o�.p��j!���;���M���AjKC	��#g^Aӊx,��)�? DЌ�-�>i�D�X�gV0��,7�T����t^BgM~XŴ>d5-�*�SOѩ&LAm5
*�*E�cJ�����{|HS=�������F�P*�~�m2O	!�c��c��KǦ S�����:>��<N���b͊�h��}5�-���6��s�ggcE��dO�ik+�ݼz!�
ڴ�L`�L��MpH'�c� W=�@��^��Oމ��X���O��>���q�l&H�����ɄY��VЙK�k�(g,�Bܿ)l�yO1/')�Ѯ^0��.f�s�Hl&Q�0ܐŴI�%��i1�?�u�
ɲY6�Ee�h<%�zS�|�W>34�P^J�r����q�������c�F.�B�V�Ή�x�K�áC{����JZ'�4Y�p��y\h��dS�ߣfQ�ԑ�pT_����&d����z�K<��r��{���d��B�"3������B����������~%K�kul�Vq�����+���E��8>:sO��\��E�aA&�Dqs	7�q3~�w�7�=n|�O��<����<v�V|�_�ѣGE�d�P�T�����^{/��
&�Έ>�F�v��c�0;�	 �s�����e0�s���_�m�݄pЇb1���Y����p���&�j�᠘������t�͸��!��e�4wH�TLkO�A���%s�(СKnc��h <l�N����%`-������$E,�%���B���,�_zq���������h����8��9����p��Q��և�����ƳJ@�E}x	�UE�$�,��r�X[�B7��}�u�����_�����=��O�|���Ñ8m^��<x@7��X�;�M�i-�p"M.a:��G�#�U�x��H�uv���qQ6\�|N�Z���ф�v�+6̮�pq����0�T��e܈�Vʚ�J��C�h�	C��4����O�t�}�Jq�k%��[����Z��Z-�!G����Q�-7��|�8�oHE����"N�8�^xN��c�;�s�N5lJ�l�8!�����
f&�Z��2򥢊�={v���:$g�g�P1����#��
[���g�N�������?�O~�Sr����Y,.��w�v�����S����P&��B��D��m}۱�-�n���P$mF�ldD��T�k��͹��a�d`A�z�z�&��+�!h�qn5�b�_n�ː]"W��[�<Z��_�;��\�ɻq����s4��NЖ7��Z"�H����\&��	�_��-��64	C�P�"�����D�ߊm�m�F[ȧ܇r݂��,�=y���XM�n���H/ڃN�}��M�nD�K�,����d��K"Y������e3�Z;wta��6���4w�C��[aq�p����݅
��v��i�]u�m�¡�D}N�H%�6��T�����ӓ�6�F�	�/
��#j�b9�����0&F1����/�,`�8��E\�Y�U��ZNc�7��vb�0���2�+%||�2.O��}�(@�50�ƞ����D�y SK����EL��>�n���A�C]*<{:��jdl��Μ�ćg.a#���δh��E����#j�g������q�D���p���C���D9��5)h�
*��6�,�l�v���C����&���@�l��b���+W�����w�Б=�t���{��P�Z099���\F*SVC@ABY8��M��5��b|��z���VI\�_��\�8n�*B3��fڅ�'�9��	��$K�f�K�پ�h9�(�[��K��q�!C�2\�\u,&�Z�#�\Cw���T�L�7Ӛ�n��m�|y��_���z	��vp�����@9�1s�Gڅ��9�l�kO�t�U���@ c�#r��R<�)W�C62y\]Xŕ�8���!��^�*XkE�R	x��!���~�\ �N+\���	*������D���!���� ��CƉ&�zqiW��b3����u5V�7Y��A����� 5:�ְ�R0�# u	p�N*uX&Fq�7 r#����ր�E6�.����^Ęp���nk�6����G��z�iO6���+�x��)L/���py�$F�tܰ�/��i����\���40R��Ǹ�!��V��I�H7_)�M
n%O-���ߍ��=���9��̏��s���y[��g�� ��`@\b>{DO��r��Y岀W�F!��|6�6�>:	z5����,Ъ%�R/�4H{#�LH�m�ݜQ���Ĝ��ݫ9(W��Ӟ�׍Șnk:GZ�:�Ɏ�Z�rV��{�������;;T/�I�i!�<��:���L5f�p�]U��lv��	�d-�{h2�g��n��{\N���و�bҮc�<���S�������.����U3ڒ�KgI��f&��=�US���x�ױ��!�B:�D-��[�����B����}�1��'/jB>�k����q��T,�q(�.�̹Kx��8w�.^��x�����H洄�i1,����i$�_!�A��|�ˏ����}�]X[_3�p��ill����T��@(���vD�AXmu,,N!����c��ppG��P͚�zIS}�at76��PE�&i���`�ت3ج9j�A=�6�*
t"�,c~j�.�`��`j���.|�/ad�:=��$��k����Y\�gqm9�,�-�S�G45�s�0Жu,oM�Z�dlJ�X��;?��_����3!�/?zu�w��w�b�����VڇRDC�x;�I +㚉q�ᨌ�]�gYo��q�Ѓ.#L>r`���j(�s�j���N�Z'b9���\�)��B	�k�*�����F��  ������7�yS��
k� pPhS/
�`V�6�f�'�?��w����MGvb��CӐK���_���,��:��?t��-/�"�LH��Chb�NY�}|�,��`sEj5��#
L���f���!�$wF��H$�<=5��s�-������L���{`e#���]X�����?��;H��>�|���9���<;��"�H �c�IJ�MY�(_(�\>��u:��UG˒,+�)@�H�"@d�.����;�;a'�鞞����^=�_����a�n� 
؝�y�����󼇛wV`ּ0L�P#��"�;��dVR���+�Q�\����f�H�z��F1���*�[0U�f��b�[I�ݼ	��Р,��N��J*� 0�g���)�C�A#s-em���pW'�{�#8��=Ƞ�d!����/��P~��B��i+�s�5��V��!�F�SIj~)!�T�&z$�Fw" ��,�!NT��Сv9����团��L�5������D�d��Z���xd��V���A�e�B�߯\�,d�*'F	�R�=~�:6����^���"1�L�޻���^~{�
��� e�Ξ��^x-M8e�gF�ܜ[��o�����狡EJM��hYA�Kc�	A��=	���s{n��w�-5e�CbѪ�J^��+��!q!ShaymG��{��ٜ������	!%!�jS�B,B��h���F3���L:�=uGF����(�'�lP��vk��< �+�ܬ(x�**��Ŏ�X�A�A�n۳'��R�Zܶ��Si�����B�i���!@}��Q��MhZ���3s�61���=)��DF'�?�@�@��"=�p��m,,m����DD�Gy93R�s�
��`\D���=\����ʺ���^�l����N    IDATr�&(������z��PE#a�'Q�L���0�݁���1�m]2I�{������,4gPҝ)�bC@��~j��Q���F�`e�8��I�����|?$�ݶ����qx�W6�!pb���&�޸����n7\>���J�<;Ƈ�1؝�$S_CA��M�MV̯�ཛ3X�Nð���`%���Q�O�m���9<|nva!|&�]�˻�ާ�����llmK(���)R���^����yn�6����L�i�6,��Z3Poh*����M��,�)���ix���bah%�N�hZ��G<�?z\|m�\�REV��l����=�|2�p7��"=�qdd G�d�æ��00ugo�{�LwH6��-����h�ddn�H�S�����MY�X#ߛ�d����3A�Ԏ[Z�xQ�3��`؅W^�.���K��Z�)?�a>S��p+G?9V�aQ��w���SM��gsBK�9'�2-%آ�� ��[2��q���k�����HCc2��I��ө6 �H�̗�;6��0�����BTR�ڐ�Y�FB���G3����BCj�����U,��
YP�˪�p���o�iV�r>���Ri�,���8���(�~�)��Z�f9�*w8�)d�I��SO=�s�=�|��?� $@ۿ���w�����/9=|��	�ܔA��Y�+�P�����_ċ����޺�b����]�%�Q�%������ob���צ����xw=}���{�E:��SSwp��$�_���V�ԾJ27�{_68�A���A�+�7�Etw&�_��}�i��vb{wo��.\|�k�F����{D=Q�汻��b)�by݃��8Ѱ�Q3j�W�܀��/j�%�''�WaGe0G�/�v.k>��X�Q�̍� I,n8,<$��������Y���cur�H_��/㉇Ǚ��d������y?z�*V��`�r�Q��f7/�[�`��hi�b�uc0�6��=�ؙo}�>��������Է��'��N��~X��ɫ2��%	�13ʞ9 �n	�	��j�`���e�-W�F� ~�,N?���F$ٍ�2��UL8�v$�-\���k��X�i!_!�ϩ�����MREi���$���Xs�^�,߼ �v`5W��D׬�
��B�nҐ�S��`�hX��C����FgGX��}����w|>/�XB�P*���ƺ`�fE0���S(U ��zG�%��2�7�N!_ؗ�_
-�	�ݽ�G���B�ݹ3+��#G�bhd�l	޽��~	�x?W��օ뢍͕Z�io�]pz�����v!Snʕv�Lf���&�Ey"����A�����+	V��T�P[�^*@��>dn�qM��J�e���i������ώ�ge�����Ob����7*�!8h��CMnh14��dX&M\���$)1�bԣ�D�I?i4ʈ���
"�#t ���7��v�%�-���������qt��<x�Ps�����b��.M� Wb�V�ȔH��9��$�E�_)����Ã���X7:Cj���k�9�]���;b-��c�8s�F:�p[��4j�<k��1���W.\��N-�.W@%�����ZC�d�zU&��p #���ܘ���֞�j�mb!�	'���ja�S�h;�)�����I>?ߡx�%���DV�"J��m$����D��BhH'7������NF�k� �9n��eܘ����$C���PN�iz?�e�R=0a������Vp�2�Q^"�P�>3B�jgS�����K�5��Ãy� �\f�����g�rC8��_@��hFGz���Ogj��]���Y�lg`�xa����r�G|85ԍ��L���]Kg05����%є���CqTt����V8�.���|�y~���dCcHC�pߙ����d��2�r����%L�,�ڴ�3�C�8�b!��8>>�#����� 
UG:]D�d`y-��y~ߺ�mBA�4�}Q�&B|�`3�"S���%+�M{������dkz.'�^7���u�#�����]��W09���7��큍�lR�i�?t�?$�u�D����[ť+���lN� ���)yR���N����S��<'8���G| Ys������b3
)0�8RҪ��Y��p��B��et��%	�
y�x�C��A�L��`��L�;����`'��&C��E�)��Hx\V���{9N5�|��M��8�[3�R\p �).�9BIbc"�^�Xפ8⹠�僠��:'DVǢ�awj2J�/��~i6�zj�7��8����-���O��^�ì�染|�V�S��!��-�S��u�[-�9S�;��<(��<��X���s����"���_v6̗>�!2f+�C,�U� م6�p����r`���f��SPޣ�2xa�5�jv6M-1A3h���@��2nT���N��� f�����䦆����u^+N~{�#�ض���� �pz=�կ}�����8����>����ׂ���������SO=����D8����v~ ��d�W��O߼(�Ê^�����=<����O���8{��5L-T��4�<Ei�$�$�����.,#�)!�-����nq��D% � �4CjD5�]_��/����"a���ο��W.!��/�[�}�
~��'pϽg15}��:l����1/Z6V��f�I�����,�$1����HX%)6K����J����y�ܵ|�mĆ��t�i�tւH8�#���!��1yu/��m�\�F<އ��c���?��O��ܜYǿ��ą�wP��K`!�M�[n()�f*HZ݄f�B�A&Y{�����ڗ>�����7�}ϟ���g��N�Od�2�EG�Q�hs����ҬR��i΢��j��YYG�ێ�|���I<��Gp��149��D� J^B�T�L��«o�bi�����#]��N3���7�"R���ݨf�Z�#�q�w�B�[�f�����6���*��$��Y��D�1��a1��c�>6���ݝ	�:{�Luө^y�!�>}ZP�4g�ӫV��C&Z:^z�ٌ0�x��ú�7y9��b���^�>!Jx�P+�K�f�O�`/���1x|�u���9�ý�H1=���d	K�{��J6?|�.t�l����h��m'o�,W���ds4���d�q���6Ѣ���4갘��B4�z]�9x���㝡.��:�BT���M�XX���N��g��ч�C�(c3�+��T9��@�~�!hO{���	X[S.�<r�e
�6R���tC�0���m���+�C,�Dg<(�}6*Â��.�S�Ǎ�ہ�ׂ�#�8{b>��9��ؔM�Zƅ�o��dl�����
X�����"3��8v�_���nT��(�`}{ْ.�Q��Q������pld�/���\4�p�������b7� !��w��+X�"n�R���>		P��|U�g�0Y�r�`��%��hHi�N�^�.�@N���K�K����9p[�����u���5l����̪|�fGHz����^i��"p���&t�6�x��ܼ���/�ԲБ�Fy�.�8��T��l���0��۫`��qH@��<;ju 
�6\J>������G_W{����֨Ѹ�>ɂ�:޿>�듋��2!��]��p��r33�hY�����iI���q:d�mE�Ǉ���BN&��Z��4n�-ana�|�>w-�U&�:�9�*|�I����l�O��S�3>܋X�+^)�xߚ���o"[n���@
�jA���9��D�Y�6�܄�]���N�JyJE�;F���"~'4)����jX��b~uW�2�*�~����u�iZ5$b89>,�W���_`s��w�M�Ɲ�Jy�a	ecրQ�!���N�V�O�.�!R���O`�X�?���R���!��*��:��ctd@��_|CW�7d+E*��6�(�����������[2�Pmv����1TzUbk�tG��G%�$_*A'��j��掐^�6����ϑ����1�˰(2�?r�)�<6�X�'w[�,,'qkzI�/*�&,4	�� M�j�*�6�1�0c��iؘp8�b�P�{��۴9)�ـ�:��Z��^��Ҁ��í�o#��H׸l}��a!H���;�F��1�$��g1�L�L��?���q��-?���D��0�7ᦀ93t�S�(�児�	�V��? �T5�K�6���%����6ى������46-2L��A��U�����Y?�k4U�6e(ԄĂ����ϱ%nh��`cv �:HNgax��Q�7��h�x�j�?�ǉ���ï�_����������o��E"%q#�C�GG,����82�޾Nh�d4[XZ^���i,�m ������r|�G�K��Y�t��YgX&� U���`ye�_������X�E>_�Q��.���r%�R��&\��^�����"��������5��%_��7_õ�kHg�������qA�ӬMi�������	V�j��@��D����$9���ﬨ	Hlk�����p%���Aؠ��<�4��!>P!�h���h�������5�J����*^|�U\9]�>�̳�§?����Ȕ�����y���/�f�C7ȷ�ׅR�.@604�Qd�[�����V��j6Y�����7����~�d�χ��_��������dw{��� ��Ύ�VFݠdH�҅�D+�Pl*}�*l5ͅz���� ������P_�t�,��B4�Z�unΧ��˓Xܨ�藆�+O���G�)"�<�x	֕O�i���6�ckaFy(���b��e<�g&P"B!���q��3,h=�����.z�;�=����J2��h��_ 	��^��E�ϩ*u١PL>RȺeC������r�ǉp������u���W�
Nq�i�$���`8�����lզ�+�XXNc7U<��ȁ�{��7��\Y�jE���&������^7��i9/�z1���J�h���F0�5^�A�
�;u�������*L�k��͠j��^4��!x���ч��n����Z�<*�z��!eZ�0����� x�v}���� eRn������v������ݬPYV6�3����C8<څJ{�j�"�'r��x{o\�o��`\
h��H8��$�er�,N�Za�
�EC���̤%� ](c��Rs��H�MՑ�>���1ĊX2�+]N\�u?~�

JJ�{9e*� �V����⡠�I%���"��24��ί�ki���d���\�����!��x�n;:�L��!���s"����t����-��,�gi��$��nm��O��,a|�[<DE����4WS�K�z��9X~x�4�I��t�����h�=s Z�v��X�Mc���?k$y65Ѭ�P����0�B�Z�լ�h�rn�Vq��&n�����fg�Q�F���A�@�!![�lW&�1=���ހ�OskN��#�����Ah��v�����0�����5�%ɥ�J��N,?��<8�e�KzIS�3�3'��bn ����F;%���?�f��q��-���p�Ip�K���x�':�θ6^k5���sxo�li~��S�y��ѡ>��t����hՉ�4���ǝ�u�,mI��DŤ*�_�eb'�U����=����F������XO�`���|���h8}�����iB6���ܸ��+��(75�Ba)�9��/>�R7���������J����l�o���.%���3%��&��LuE���e�!��""9��MhJC`55P/�e^ۉ�~���vI�Spm./�R\�:���s���h��d^��"�$M����Ȥ�;�x���q�p7�hg ���.~�d*���2�2a����ቲUYN��ٍEC�g%��9[8�IK�R�f	N��
�P�Y��o�(�d[�s9�A1�t3'����64��"mg(��j�Y��L�4>Ϛ�^��L��Sn��b���p�/���;`�@�Zp&�>����{f�ʟ��˵�|Gm�����|�"2Ez��ז&�BW����)�#e&�o�O�������H��5�7�����puϵ���I]t��{df(Xa6K_��W��/�/����?�3��V�@h�כU�E8T�c�>�s�ߋ@�/D��.S~s��Oa;E�_]�Ň��d��)0��m��2�ze/��-�g��AVf�,$/�vYx�ڣ��ܰ�sXѐASz� ����~gO
���{p��5$�)������`����D��"q#�B]+��(A��(�K�<=�bN�|��m�o��������;Ndk-Ec��{�`>3A3�φJ�*Y���\z=a�!x1h�b~j?|�'�~y!g ���g��O~�@'�����?{&����e����bC��Ca�`n�`���XB=�����_��|�D��G�?�������/��'�?�ć�K���Dj�h�!�
����uW|fI+e�"V�Q�T�@����c5��H�d&@[�-x(��&�[2��|/�6���:�.�,�n�qe��6���0��f1r].`s�:�'/�YJ�(�`�e�*%	�0x_X5��a�s��=]��E��+ԡ�8�O~�Y�vv��Bo���ޒ�bnL���"�!)��"�vv�L�J��p���yD6ņ���D<�!ʐ<^X8108�Pz|\��m�*i�g�37�L��@�S�AK�i\�\��V[I�j����� ���C�XE���fE8�b�\����I�!6&��"�B��u�6`��톀�/]$
��SIJ�r�|ß���uR�]�1�U��H��g��a'�%F��^<�ܓ;w�z{;���pXE���A���h���F��0RU�}���߄�"U9	ꎋlȦь�4����Ltg6��-�����='��3���E���ֽ��~��e�#px�"��"'�⁠Q��~C��><.�.�<#<±�<�wuB�H,�@Ѝ�ׄ��C�(b>�z�h�L���vy�޼+XY�9��C*�Js̓,ld�+R�X5!qp�}��gA"�]�)01�Y������~1?"�A/�A����vj�=��յ	�"��LluZ��܇V�bXn���a7[��A$&Q�7�� ��M���h�*�ߡ��!/DfV(U�$�� ��nH��b�q�+Zd�-l�,�?����b�#�
�������L}z}A��r�$�mu���ۘ[�E�cj�9ģ>�+�I��U�9 Zӫצ0y{�Z]&�I���gp�7�V>+=��Ŧ	�J.H&�@�W��. �) S(K�S����	M3�M�.���� ���f�k��X/���R5^��[���u۩�K�}ܐr���G9���S�^,������ǵ�u��4▆���٨��p�Ό�'�E�XDS7!�ӱ���;��X�L���u�,Zl&�2e��uvM�����0��{��fӐJWq��m1䕫fج^as�D�؃'���`u(�-�N�bק�p��*��� l�vP�M|$:n��f���:q���z�173��Y	��;�2�㦐D)�b�^�ʪ!��Ŭ	�efaؐ�ܪ)�Ǌ3GFq����L���	-�6i޿9���hN��Jnm�e�6h�5d����1>֏��A�;�(�,-n �oH��Do�����Υ b��$�$�4uZ�*�@�~pN��B���j�I�;'�,Λ(s0�
�4t�=X�����h��pY��ᆋA�-��K�7@����L�Y���4�ag�k����Kx��?�$Ų�:7c�M��O],W$�@V�1;��l��)bӬ��k|ǕY�@Fx0�� %��{B�J��m���-�L�	I��y�(���f��>U ��/T ��P�H�N��*�u�&`���E�	��ZJb�3� ��[�2f�f���>e�5�����K_��+���o}��d�bvXPmV�)������/����7~���Mt)�d[�TdyQ����}�v��2�����?~?�����+���R5�3��    IDAT��סY�0Z�I�S����'��k��4���1��g�ů���dj`��ܸ9���5��U�|nDQ�A�������@��C��|��=hXjh��(1���$�\V�����M�ڰ��)�x���->�J�G��1��������l ��0À��.������ayn?��˸v�*����������z�'/ /����'�3��I���D��vC@.=��>������_���|�X׺*d�~�����������9��O|���~�ӈ+p�$ �CUjJe{��]� �D\�'fs?�Fڹ9���[�(ds�y���q��'XUÊ�BW��A0�Mfcia��.q�7Y�rE�&j�!z8���8l�^�.l�\���;0W����s)r)�xP�l���(k2� ��tX����������c���w���V�p�u��6177'�Ξn�a)VcM�]��ueE����:]V�vv�;�"����OG� ��4P���dm'��YGW���l�YZč�Y즋�[�.���<3LX��K��4](ևS�L��A��$��zE6n7	!�sw٬��
(���Z]FugMi�qh���.e���(���̦�/�2x-h�����%�P�ŉL��<�1x�8��<�3i�Tr��U7�Kj���	�P5��o'�<��u���62�2n��a$"�:,��i4�ڭ������n��\7��;���.�Bn��N�1Q�Pj���x�'�`u�����?�*js�*4��^�rp#����h��.�.#�˵��:�5��:z�!�F���»_K���\��e0�"!NMa��sapͩ��I��|fɈ禌+Y1�x�RS6�^U	b�"*춋T�#�E<ꃋ�%�Zykܺ����cs;�+�/��������*#�40���P�Lj�5��^����i�;�<-x�״���R�U��֎�Y���8E��r�E'���.&)��s��􇐌�٤��Hn�O�P)��aaXڑ�N�%p���2�rzBXZ�Ǜ��ܗ 7��Z17N@Og>J_4�4�l޿6���T�u%;^����Ν�HĦt�Ōxjf�����v�6�@!�B�RG�Z��KJ��vӨ45�H{���*�t���X�%� �j�^�j�6S9L�Y��ZR���vNo��(`���=t����{��n'K��WEx�!%�J[g���h7�H�`X%���lV�9��<!8]�x�0,�Zv[K<(�c=�i@j
��l7n�a�β��l��86��S�݋��@�Z��E)[[�2��Zč�U�f1(�̔4G��;5�����v���0�>/V�WE�L��&yf�L0]��6~�l�H�t;��n�	Kd���w�3��q���85�@���9�mn���l�1���;K�QvdqJ�?D�̀@��6Q�g�T��#�0�ad2,�]�Ѳ ��㑆@B�^�2��Ɇ����[m��A,+Cq����&��9(	{Kd*����
�������6s���L���C�;ͅP4&hO������b�ڔ�����5��	;�fWk*��r"�����1����I�H�:n�W��~�܉LGɞ�p�B� G@L�jcȉ=,�?�W�>+d�k#BEn	��.Y8&�;���l��jC������C~�2x�(mj�YA.�TK�Y�pe�B"�Wάhp��M&���92LM�!���v6��F-�_����_��H��y�}|��~��t:?���A?���'ŵ��1�ׅo��_Cg�l;+���O�UT5��UQ&P�Q,a���$1����x��Rh��:�����
���fBI�D�%6�a��8rr��?����CG��p����q�*�FvB&e�4��$���KHv���;G(⇍�o�/�@��@�M?�lL N2 $��5
�H��猍@[r ���_��a���Z�(���攻��
�Ll:�l\5����.�\<���t��7~c#g�ÿy�������6��Ț�$3nø!�ĩ�l�AOX��Zn���s~�_���|����GC�O��7�������=1��ǟ�֬��������REBk8m$ݡ�-�II�jECg�[�J�R��K����#?,y9!�u^��s't^2yS��x��7�МQ1gP7kjT�Iި�f4�K礁�?1����ܾ#�������\J�uihdke\5��v;�:6܅�}�	;:��ߏJ�$]8��<�I�����y�֐��p��Л�]����)��e�n���Tj�lZ&����gN�������7�4�-�N���:*5R_�x��ܺ����$��5*��F�l�+%�A�AI��j���B\i�&,]g������{)l��#���Fr�Bh�5˩7Sa��69�~�"TSf�H#�S���Y7�ϏR�%?4 �u�s�������V!�L�(/g�ȕ$�H,jL2��j�D�e@�x�L�Ĵi6�ed4a�Z�AN�]�B��C|���=�H �]��U\�3���e��?;ћ��#��`g~��^����#��W��{7���O�
��Ϧ�U�ܸ�M��gC��%�,�@��{���`h�S��z�*��]R�u��p��R��v	�(�_��fo�w[y�\AXܤǰ0�a��o�JY����eij�����.A)�P+W�;����\�38�	��@��BW4��nI[����4��� I)��1�������Y���n�����C}���4���V�^��:�YJ�8q�����9f0IV��u�{y�v�ʤ)1Ι�qM^V��լɆ�t��Bv?�A���Ō%�d�a�Y����'�`�3��,h��uY]�,.,m����[�_ޕp=��?���(��A�u R�
Na��H����%]�����pb��!'�Zz�x<ChB��F:�wid�ƺ�i��:r�
�u���%�0���I��;e[��J����#���[9�������3�_ޔ�:I�m6$���?�8�Z�LCY��\��]��~�N�s�io)s�">��<z?�A��)�h̝�����l�����I2p5vj��	p����p��0F����ƱR60=���������pt0��>r�!�RV�M���}��2���l$\>�|�Y,�LVE�>�\A�T�m��M��� ��Saj(2�x��)=�.�g3ٻ͖'��6٩�ef[��If*�ڪ��5����C8�C�VF��-L�]����Hf��G:��A�L�Y�r�I=IR2٦Ο�|[��+�;��v�3�0���'��lr�˂�}���)�v~B�kû�N�h�U�!O��R�Ӭ�e5�h�SX�|���pR*ܤ�W�qcG�>�"90dQNz����Ҋ�w���>2�=��x���af	�`�[I�<�L4%7E�s�|6�_/	V��5~-2�����J6���+��k��
$K�N�g�Oj�P8_���ޮ� d�R�����������8a28�	rذ��%�nz��/��9��簋�:��*C��;d���%2?n�[��x����g�q��_�,���G�{���o��d�$���-��빧��>��݆��*�zG���s�y���"�p������F�(\zB4�T��3�D��^�O^~+�ۨ�L0D���%����H�݁Y��	pB��p��8��+_B�`B~�ć޽;+�a��5����Eܞ�B���/�Dw���p Vs58��ň����Lm\�`��l��.��| �����=�<#WlĈ�&��M�����hK��ŭ��O�e���#��i����0{{���0�N᧯^�K/_��t!]�:���l�d�҆f(@��n����{R/�T�y���|�+��w>�s�|����� �wh���SJ�ު��2��{p��i!P�r���������йζA����rZ$Q���x'���n�� ��� #���jMRtÁJӁ[s)����XX/@s�`u2����W]��q�*�حnx�N9��]�޾���@n��,��<X<`��E�Oi�������O���Cp;]��rr)pE��6�ړ������*\�1!S'^4^/Y��3r�[��l�H8(	�^�f��9���^�@9�p��,	�-TY�p�Ey,2�M�pub��u\�\��rJ�@��P �@G�THV�
2�,�������h�hH\�ɭm,�/ ��s.-�a���e<)B\���R@>Ѫs� ����ץ(�Nf?�%V<v��J��o�s����g@�^C�\�iN6_��@r&���͉2u��K��ߤ6�%���Y%X��?7l�4��&���.1fE�NxVa.;�v	���qg}sk���c1a�+��xHB��6���\0<�5`v1��߿��}I&< ��^r8mQh^{��p�������	ٌ|��\똼5#�mfb��ѡ.xm��0��&>>W�?x��+xj�h�l�[Z��h4JJ�f#��;�r��0����-%�c�5 I��9Q�l��&7�Q�ëݱN��J�kXT���&R5̨�[��X��ce#�t�
�n�����;SN���{���ݪ�}<p)��	�㦮Z��1�N�';V�w�<���/N`vi&+͖��I9�{nG�&ʺȑ��Rf�` �B�6H�rH!�qScn"�`t0���[��	�ש�5�by=�K����DV7�^?�VMd:D�����ʳĳ`s{�gW1��ښ���Ɔ�8��ȹ@2���^�2}.	y��H���*C�J͌��K�<1�L�,��:"-$��]Q/�z�"�
�MB"�aniM�X�˗ȗ����Q�=yB�++��M2,�8y{[�2�U�$уBS���<����XDg΂��37��1��)�Z3#����4�,~�$����&���H.��g�e.�cei�]��b�G $�'F�����$�XL�fn�o�K7��.ð��p�9�_����E�.u�ي�$Ц!
�y�/�|�Ď	�*j�hR����5b���`Qa����j�̼��܋A��K��Êýx��a٪2`�dwcaso�w�۰���yê!hQ��h3ͺ.K֊$��[�J-%�`��NL������ިF�@rr��+uO�Wá���*e5���Qk���-��J�<Wex�M�Zl߽�����c]ȥ�������HK8T�`QvK�x(�R��0�.��ϊ�R�X�9�n8�Ԫ,�lajzK˛����3�p3&]���ߓ�>���A��'�ɼ��P�V�	�����&��S�ln|�P��g U��Noo'��Hb)�-+��
Bѱil�O��3��Ѱ_h:3wnA�+�(�i�iW�L~�X)��C�9U��FP�(�7N��p��Ty>Rw����7~�x��GP�+x����O�}��z�y�|�ӟ�P"?��en[J��=��������S�ܥ_�d�Ѿn���J~���ە��ʦ�*���z����/���E��(�U:\���aS�ϧU㠉��z�x����y�˥���h��]�����zVB9Ý^��ek��(�$�<r�T$�_�Ī�i���,�=Rj��j��Ć��8L)kBVD
�������t.ލ�R����1Kj�>w>����v�/��>_��fU<�w�����@���IS���&{���x(�oq�M_[��f�'���o|����G��N�_��o�З���ċo^����v�iG�F�G���'?���n\x�<����He��%�GUΈA���8Wo-$�<��S�;��;�3848��'OH.��K2<��y��ݘ�I�7�qw�(&E��Z���z��V]&B|H$�Ns��`ѧ�\ˉ��MAy{�Z��t�l�x��?��`?N�:���.��:�~3�=pV�F�r�Y���ؽn����ЦT[�����c~~^�8��h)/�A:��ΞN|��:r~~�tZ��9�9u�`T�i�%��@�z3/*��Z)˺:����o�o�{�Տ��	8=��@�gu�_��&�3� u��h��x�F�B�hTudRIl��cc����lC��L��t��U���5m_:N���*��fv?�g>�9�C���hU�Ɇ�Ŝ:�����02���Vs�Q�N��U��4`mc��,�`c���������<ڭ��g�y8B�T��>�7�0���L�E��]��K�7ꃏ	�v���Yd� Y�*Ȅ���*�ޠ�l�Ĭ�-�M�\�<Hh u��l����فD",���s�e�W�&�q#�V�=�ΰ-��kEŽ�9�!x�wqmz�D?ܑ�$��Y/�U/�D�cL��ᥬV�r���=yl��J��(����B�`3��HL�:'3u��ή0z�b��IJ9��6����uT����GnU����v�3�kN�y8;�Π���q�\�AB��/�!�+lؙ2��^�ko]���&b��~U+"ܭ
��@8�B,��3�ٜH(��n?[���Y��b��A$�}G�	�ӄ�ǆH��ǁR���5�,cq#�������*�D�+�x�9-J�*��7qsj^�k]a���D���a����i�E1��_� ������4�C=��6&����*5�u�Zv\�<���I��VYE3��͐���k����;,R����/�
�2��I����Ӆ=� �!'*�*�
i*��y	�Z���v��˯���0�uil��$�^RW��!������]�Y�B�Bt�]?Y�)���<���]����0�����
K�/�X[���;7Q�p��z,83އN�ok�Y/�t�jXp���yi٪	�PL��rQp�񈡙��ĝ�������&�"rS�T(Ѥ���OE/���dg�AT]��8��u:0�ޓm����I��b 걡+h
WG� \!?�6���[q{~6�a�A��SV(�϶��  ��)9��ͳ�dsf�����*�x��Ta$�9�I�N�vC �kN��4͞I�,�ITAY�Hsۛ8���0���<�#ý�A[Y_���;�[\�~jO6�����R��*:>?���8�C#��E�z�
bP���e���-�2��o�/_|	�;��=�V���j�M�
#&���42����5.���8�� �:{�L����I�,�9��D�թ�αC�������H$��[^Z���VW6E
�-$?�H0�H8�B1���9	�c�֡���Y)�����ո�f�J*#�v&�����W�4��=��3�`:aK��H������{T|�צ��;/��_G���'�{
�|�i�9|>*���g�JY��i��޻���^�3����P�1<��C8v�d�L��	u���=]]���)�M����_��w��]��f�0ds��Qc=��� ����8S��Y��"���G��x%�/W����U�	:��$"'����4�+U���s�*���K< �?@L���@<��"��r��~�so��I�w	���^*�#�-Qa]�sE��,�+*�<?\6�����3���^@���݉卼dҰq�ei�(�2��B������F5�Va������o~勿�s�����ߟ��7.����v�;�07��jY�tE��g���z�����)��Wߕ��x� �-ME4��v�M���|����ƕ[��~'�������r%/锜s}N-|�i���4^zc�|q��>9�T��$W7��9��R�p��I FӨ�P�Y���$�'QJ.�lƺ3q�*R�@$�ϝ�Qj�qy�N�R�����/1�?���^�D���Yt��?/^D4�u/�gawθ�|�>���lll���,ҩ]���s���Ԅ�k�jM./o��,��8�E6�Y����-���7h��Q7�219|�� ��M�gh�2d�*�/�C��L�(�p:��Bg�J�)��R.�b2����M�`C�mU�c��C��	}�*_�����r�dC�9tAV�b#��qs�?��M�T�:��]�8�E�*�N��RGo5a�Dj���a	�Z	n�E�a���_�Ύ���{Bza�W*_�%    IDAT���Agȏ��wE�Z�JCL�4�ڱ�,���S�r�.\�(�ހ��(S�AC�(���y]v����N)V;bL_�粓����*�7�.�u)Rϝ:$�׊&xԑ@i�߹t7�6 G�jdZ���!��:�#N;+%5Mcs�ل��Ï�i�� ���
B�ir`!%vɶ熂27�n���Ɖ�#��G�7'��ݸs��!r6��L�'�дj�ԣ&l��0�S�2rE�f��Ҿh�]^���\�/�nbu#r�ܾ��_�l5j���튊.���|Ge�ca�d�L^�׻�+2}��x����슊|����s[��A	���4��Z��F-��$
�l���7���8�l�\��1;���yR9���=R�r+46�'[*���By��>V���/א���V��ǡ�^����R����'���n�^�N�ݰ˴Z��u v�������C���8���dSJҶv�E[��8F��$h�RR�J��ť5,��#�.���aw�d��kb�w������}29�3��)b��nͭ#_��`Ѹۜ�� 5)�(�1���&]1��bl��D����6�_�))��$�C�s��B�����R�]����Y4L^x"�T��Le�&"d%:�I1��ud�T 6@ɿ���FN:=dz�@��􆜑~�N6�� X�^m�yX�A�fT�ڑ{�4P/&��׍��!��Y���.c~ynoW@����B@a�5��LX�F�ŋ4<�9�m��=3dA&�b�A��LnUک��w�R�{�)�L�ą�K���"�cC�2��!8��g>��c�53��i�lobqe���"{"0����bA��7���phh��F{e��
n~��^Xq��\��߹�?y�y�n�Wʫd
M;� ��g�yp?Jդ��|�j��|N�1���!c``H����|��ߗ^n���ڐ�rp����O<�s�����͛�����vm�r�*jٰ����K�ڡC�8<>���~��.�����g�g�<��\��D���%��7�/���x�|�(fj������������Ҩ^�1���2�M�F$�7~����
�ɛX"Z�[9�2�X��ҕ��7���q��5ģQ=�U �x�i<��3�m�����		H|����G�BggB-�L�m�~�o}��v�$�D$���%���V�ۖ4u��ǃ���?���)yL��L�cm{v���0�a�7̎�BL7Mr#	��́`\�����`>n������h
IN�=��#F�9T�Q�7�js��za愜!l��Y'���f�m�`j0�ʅh ��H7n�|�G����%HRd�`�p�%�Y(��f�%e�¯��3��V9�Fa����|�W���sG~N6_�_�����7���LtۼQ9DMF�V^;>t�>���08؅�S�W��oq��|�"ݨ�*5.�����=�q����bki'ũcGEW���*�Op�&�U����񛷥!����a@�T���n�8iN�a�_X�aC�+�,��˲�L�݁�ߖ�B�E� �l ��z��̧$�~bjv���W����HD���"r�Q�O�P>�h<�9�z뭷�+�p��1�1)�Z�����b���$��,�t��#,���!�����Ԭ3JJŁA�����W/����2L� { �O�CG� s�r>�M���9���Ϥ� ��/�;���s�B	V�,����h30�ԊS��B�g�!u��喀���@3a��q|���Bl�i���tJ��5M�<`|�
Ѐ�0�L��.2���s!�tI0�L�`@pl�t�b^23�x0��-� �T�:Rْ��^�^�V:/SB�ӎ�xP��� �Z]hAV	@2��,��&qej�H�4��t5D+Z���ZY�W~�݉8�:B�����2�����˫k��	�T�-���NFWN= �wM���Z�ݘ�z� g0�7 [6����4��7[�d� S+�W�y8re�I ���Tq���I
"&��Ѧ9��d[�n���&yj���ǩ#C����4Y�X����w��ʉ��H~��!�Fw�)�����5�WӸy{	{���6�z��BmڄN�
ŪhWC������#���H�#vH�mC���Ε�%��d3��U��.ac')����^�&���l��ڀ��eʹ�����X��V��G��Ƃ6�G� ��drH����*�n�I(U�ER�!��D<�p�%�"��
{XX[�l�n��
��{0���'�q*==G��v�*�T���aG���a7�������iwV��ۘ�����4�qy_x��x�w����L�cquS(C�`�b4��*e�|1�vF�8qd�	7jzS�|����W1qkْ�'(����S�/���6�l3:��I�p@���ĭ\�:+�)nr(�:{x��B�G�'~&�x��MḼ����}Jo�@'�=B�%~l D�HiY�S�>l(3���Rn�֥���j���g�yh6C��1����P�_X�̣��tI�ު�{1>�-~S3�`�'��|�!�'�,0���%\{ɱI�R �ۍw��ҲcC��� y�%�r%�-	��ɭh[�d��!	Aj �麨V�m7<���
Z<O�ux@�����tx�x�0���Z��T6���M�R)ih��vwS��:lv���0Cx�6��A�[4�tVJ��˧aW�L����"R�y��r��m��-i��!
b=^�4"���=��U�"M��(c�����>n߾-�gJ���pX��!�o(�=r��s��˫�X\\��Դ4��NJؚ�)��Pȇ��.><����������<��{�m .:@ {'ER�DK�E�r/��L���dw���nf����8���;��[�eYV�,Q"%�^  :n��}���}A���svN���s$�p�}���-��y��vX`7١��pSL0;?_�i�dL��+�������7�~W��7`�V��G�����Ï�'[��O��ӿ�-ܡf�{�}ػgBV��[-��p��udstv�J�/���ׇ��� o=&�N��
}���}�Q|��F�X��?�#�:u�l�<���򻧧.�n`zj����׏be%&o6�,r9��-��e��m��i��F���C}���M,bauE5�p[ �v?�6=�.J�|�,�;��H��k`m3 )�BZ�wUC�s�-[!O3����,�~=�O|�g�9Ai�ZC �~kT1�J��6�����t&�5UE���49��n]��į~�:~��W�J�3�dC���b��h�|6M�m����HlZkjم�=���?~�?��4��߾��S�����1y�Q�s}>K-aܷ�s�<�^{�M|�;���|�H&jک5`p����������~����s6���&�5���7��8S1��d/�}�s�Ai/%p{-M���J�S��\�$/�_�bh����ZDtf��	d�3h�@9	�$X���áC���|	]==�11����0�yi����b��=]�p�.��U!WL,�9y���y155%]lww'��x1[PU����Q;�.n����s�㴡�+�Gy����.�<)� �po&�ǵ�Q�����׏!��
Ҫ��Q)�hݸw���3�_��l�����-�kfJ�D6�p?^�����(��H-."9>���^T3�H�@��φ��G϶�8��� ۨ#Ỷ�I��S�)�����M�C�N������*Bojo�5腓i�Z�z��cX^\A���^l�t�;F{[H�<��"������i��q��L[wn����V�,��a�Z@d�b<�������a���_Kcq���R�bV������<��-2�"W;�Jcbj�3�P�^椫���f�������,��z�z�M�^;v篍Cos�����Jæ�|�xJ8������DkGX
N��n-����ނ�x�D�
�M�l��g����Ј$��j�&�"�[�w� |N�0����-�8s�&�^�M!C�����{��ju��g��㖧a:�����b�eR1�l4���<,�۬y�k�x�'y���p�oB/���I��RL�2�����[��5pct
�#O��tώ�c��m�f�L�������x��(�r0X�r���I�w����k�b�`0��U,��|�&Ƨ��0Za��Q.S�O��v`��GTj�\NL�,H،�8��=-�}pڬ���M�j<%Ġ��e�*Iu����[��Z^��͛z���$�8,Hkaj��s�$���H�Ӂd*�D*#Zv�ށD:�م%��m�B����z>�~���CR����|P�֐���y����n=\���J�2�JE&a��g��o �6c�`�4-f��Ê\��I�<7*�)��#��-�طm@<�l�Y��p��(�O,��s��)Nۍ&!gq+���]��pBh��t�;��>��f���b���`$�,�k��:�Ӏ��?�`q�
Ҍ�x,�|.#�dܹe=6u�Í���Z�pȧc�Z�R,�R�([1�t99����2%yl
��,��Fn��D�c�(�F���j��%�-Z;�)������X�M�5}�I�,�F�r	c^��F��N�_���=X�ւ--FT
bɄȧ
�<���P�Z"���d!�Mxlu��/	�s;rngRi,/3���fRɜH�n����4������d��sa��p��G� �BIDJ���g-�4���/�r��lK4��ccks$���N�v�i"�4��H�����3>�FGg�=������R�8qM�2@�G�@t�r3T�E΢���wpuxL|K��/�����4�a��}�� ^~��q��q�݇��}Z�^�J���:�.N�:�T6�C��'>�	X���p?���8��i>0ȕ�_��gg��≧~���/"K�\*�������>�Q�ݻO6�\Z\�:��|����ѷś�&q�gJ2)��u�����&7�fG�]��k����
0"�O"_�Cg�#�ꅯ�������EE�ae���ѐ���PD8�ܮ���
G�v����m�O������_�"�%Y�!���D0�Z��p���sF�aҌ�f��*�J�K�����E�Ջ�ז�Ϳ�1�9>���a�:œ��q؀����GC@�BSqv�������?����c*����#?{���=���u�Uy�M��Ղu|��b��~��<����^��J�P�ٝ��u����ۺ��_���	<p�0vm�3�d��ë\Y*&�kfܜ��wƤ!�ٚd
���v��'��5<GU�5|�Q߀�mA=�Dry���K�d�P˭BWM�VL�a�?0��|�#صg�|���E�R��&/��;�������h,,yp�!��#/�B!'�,���H�adl�O���p�ho	!����K��;�J�;(*h�I� \��/���^9�d�"aXd[�$s�Ύ��~ ����JW�'h���,��\���4 ��x\q��q�����ͣp��!P8��͠��E�ʉ���ZC�A�j0zT3�j�V'�fv땊�4x���چ;z ��J����Cƴ�=�E�()����5�c8��ʍY�~Z���=܄����fIN�ԋ���."��\	�ဠd�[C�,�т�Dg/�alv��Uѣ�I��|C_���,�8M��S2�p����x��SH��"��p{|� p�N�k:�c�Ⱥ�[eZ�I���@�R���<Fǧ�L��4_)��q0��n����֩$[`�;E �ڱa;qQh;n_`--��Q�Zuz���F���b�*+��]���b��B��=l�Y�v�����8��-Y�mN�,�JaWGW؋ݛ�	����CF\����W�P��Z{%'�
�:��	 �w���h�"�R��ѳ8��E���~)[+-$��!PS���qMC�1ӄ��I��l��A�`�&-)Spq$ި�.�S��sW0��"[��c�z��� f6�`ԕE;y+�S��DΆ���tf��m��k�&��QR{O����(`bN�[�s�����B�lTQ,�t�s�iԨ�%�dC�a�:d��8բ��K�'q��$*��fu��D�Q.ee�?��C��=Z�������0|^�55�0���l� ��T19����8T�j�BAҐ�U�-:��$f���F~��H����*�]�"�M4�W�fT�\S+(�3p��R���Aw[lf�ה�4pad�{�ȇ�M~��l�iž���p�f�|1�d'�]å�3�г`q�$^�Ɯ�����DL�4����R�+��o���"|t�{��FD�-�C{�ґ�ԗ+��9]n!M�j&���.�q��5AS2����m�qh�D��^4���d��K��<2��X���n1�k����y�3K��g6颁�ba�����q&r��H_�{q-�MJ5	!7���vC �Q�$`�_X����Y���jT�4)p�k�M]Ctj-N#��*�v�Ж
��4���@���L�I�a���Kp��9�s�� �ER�fff�P��4���JB�?Y�(p�E_��)��Y�!�����!�)!U�0�k�QRDZT���x&�>�2h��2A8%#Ԃ!_V�:�[6d�"Zd0r�����ٍ��	\��B9�P؏�&�8��jÎM[���'�"��ԋqu�$.���XVp��8���'0<6-�,R�L./�n�)e��|�cl�0��W�����w�×��%����,��;'q��)���L>�<� ��/�f�/��:~��pmxTR�+�4j_����/}Aҋ���8��),��I>T�V�?Є��G��c��@�<��Kx��/���R�H5����g?�q�޻�ro}W�_@�% Ԡb%/hӺZ��[sT�=D0��0)�zL2P�ץ�A�mk�}�!�<$�g�h���
�Oz���`�zQ���[�%c��.H��'h�[�� y�Nk��6`C m)�F�B�0	i��?�3\V7�:C롯7���zO>�<�f4�^�6 tˠ�y�Tl&��G�IÎ
eh�|䑃O~哏�ׇ����&��_}���_<�]��Qm.�4Peq��J.����A|�Gv걺��o~�^��J(�A�0���G���!����qkr�uw�C:��h}5 �Ɋ�yj
�Y�����E.5�1+d�J�/u�l�	������H��=�9��ƠdW`��_G�)�-5�������؍��Rٸ�y�twvb��mp9�+jF�N��%��� �̈�v�4�*z��������Sr��ChmcrlW/^���}�܍�N�h�u��
ΜƯ�y�.�`%��7�O����h�k����0�ܘD<Q�8����/)=��U#֪q�4�x�R'��NQ�X�buz
j,!��$���,�i�&I�]�ZC �f>��i��7�D�Id�I�
�����{�!0�(4(2 ��;�r�/r�\hI�$�[�Va�D�@Dhg$�f�K~֚�.r�sK�|�V����;�zDjR�2���?we�t&/���,�t�=���qKک����!�C���W���A8ҁ��.�47�,��,�TY2�Ը�"��4�F�L���ctlF�����*�V=�A6�wJ�H�47D�����]Ǜ�OI��?�"�vJ��^�5�u�����P�W�p��A`��|^A��ex8������hAs��ф��e��Ob|��h�C֞�d�uu�����z�N
y"dPl�0����%)�t�:�z[�0�ĺ� 4�JCjE:���%}�jz;\L��4 �4�Ya��`!%�D�O&��JI|=\�:mF��6�����D�ߡ5A:�� jUZP(*�[����2V�I�9�=N��c}o����*���u������	�.fDUoԐˮ �d��wlA_���g#G~<Q��xWe*    IDAT�1��C5R�g�{��JN��a/tL"�qWH/��U.�����عm=�������[Ņk��y�@Q�6�mF�i�U���)��x0m۽FIF2������!��0	#{jv�G��Ӣ7{��9P&����zE6TNka�Mr�m@k��tK+)�Z����i���03��G�d.���*�^-���B{3ַEZ�vpU�G��������NH�:'�0����Chi��f�ߌL��c�.�&*UPaq��Pe�� !�N��Uy]��qᔸ"���6�߸�DT<_,"٨����َu��h�8�����A��BCW��!sV�l�Nn-6���S2�6!|���}[���C5��D�T���WnJC��q�i���b�I�+,>����"d�k��Kb��k���E~�,d9��3FH6U-���?�D�5,�y~ަ��t�C �7����7ZCE�����Z�F٥q��'0��X�y&ݯ�� �"��
�DA_ �]�v�}�F����{�5���sB���l�P_��w�bQ��Ή��Ɓ�ΈD.���Uԩ�2X��$���96/,f�bCj����|��->;j�,��P�yfp[Dꐃዒՠ�9��I�L��,��3�u�y\�aj��� �L!�� �N������8���	{�m�̎�l3�㵣V/��=�;v����	��f@B��3'�l���42�"&f����g/��T7����d������p�TH¢/�s�>�ǎ�'��g�*~�ۗj�����\��#�8��q���jlI��x�A|����v7~��/��s�����H�wQ��?����"ҙ~�̳xᥗQ̕Qa<�Zm���o�<��cطo�3���8v��z�)\�~]���C�җ����ӈ��i\��+�����%�I
ҕ o��]��Z��m����cA���|���|n3����6w��$ UkXgh?M��4���"a�}R�x������L�:7Ԣs�4��f�Ѐޠ��;u�L-F6��Q5!艠-4��o�x_�ۧ��Z�����mpka�N�	Tl�Mk�BI$�qv��|�˟����`�������g/����b�r��Z�/�ػk#���p��5�NNb�ƍ��G���N1t��c�t�:����+7G�/a`h ����ap#����`��}��g�v�N[L��UF�HZ�#�Zpu|o���|�
�3�1i4635���"��������� �"��3dE)�Qͬ �(�Js��4}:Tdr��F�� �{�^�{�]���2� a�r!��9U�f���!�!��\��x"!�/�f��a5;$`��9�/�N��]�����AM�¢d��y �}�.�v�DL�ȉ��O����\3�������"U�!�փ����c�֊�kD���/�#�����b4����\��O��n��y��e �jEi�����^�f����<b��$C�ܖ)�y״�lD�G�h1/��C�q��5�$#�՚�����!N4��h)��\M�I�#'g���:t�i�i��~���4�����Wp��9	�9x�4�L\)��'�-`|fc31����z�se���lj7���a��n!�XL��K,x�]��KWoHb���Co��!�:�bx��Ve���U��&F�����E*[����b��*J۷`��-"u��,�a���\�"�Q������U.�H!"]!�Oc�P�mְ݀]R�W���@u��p��u)�ns�y&��V�Hwu��f�Z ���gf1<>��ŘH`8���rh�qp���v�`�!��a|~��I�F��pꭖ�n®�}��l��a���hr�	���x��5dJX�~�1Q��TX3@j3M)�!�R��$2,�lx���pXL��]p��p8��;��@a4�Ɇb�&!X��X��9⮗��ƞ����T��崊�ct:�g�ca� ��J���upϡ����S�g@,���r�n�`5�ȶ�����=vA�R��τR5��UjZ��1LJ.��Adm�7���)[���U�<���(���80��:�~5�%�5�>��>(�o���E�V���� ��&��AscI�r&_��+7$8+���I��ʷ�%y�6`S�m�Eo�咦�^YI���IA�V������6���̔Y��MǱ��w�؂���I��ɩ�cs�x��i\�X���l3�&�4�X�;7���X-:�N��|GO��|4W��S&oܼ�P���BslNB���[׉��v��dB�*�ͫ�#hf��^��l��Gw((Ġb1��Mj�M09<Hd�ȗ��'��62)�ybt��~;܁��I��T1 S�E���lL��-nz���>]��A�T�\ �e)`Y��%	����L�e&�� �����4]�1A�� 0�hc�[iX�8��ɴTy��<�vH'�R�bת��U��%��8�+�(��V+hr��� ���P�U��U.+�)j0Ԍ�W�#;6�����w�!�][7bۆ��{��Ƥ�#���J*��3Ө[�*:,��"��ٹ�ヽ!�*RrZB<O����Bgw���&F.c��)Xem�@ο�+)1Ƭ�P��q���?@� �"�ŎhYA�4�jYd��o�c1�7܌��կ�����N�=��q��qXFX�FDZ[p`�l܈�p,F���VG�vZ�K�!(ab~���O�։p�[�o�'��Ãl:���q�%��
����h4jx��w��K�,6lَޞ.��/b��M�,. �\�R�`߁�x��'�7Z�~�_?��旅t����~᳟Ɨ��EdK��?��G�B1W��&�k"��?�ٵ����{�l����ַ����>�u��ԧ>�{����,��$�Vnaai�rV���R�lV�V�5nc-@;��AR��4�T/pj��'�qY�Q˯�h� ƭ���
�+<vE� �5����	�F���V�p~��� ;B(�k�P/9��֞��F�3ə+��/�^_D��aC�^DgJ��7�׎^E]���n:JY��}54dpɟӠ�I8�Zɠ�Z(?�ȝO|����i����=?��K�.���;ڠ3Q�a�G>����^x�E��������'?�!�`/Z���ҨR\���b�<p�A��<��[J�޻���A�|:�6ԉ�\;��	M��=��^C��7ɴ�:\-�Pk�v��r�@,�rX8r:̂�4	ư��Pz`V
(�o��^D��(�'�������V��䰣���'����< n'�<y�������s���%��7F���o���������dZK�t9PQ�_Y�j4*ɪ��I�7-�+��6˴cqi�8��GO���<�Ul�f��r}�7a��]0:}2垚[AMg����x�2������z���D=��Y���t�Eo� �����WQ_^�W4�Q�7�ZK-��V^+eN����pǃ�kA��|��vX2@�����^C`P(��x�Z����b}_����f�*����8m&d�u������;W��5B
�ɹ���
��H���������`]7C�X�8��������|i9�D*'>���>t47��)�^'I��	���)�K+1�����*�5�LmN���"1:v�vo���"ԤG2Z@*_�U����C:����-X�e�4!����1c��,и���bu��a�23՚�����m^���mp� c�S����)�y��E�Z��4��`w�{?���b)VXM�02=��sX�qC�09�z�-^��>�u�A�Ͱl�������x��e)�ހ&"��v��b�B�i>�xa�/�f,&+��<�p8A��%Xmӄr1+�xCt&!pXm��r�O�xk�;��앇�;�Ã��,�=}���"�@�R1�u�~�s����ü�T����E\�:��x	f�z�*?��P6�����1/F�ə\�2�|�*�D�ɈJ6.�����:)��Aob���R4�Sg��}n�d�N�u�b�f(�����m"_	5��T*ȧ��&㰚M�[����^c�K"s��
����*�!�5�Px�p��4Ў=�7 �Z���8C�N_��|f[ v�_��F�u]�J�ز�6n�ց>D�v�wч�̅������Dav4���Z,*������;�wkg;�cL�>q�"�o��h��hq��=W�m�#�ZA1EK��{�> �n'��: ����gp��E���8CD�֡!l������*t�����(���\�[����y)�MF��"�~�s���`uaJ��ͭ��8u���b8Y��Ch��Pt&1�k��<�k��K�d3�hkFGG�Hʦf�1��(?#	a�ru��5l<D&����FdN����L��X�	�H|Z%2���L)�j��i,��]Eq�t�$,,Y+#[*#Wִ�e	��&�,$��ߍ�®��11|��铰�뎽h���%�&O�nu����|"��K������f��!`Cύ<e��|����;=}w�q@R�o^>��ѳ�-��9�YBU�m%�פ��P�A�]�2���A�T+� R�%n#�ʊ��#�������׾���N�`\���7�b~iZ��`�	�6n���m���C0�f	��JPaz�J�B�|����_��Is��&yR�N�[�����g?�>���1���N�;?�1b94�u���Oe�YI �����I|���η��т_<�~��066!�S�z�M:|����t
?��S8v�42)n��y<P+���{������n����w�7XZY�y?��.8�F��sP@	p�RK�E��W�H'�/���s�cEMGJd	����0�V=2�l�6d=p�3��/@	1�^�2����NiYK�L(h
H�U��D��h�1���B �$�&��+���F����vj6�1#��m�{԰���@�v�y���o�?��Q��F�-n(�f��R\��󆀞�j��b�C���W>s��`��������ٳ߿5��>��ٍ��G��o}�{x�wG��7a]O'؉��v�]b�
�]�B4jF4�Ə�4�9<���~`PX�&���PL�:��5�x���l`i�a-�Q�Uu�CR���$�I�bQ{�B�VT>�Jv�~7)4U�D�ƲL>fǯa��48E�(]:-�ڵ��>���$^|�E����b���C����;q�}���r���w���c���hk�ȃ����N~��5�D&!���6��^U��eF~:�%��F����M�FT��W4�xL1ٰ�ni
��{s�
U6��S
;���YX3��͔ɪ��f��>��L)�P�I}��*&�_��J}u�m���������5�5�4�1��C"4U��`���)�P�\�W���#�ݚɕ�T�e*�'ΰ ���k� %=m���h�8����DF�	|4���|%��"t���(&oŐf�Q�꤀tX�����+yD�.��@OW���4C����f�X^��������!�^>N��ʠ&J{FL�.bv�dRLNXln(��T��`p���mEW�I&K�XU�i�M�g/������J\�P���mX^]�j�����ZqTfHW]��79��>�4[f�*䟽���uc ���r:)h��LV+�'�q��,�&� �44���؉�f�a�+We�2<qK���:i
F�x����D[�~]�lt�Q�)��ur���|� �!MB��q
�BF[k�D6���R�eBKEW$ѵ�w֨I�*`��d�\���u�&N��}]a�t�ć���Q�\�>���/ciyU���K�4Љ��6��9 ��b��J���Gp��)6.��X�
��ހ={���-�T��	�~�,n-Ť�qح(���j�����l��9T� Y$����qsbN<DLj�ё��)�tj-�.l۰m��}��[/�`ZK��a��X�I3p��5)���&�%��bF-3D�Q��m��C��l��e�89=��g�bx���^�/*�JI4�j�&��}۶��퀩Q��b�pĺ����$�<yc��pxCp9=(�pJ�����]��a��^@i1bnq	箌��M��8`��&ic��𺥡�R��g>ý�����/�Z^cD�}�4%�v�����҂��6��0�k��`&S���FFnAU9Qf�Kdz����l®��2��p��9,��Wf���3�_M��jt�{͆@t�hC�V3q��nۺ���XX.��눧3b�%���z}�\�7�L�g���[�n�I�X����U :i���<�}Fm�I�^��U�Of'`(&�_�A%����_SAe�R^K/�P��P�eii���z�A�ޱs��x�g?F!þ�[1��'^'N���l��ï3=���xK�,R�:bI,F�"1������u���j�"��-�v n���J���j���) [=_��t�X��T咖��T`3}'D^+
J'�5�RY��+�c����������8x�a�s\�.T��x�	c���Է	�P|,z��q�3LA.G<��P�B�82����BEo��D���r4)�j�����9���gç>�0��{�wx�����/��(
�<X�4*TJIɤ������׿.r�g�{�z�\^-���b��~���g���
�����ɳ�V5�����<���A1C����0>�ǰw�.��N��g�����G>�A���b~qzSu�;TmT�Χ1���X2&$���6؝v��E��::�[�)(�2��j���\ߒ�I?$��!n��<n-V��>�u�\�uŢ?��%��������e�p�()�uɦbc-�m��-׃�~ �׌�y�4�ZF���ܰ�c���e3:}���~���Ë�,fkB]1�nk��9��D�?��v6�J���<�o>��PC�w����|anu����{6��C�`��ܚYē?��h�9�t{����۷`]{��:e��v�5�?XU�I���1<x�Cضu�pQ��`�K>+5d��ks�!X�ՠ��a�:u7%Al�uB��g��d���2�J�Rf]^���R@l~��W��.��]� )GE�T�]�cϞ=B�x��$��\t⩜.��hq{���u�N�!1Hi���$y]��@�E��N�8�1B�J,�/cnn���+&'���bs�l���E��#��%ŀ��n�"�Pu4ff��$��h����5w�L��{h)���ee�V(1��m�IB����Go��{��=Բ�!�2�ְ��/ɐ���M��G�����.�)mp�n�{�~8#���!�M�5 5���I
0�>6�M���"��bY�֐ݭa�\vX�u	�bAϭob�ix}q@z%>�(dnW&gWK�`i��ϔp1�O�e�6��ٌ����8�6���xH���� ����|M�� ؈�3�Pd��^*��j"��xV�D�$q�Թ�l�`<���͂��0ښC��&ʔ�}��h�e�L�P)���у`ЇD*��6�� )�8="�J$�x��Y̯�`q�œCJ��QX��]X�.�� c�\O�:4����9:� &R2���5$�}��r�IܜZ���tV���s[H�#����6��+ ���Na�p���Q���E�F�A�Y*�e$hi������RR���
�D�y��/ѳ� ���-�j4���B:�g�l5x�z�v��܊`�.Iz�|n,G�8u�<.^�������9�����d�(���N]����8Q����ۣ���[�s{��ADS�_��q��0N_��L6'�M.�n���v�א5����?���(����RQD�H]�A�K�]zl�Fo�E�T4�qJ���9���<�=���	Asz0�d�V4��%Swkt���sK?z;�0�j(W��Z���ØY��h��$[_��2�>'z{:�*�
�N��Z^WA50�����c|.��P���,��ɨp6�w����r��F�����1�F�y���f�S��l�>�Ⱥ:Z����})YE&+�&�p��,�R�0��0�$lV4�U�i�SS��N&]�R7�j��V��	���bN��a'�o�BogMO�    IDAT^���;3�ɳ�F�.�`sd����1���I��E4�Y�fw�ڍ;��,���g%��Ave��IksJ��	���Lf1s�*�����Ќהn��]�Ezy��֝A���ʆ�ii�m�CI/ˆ@�ĥ!��V�tȗK"������
Ƶ9ģx���عu��c���?�č�������P��ܪh��0lr~�	dj
��ӋQ��.�LS��JU2b�	������!R�R����h������x��`�J�<U�ehztI�e(b�($*��
�7�\��مE\�>��7obfyV���o���=�L����I��|
��G��F�=��{�b��6!�x�>��6�I��t[U���$�T��k����������P.�٠��X,�dH-e���/��s�����Ͽ�_��e��>TUn�̣�cM���R�j�|��}���7����o^�/��-n����:]��bƟ��?ŧ�����Q�Rr����jE���U��R������%�r%���v`���h�'���/��ʧP��Q���$e0�{����(P�>Z�P�U$R1ijl�׈[��Y���b\�[E��L���!n'S�}2l%Q�>�/ZBa|>4�(�M��.M��O(���YN�iݠ�&�l��ƾ�fH���I���1���ч6�l��iބN��x� 0@Ͽ�����b�~8/*Uf��$��V6�A����ɮPL/��<����|����!������^;��R��im���߉?z� ���<I%7nB�7�j��Jӎ	�`]m\�:� ��TK�k ����ś��^@�ߌ����u� �jU��t�� [�����P���,�i��d���u�!�;�S5���s)Y�3��^��j-z�L�l�P�%��8���"�2��60z�HD��Er�A�/�Jo��,Hx�6������Q&�5񿩩Z(/:Ѭ��!��)�Q<�6�ml�;�����DĘ>#�:�� ӻ�j�#�!I���D:DD5�<,]M��<�Vƒ��N����5�$�Tu�0p�c� �Lcuq˳3Pb�����=ɐȿ�yQ4�(���ZL�x�^��0,!?��"
|����	W�Eqa���u_%c�r$�Æ�`���$=�M�niɅ�I�A60�(�ilt�*5A%.ǳ�ƙ[A4�󟞅���D*0rMHҒZ��iA$��;� <|X ��F�rr�@d�r��A�3��R�WO&QS���r�0l+[�����k�l@0�/M�N�	�z�%Ԍ�}��xQ�J�d
�L��P3����/_-������N_�]��o�uK�,~��H�1�\̠Z�	6���3kk( 2lJ��x��,�y��ӆ�21�����k��ZH
z�� ��+���f��X�H���"Lz��]*5������y�$ƍ�C�O��N*�ľ�Y��M��S���#DݴA�5 r��|��8	.�BB���{HJ��i�,�>���U��H�	f(dK�%������[���GxƵj5��\�*pk9!Z�T���'dM�#���C۱cKj����`P+n-�p��y�--�������a]W�'QU�V��[���k��R���l.��E��Ȇ؀��m �����ކ&za8��iF;�a�bY����8{i�*?#l6�ݥ�)9��ө�����&�$��js��\�1%�3����y�tvE�u�F��#�J#����M
�?�b�0<�h�o�U"�^A5�Ǒ�݅pЍL*
�ہ\���XR��<�LF|MAēix��D�m�zir�٤\#6��r���1<6��ފ*osru(q� ��mSI&�f�ր�I冉�%����[	���+�<��:,ܾ���׌;lG��%N��������\z�K08Q��~!��3�����bۮ=b�>w�*���ّ���Ĕ_��rI�-�)�v��v���L����L�g�4
ZF����<W�i��]��e�+�rl��`���Rl���[j��%i*���W���G?��~�#X�ہDto��"�&G1�ӎ};v�mwh0R|֊s�&r9�zT���f���-XZZB<��;�����Q/d���Bkg��
f�'P+���ej��i��,>9n�%qV�Zh7.y�t�a�a��P�V%�����q��y�����k��v<�ÌD&�w�ǋ��K���������@���*�)u�^HG�f$	1ٛ�.��~�s����g0���j!�Ɖ��A)WB��F{Њ����>��$Y}�~���`%]F:_B)S亁^�%�ri!�������o���^����J��%X�ZC���>��D���Sx��S�-����l�Zn�j(Y/�6U��F�ۿG}����,`�V �d~K47�rh�A��_��-GC� �:[`u�-�a��V�e��I����C7!Hմk�9<����Fx]n�<�B���d^_M.�N�ȅ�����-�����JA� 2J�(i���5�����3�:�o��KJ��d�S,p���ڀ��8sz
��o~��9nH]�����2����\������)�T<r��'��˟������	��_ki���211a�_�|���\�+�����������E��:�0)��ڧgՊ<����,<�v#�mb|���sϭ �)J�#����QJt�#F;
������Y�؜�5ê����W��!�Z �/���"2L����RD����C)��B�h�ULܸ����~��F��
�v�)M"�_�� ��&T�L��ɦ�]/C�Jfh89a�ՁwmK����f��)�,<��D����U�X��8'/�2`s�� Y�PK�F�$gs�#���QB�Dg �_#���g��bQ*o͸,���Z~�WT��]�!1?���P/��/�h7��bN�9!�x|�sڱ��>�8|t^V�y�(Z�Ь2��S(��9�G,�J�	Wn4☌2��V V���Do���.�	�r���Ax�L'ҹ��a�$
�\��|T��Ē� ޔN�@6�U�ߨ��PUbwb����2�߄;����˚(�5��FCb��%�r��{�S�t�(M��bL�Œ":h��O��bѕe�l�@������D�"2�d2!��j��	=.�
) 
��"I	3���8VSYxB��9���,j�4�J��o�6lܲ~�z��I1��بq���6 N���f���㝓�MW`uQl5�?C����[7u�����rb�BY'\��7����㚱�4�
=E�Z�߻��FLT�tr��;Ԕj1�Zc���?�QWE��V���L�Ђ�T��7�u�*yX�5�6c���t����\B�^-<b���!/>��&�l5c5U�)���Fg���aF �'��$3o�Ѝ�C=���(f�rM�+
�FfW��e%���5,�7&���N��.�,6�5����^��$Bs%N�4�>�m�䷷��a��\m�c�Faܗ�����3W02qWL6��e�	2_/�WnpQ�JQ�����M5I]��5���fB*����"��q����E�3��|]F����쉷�Fbvi	7'g1��F"���h�n�eb�*�"\��ܻC��s(Vs��aѦ�Hk��y��3E��_k����$9�����p{�҄S
6���� �)��O��P�$�D�I�yC�ٮQM`Ҷ7"a�GP���8��p����l�I~W�4���=3����y�/ŰMJ�¿�v�%�v��.��TJ�
��0�{|��%"=}(2[�������4;m�d�5b�ךh�9�`�πSv��T��VihR	���
�sN%�&wC-�jb�Z�*�	�2iJE)�\�	�%��0&��c��G���=�t�.�}�t;6mD{W�l|Q�s�f�g�P�4P��*7͕��(2��q��2��|���(�cHD���BC��Q�'`pjC5�s �5ɉ���&���=�Ao�����yx��//���x�7�֩S�_��lݳv��F'Ν�ӿ�)斦io��m[�~6�5A���	ה'����1��09��:�����\��bt�������w�����?�>���(��x���/~��Ÿ��T��ެrKdD��D�Vl���ݍ@�	ӷ�$D���ⳌF������'����|�&�s/��e���X�h�\�(�m?��@>�Dk[�~��8|x�x(r��N��,��0�0+y:��Z8��fu� �u�IN�R0*P�*��5�$N6�Ź����/)bZuI���M������s�.��nc7k�ɬ���i��ÊJwI���^K�1���R��[�p�G;�!�����W���h����y._Z��~���dP�[G�O�wX�C��635�ej9�jf���G=�������93��_�|�?��6�eWS��)���|���.��N�u�u�C�s1���|�zK�*�����UBH��X]����4�͓�;���0�6nl>��_���(�v�^��'A"ٵA��P �<��R�����e3��<״�\�il�*v��<���0#[���U��E!]kxJ���hw��-:��pK�$`N��C�U�.��0��L��e�bܲ�Hf1Ia�Ɓ�����X)��r=� ]*A1���B��FX�!��4�5P,�u0��|�đ�� ِ�@�iDr!+b>��n�Ĉc����$�,����4��*���ↀ�71d�/��g�φ�Jɐń��ޅ=��i�b&�^C $��V���b!(��rzY����Y'r�֨�<������j�C=��w�Jpv�8�"��X��ϔ�A(zon|$���̆I�Z�m@I#�k�UT�s��u;	�7����b�B��,v�3��Z�t���vx�MBhᦢTQ�!��Y@2�	�V^L6OW�,Mt$��=(��qM�׮i`�VN+��ɔ!�6d�y�W�XM�̂��D�TC�\��K?
ѳ�_�aP�b�f7�i�f��ȯ�P�����N�[��Đ�OI���L�(����s�(v�m>(Fʣ�0�*�$��,����ÏP�)��U��a�RҖr�2�6����E˼#b��υ�x$����IC�Y�A�\�]^H?��tF�����4W("�a��}�!�9]r�i%z�&�z�)Ud��m�ӋE\�9���UD�UPI��}L�IMp��)2�a˺v���1��V���CMBӌ(I�jȔ�[/�ՁZ̀��e\�8�h��M���ԙ�K]8e2�����w���;vnD�$3�.J-U�(��z�_�1��O]����b���y&[s"����M�ZEKЍM�:���e�	��Ny��$��%�%4�Y�Y�~���f�H�v�{|�U+��gg163�h����U�F�	�LE-f`�)0�d}W�q]�n��eF6�o%>&	�
@O$-�������@ZH�D\66ަ����L�5_�V�l�x�ː�c�͙�+�u]�Ǆ���\U�Ar��g8�����|���9BFڴ~\V�H�L̝ ��`�b4���[��mIx-�l�GO'|^R�*�p�0='6X�>�pQjDj��x����$��g�������ֆS�]��������`H97Bl�J��L�l�2J�u��(�����(�,6��L�T��0>�����AoG��".�9�z6�ݛ7���]�F*'���|V�9��G�PC����̒��׌6$�E��)�<voۀ�����쪮E���ԩ;�A $$� ��c�ql���66����k����d2"#I		P��[�թr�:9�{ǘkW|����]���Vuu�9{��֜c�p��T�do:��L�7R��  YZK��s��:mrCR��	#]x_�F����W�P��q��Q|���߹�C�����Ძ�]�ܨ��G��}�,�.bp�[��(a��[020�T$)��R���	���L4�Ӌ%|��w�އ�֡aA�j��N�ky�@o��W��/��R���W��o��K9�;�k�e'�gֹ�vMZ4�htw��.��߇��U�K��V�Z�/��f�|�-b#0����A1ϳ�붮5�)!'�y�!�3�+y\|�y��׼����%k�Ad�8>��O�@�����|�`(�3��Zڷo�2�={w��R�!�,PC����|�h�k&#�4d���@\��sH��Q;	���i�` $Bܐ%k"N@�l5z�2���7�&�V@�C���Ջ�R(��U2�f;�p�����;r!�?1�~�N>��Mt�M�7��@83��!�3����6/�w�'��G/������_?!���]�~�����Gސؒ�"$����p�۱{� :��Ɗ��G�&�	4C���A2-_��]����J+�yZ�����S~�/�EPjt�&1�P�7��}r
ɞ��$m������~�Pov���刔�cفM��(���?�Qi�PЋ��E�S�@O=�8ٽ8���p��C��~S���LB�� �(~�|0."��Av�1-�@4�y�6c�	7���\|������rŒ�C��ڦD�@��Cr�c;v!38�XW/���
�z�>G�I�|.�Z��B������Ի���*�T�&PxJ�f܋3s��� �"��&oB`\�_�X���KطC��a�.~=�+^Rp�����3_xZ�����PD�)
p��(�@�/{_@c<b�ۓX��5D��þ�"d���16ҏ/:W���0��E��3_�0���Z�nD�wEQ�������Э%� �`)k�JǑJ�{�A�\A�X��ڊ�;�;w�ęg�EWO��C6LDeNOLcjfAM�m~�RB�B���""VXy��7����ү����,�2�^,,�`e��we4k>��O�B'B�vn
z��kiR�j��4�{I��א�Ǳg����+ǂN<�T�uK�əe��A���Bj����c�0���4�ڹ�[��k]�+UL�,�#��T����E��,#�a�#��R*U���1�C�T��/��@)���D�n�� �0kN*���fӏj���"eӞG�^P�pO<�g_v9�{���RXJQ>kR��#�Vs�c���CǰRn(��k��'�PX\�Р�����Ͻ�
��1�[������P�D�H�v�@Z��ࡇ������
�z��P�h>��uk�;5��5�K/>]]�9�i�K�y��u���_���;4�H��F��Me��sE��Q��h[Fp�Y;d����T_�5�$�����%,��o�v$�|��l�j5DB$#)q��V��8��i�+���_�!�U�p��SA����0�ҡ\͕�:�̈́CZ��>�حTY�
�W�@��o�|��P����#���c*�c�^�q��4���=�9��x�Iu��}����s�#��Ѻ��"��G"TÖ�.��<$��K�twi��5�c%�Q��Z>��:`���'w����C��+��� U�Z�>M�Ho��uDg1;l¸g�[feK~<�9�����BH�yDku�=˚�H�`ڬ�Y�}r�]Ai�:�UĚe4
9��(�ٔ+�D|�r��
j۲m���|\��8c׈�~����,��½{q����Vf0}zB��&�g�&g�Pj�����q��Ќ�����0�}p�1\r�^\t�ػm��RFR�.Q*[�U4�g������3�v�h_�Ã�d�4����!����R3>9�o��'���~��-;��{\��g�P� _.�!�Ɲ_A����X?��8��@?{�0�?�L<�&�������/�F ��sE|�_���=�N�[9 ̋a�º���T��	�+_�䖗�}_�򝘚]V�&���I�b)T�uQ��8��u��tR��k�V�!�I;�w�^�ܹ[F�'籸X��bAZ:4�p�N�>j���c~a
O{����7�{�؂���X�. � �m�����iT�M�Lt�sV(�4�Ʈ�����-��uPiW�,���,=R���F�D؇0�L�f��ŹC�e"20�$iOʏյ5MX�|p�%l���lX�(L��"
p*��It%NФ?h*E���$x�=;    IDAT3�:5}�m8c�%x��)|�cw��x�e�hE����KVWc��ۄ�݄ ?_��W<�S�����s���X����~+���G�����n���ߘK%�{����W4�>&F(��(��hIK	������������ف[^�<�{~q�/�����Ϻ�[��{?y����|�Zl�s_�NLUˌ�IX��dKH��8�<��8�M#ZCݪ��*XTJ`j��5ڶM���V)���X$��t�v���ǱCG����y��˔/S�k�1܋�5zM�P�F3D�h������0�m��1Ca4��+1W�z�b�lX��G�=<��;���G����_�-���Ew����4��lz���r�j�,�Q��ksGB�N�	M:G�T���;uX^�	������Dym�]��#:�O<Z�����'P(�m.�'��|ޛ��b���y6�}�-���EI�^��^&�1��)W�FSv����D�D���(�������P��<����B%X�s�P��Hui]S�G����7����U,D�8Z�JKs�aAkF
��l��[���^��E��7���k)���_b����M1�+�h��S��曜h�tO��bll�#C���R�>M�����F .���CKU����)_�	^(��,�x������a�B��n��-�H&�[>77���YM\����
63���#h���,���<Ъ�ZE�<�yJ��29N����&u2�H\�;�� =����k��`����Xo�m��5��e,��\$�޹>[�?{PIǺ�������r+�4HD����e����޴@���ݦo��jk��C/�@4��?Lڮ����^ɪ@ٳ}W\r���%"Sh�Ȥ�Zi��bl���p��Je�ϸ4.��^���,��Ry�誔�N ��;���~��!���!�23Wŝ��f旐���i3\�����&`A?�&y�J����at���*рhr�!��I��5��I���g�S�B�M���)<��I	@��(ڝ r�
�nd�4�j�����zi�����k��3w����`d$f،��fgW�i�Po!ݝԳ��k(C"�����I84�t�H4� ��~��X�9��Ŵp�=Q�ׯ}�ɵw�ʖycM�B����I1�*�|t�;��b�����E�0g��dJK\���}��KE���q�}HT�'Q���	��
��h��'�v6�4-��g��T��:�''\+z��y��r�����D 5'Qq#���⌄�܏4����!���0/*���nz��x��W#��QX�S���O�/���lIw����J.���0`z���v�tE;vG&'Q#���Ș����d#�]8o�V�F����mx�}�q?�&Q+��E��P��|����ए{��9�ǰ`FcPߐH��\��%|���G�x�.���3�?�J	��xt����]_���i�{�Yؾ��#���8��$Z�G�F
F���7��?�Ǟ�­�~r�~b��,l�)�6�KS�>�����<�9W������{���;����U*t�4ې}R#E���HS���t
�v�/hw*���)܍�s���hu���W��k����J�!N�S���i<��k�xF�����a,���i��)bfi�(C�"	s��ҠK�R���k۶1�¼�YMF�4I��3ò�H�V���[�xJFV��c2q"�fneiYuid�D��>�,v~��E�0s�se��:�?��Ʊ:�V��݈`2!%֝�~2͛�>JR��X�}��8s��x��Sx߿'OP���K9�$��R����_�Sɦ���k��W��E���W��^}v��o�l��ߺ!���̻�?x��C��/��#8��~�L̠;��8��,!ߪ��fD�NA���l5+���n�
��W��[��_��6�+.��#;Qo0��iߐg�F��C#���d���>L�5�ي@4m�nr���ۑ@�OT����ʃ��,u87[Y��jS�j�R��A�� &���o�0:FW(e�8r� �<���(4�U�FQ|7n DU��|�8�Q.zң���+VE{a��!E��0gdr�;@���!l=��lA ����
�W�*��Lҟ���ܺe���Wy&��V���g�!�5�k`�į��8���	��-D�����)̟:���,|�\�\u~7K*�]�����j�f��ˣ�G�Qv�D�̵�<M.H^��(��q����Y/|��S��(�\H�����vGw��R��L��ZMt+�Ѷ�vݎ���Ƚ�겙 ���������MFu�
��	?x}i�G��l��_�͠�
xE(@$B�9�$�;��<�nb�#�(�C#�~�a��Ƈ�M��!*�ü���9΂���������'�Tʇ�l�؏ɩY�3�Ʋ!3��o}��b���Z��J���,{5>W~Dšg���KMEV.�S�`���#�8�3JNKI�~J5��$"A��t���p���ȗ+B�#Q�s*���^�{kٳo��z��oBn�zIk�~�΢T�+�s��Y
�/d�G�ߓ��F}��z�euH���+zݬ�ff0;��r<���V�

>l�]�i��B�{4J��v��
��Q H�b�Q'����c�g���&��lie�E�tsb8�z��Sۉ>1M�<�$���F14Ч"�rww7��'~�q�i�b����	�[]7ڮF¦C��)ãx��!�am�aRM�kei�R	
񍖢�,z|���p�z�\�s�X\^��V(��Xh�k���B*�h�L��P?
���%z�Uc�������4]]=�Jw�ȣ��t8"��(p��
���abzQ���$��қ��� ��xM������6��g��5h��Zm�f��c#����Y�v�����RQ�O:+��\�4`���P*��G������R�%ŏ�;�?W󦡙�Ϛ�4����:s6�ux���+�I_��_�]v���޹����h�_~ťi,O�DquA�2�P@��+X0�"�F��7�`2f?�Zu�?��?���q�jUlK��5�F-�&2M�� V;>�ZXi�pbf�,OJ��tm�]�v]�r��q��b�N�@���yg�Ǝ�ў�����V�ҍ��>��/�������N̓IT�ŒXk�q|y��?����ĹO&���wa��]�����������/k�u���c��]�P����;���QW��Ъ����Gw �=�pt�sY��c_�w~� *����C	�VZ���Ǟm��m������Kw�_�&��
:C(�%r���M��e҈��₾IﬖVѕ��}��%/�'��w��>��[XY��i	m�n�)�r�kK�I{�v����<��k�淾[��bbn�jZ����;���)��@�+�`��y�����M�R��NQ��q���_�d�P��ɰw�s���5�@"F�v�� z�z�5�=tmqqݎ��#����	Hq�6z&��s-�eC@#�H(3���6Z	II�F��H �X0	3�d�Q��\��<�~�K89YD�у�?�N����݅*����r��l�y��_�ꗿ��������[5����}���u߁Coݱ��ƛ��+݋;>N<y�==��"h���*83�P ���jL���K�v�=�R��w_������]�-��ܳ/���Ս�X'��V��$����ů��+>5�D�.�
-�NZV�I�Q�������B2�Kk�RUa:��'�A$�X�Z߷V�h�50<Ѝ�L7��Nڏ���xh 
0k9��(|$7���l���7���)��nK�3(8.� 7�t�]=�����g"��'�A���J��2�1�	�É����{���R�u�z��F��դ�!��+t
l��$���Cvy	s'N"w�4���Q,�����M��E�¦�h��G�+RGQ���@�=��`�a�m�\z�5������&��a���6<Є����tX���+�y]]� 	�|�M��tB�:���X!��
G�|}� �F�R���g�]�r�,ʴ�؄IX�`9���0$��M��ZԄ����j�/�YD�y�xp�@�3V��I�D�גMU�]r2�I�#�?S5~�(f�14<f(!�$�U�5�]�&N��cG���y%NxH��R��U���p2��>lj��Tij�|�Yҟ���
+"��s���W.&V�(�^k( _��A���gh�v#^�G^'�v�mt!7p�Ŝ�|*�%�tk���x>ּ�j��T���o��m���<��6�H��֝Cq�����D��AD�)M�x��Y�r���V�̄�h�(4SR����J&tٴ�n��Q��~�����~2��b�IoBE����d����N�V*�eu+*�\�8)�h���A��Ҋ�P�:P;@��E��+�Q�$����6�G��g�V4[L�>����L:�]�v`xhH��ם�ܫJ�V��8��8N�:�`��}F����p=ЕJ�p�n�AK-�rE�n~uk�sx��/�uϾJ����8uZ[��]{1<���k�5Qz�s�����CU���U��}\�v����4\\o����o�������� ���<-:�U����;�{�,m���i�\�>�:�Y��0���O��%N��T�B�٦?$�)�nL+��C��܊�i�KQ %��x��F�ͻ�?��g��:5�|N�E5�1 \Y���8�OAiuyݵ��L��,������՝V*�u�\����Ï=���Q��@�Q�h,��d������<�/�"( �'�X����-"W��fD][��@��^Z��S8k���vcejkN�q�Ȁ��,���2���A�X�󓈧�n�ĢN#�G�֭�j�0&y�/gql5��bWߴo��D��&�p��������v��[�� !�L`��GYt:Z���$/��``p��#H����b	�����z#��w*5,�>�s��߽�Op�U�cvn���W�;���S������o�y瞍�5|���Ɖ�	��J��6��֩��K��߼�-��Y�����]?��?�q><�f3�r��)w��<�1'0���4�f5���q�M�ƛ���غ���Ǳ�:�N������)�,�e�!���^�����F'�S�F<��8�ⴈ�3C]5��Yn�����.�uL�u ���aզ�SZ[XR��6#-ȧ�1W(�P*��3Hx�I��$���sȥ|�X�u��U8��TE��-�)����!#�p�n���r<��c�Ї��S�e�Їv+!�.;g�׭7!^SN@�!������/��?��[>p����߰���[5?}���{?�xrr�5O�����_�bLO��}��>,�ߘ�^RX�����D��̍�*�d�2˂���L"$���{>����G��#���kg�9K�7����#�[�A�R@��W�� �L0݂P*#�o�]XR��.d�n�
p*�k��=�8)ЩqL��hG�~Y��S�A�T;Uu�݉��r.X�9������x}ٕYTJY���	����ǝ���,$����X(�F��G�A$ҽ�CW� ��nDI��81=�%�:�[�P�L���QX<P����m'U��Wo^6�6���)F���5Cb�S�J�=1�����5i۵�H\���F�-���6���98�{�r":�}������7\��=�F�2)�
(Ӊ�\C���!�l�q�ǃ�cwE�
[�at(+\YX��d���ȭ��C�Uԓ�E�0���II�����ݐ��/*�SE�9��J��9Nn��t9����Q�ń��p]���@2��ь�z�\�?����(�
��lB[��P�|6'��K)�t��J��?����b㵩!PQV��o��,���LN���p��b��F����p��}�z�C����M�jU�a~��E�$ø8L�U�])�D$�?K�ݽ�!�����ϙ�!`���l��@��bS�.d�RǾ���r��1��^�MMCh������W��PXNI�a�S*W�8���4Z�A�\@��s&�x"���ɉ�դ�D�Q,���6"0�M$q�^C��l*V���!�V*�xe���zPφ���f�� ���J��!�5��0
�E��{E]����r)���y���s�v\t���A�R�m�Z6���
]��g��0�"�N"���&��k0��8�2i LG�BI]$k���9&�c�<���%�����H���|aU߫X��JsqeU6�1�q����0q��W�"8����~{���͵��Ok�t#]1���'�����L2��=�v
#�P*���ī�D�����2��Di���Dj_!6���GU��ܢ���66]�M<�'f�����(���O��n��Y�̈́�
�(C}q�s�p��QZ���9����5�5ņ`yyQSXNڸ?��9���Г�a��A�?���<��1�&��Z�f�(�r�6�ҜpB�X�`�,��X�=n�fU��t�|H��K�q�9g�9�|�2]�<~sǏ��4�P��&�m��L6�	�(�j!��h��K�6����j>�D� 
`b-���U�q�K�y��=��O�Tex�y�O�Rn	�D]}�##�/ӥ �z!���U%�!��2D��3pj���}�s��g���8�����q6Z�"r�'q�����<��gcnv�ꋸ��w��=�N�%/�	���W`���8p� >���p�}��Q)��4��M7]�w���18E��ƽ������ؿ���Mu��&z�����`��F��F��*n��9x�_�[��cf���f��S�U�R\����V�e�@�fp��V|F��04؋�~Kv'�����P]Cs�.�ӝ?rVc�I�P���^�h`S�+,,�\D�&p�Kӳ3����Q�@)�*x�=��s�#�}f��Jd����C4�@,ЅLl];q���q�Ç?�U��� ��C�F�B�R�hT/M��Il�Y̡�6]x�k_��7��-��ߢ!��/���g?��f8��}��\y�ex��'�o�ފ���hJ#�D0�/�7�\��z	�=	\q����׿
go��B��{�� ��{���b���J�&��f�<5�;��fWۈ�FIuK�/��g�E�A�Ad�;�y0D������榧���hM�QdW��H*�
��Z� �'@2B<�F�W��#�@�f	�FY�`��
ْ4L��IZWN�<�3���])t��#�A�XE<�_0��M(�nw0���R�j<�5����
��ӁFug�`U�FC���졾B���-���O鐤t�rY	 �^�NG��I�i�7~N����[���J�)y�8"��J6鈎dC�bZ!����o��P���?z�"�憀c^wL2V��ߞ��C�77:���خ�E��B�beM�Dx|�u=n�0�j�jU������}�)���h>��Z7gY���7�B��p��95 ��)�������(&�*��r��i���H0��	��lb\+�t�F��_ȷ����H�`���c��H'�I�j��me}� �,�u ��P +ĕ!�Qؼv��z��dQ�5�j�_�M��D�r����5�,���r���=�b�*��G�����A������}�~�4$v��Z�+�c䡛nAt�-NmBTo�T�3���޵�O^Q)�g(ײ�ȯ��D�H!!6�	)j6��>wZ�.���{�uR)�^g2,��vm鶢��=�z|f%�5�A���Z&��G����
ͺ�N۷o��m�����氼�,���0���.{�M��0j""�k�y-��d��
�n��ygSI=Cw]S"(���>i�+M�>�Fe����g����8i�z#h����Z��P�c91,�]��@k��A���;1��(��~�|~?�S%M��A�)N�lrM`���׈�SN��E�W�Jk��/V��Yl4-��h��f��+N��Y#Q�%�('���MSb!�F�uBM�}A6%L�f^�p&��HSO>�����gA�    IDAT�"���A�R	Q�<�pf0��k�b��;��*9���]Fuy	����+@�t!	�2��I���c�PD%��|����2��F��W�Tfʢ�ר�?W *-H����..������c�S*��b��!q�9�6��\`n�")¶���<K��Eb���J��㫫�(�I�����O��z��Q?�ӳӘ^��Z��P<�toc���đ�aAH������36	!�B��6��<�S�x�Ǿ�_>z�U�<��p����4ιd7�����q!����2���_��R��܋w��_����?������|�'h�\�Ą�eUE쳮��~�;q���n���?��?�Y8p�F��x��J�}S�����"��ny��ַ�1������r�@��R����i�:�٥	����
t�wޤ�R�}�`tl#��2����t�&���n�`gO`N.�+��3�p\���3�@����`H΁j��1M
r�&gg4)�B��HI��<�7��Rꮅ��63���0��A�݉At�GћŮ��q�7���?�MLΒ؏v;�L����࡮�{S`���Gem���/{����wny��������С�|�+oٲg�?��������y|��_é��ǰR(�Az��3��}oF�FMt_���ع}ox��a�7���"� �6v��k�B���� @���0�,��=��3%�C*��<,ĩ5�@6<K��%�F)�mӬ+���֛��mሉ.�x����!'��Q�o>oRF��i+�5�Qǎ-��>6�x4$����
*%&�$2eB"���(�!2�[)��a%�����rE�䊨4Zu�}&L�k�R^E+��9&%��r(b2��1��b��w qC!UGŤs�oM�������%�Q��r4Ŕ�F3Ǐb���&�e�nN>C��{c��"N�EK��Ԓ��.��֡��RC@��,�g<�\r�5�D����5!൐�P��͙{ D!X�7�K�����¢B�̡��f��󺒲So�(�}��+ҽ`�JdFW�g>gŴU�j|<+W�oU�q-̊O5�,��TE�������\��ϯ7l"\��'���סx,��*��L[E6���Ԫ�oQ#���I��F62r��F��"�!�}���#�m��Ǎ�-��CU��#킩�F������MK����o�gs���G�5��xY�q�z����1^a�{�5�|���΍�g�+��l8oy�A�4"�<��l�5g��fg�R"���R�6����5�,,i_�&#P6	ך�� =������J��=)S�#7�QԞF�_v�ɻl���E�*�u��.�F�^�YZz}z��3�=�Q`�xoǗ�4�_�u)޹L	̉̚G�"�U��{��9~=�/�;)#ٵ5��e��|��s"��1��0�="�^�&O�/��X�aɻ\�jl�ia��Vg�YG	ȥJ�٬l�I7���'�e�{��B�B�5z�8���eMAM�l(�P�E��f�mk�>멚=��[�xI�I!�@�H���|�糺6�PTS��!���(�Kj���A]������'v��I�U�l�k.w��Mx���%n�p ��DN���׉����ԡIA|����8FR!�:��=� ���&���kNg2�^�s�j[FG�m���r1�L,��߇`���C��K(.-�������2��η*��P3ky��K�<B3	��+�H��XE_*&mƥ矋K/8O�Vav'}��e}R;�,1�L4�zC�n�_>+<#8=$�W����Qqzu㴭q鳯�஝�DX���ajn+���n��?͆���~�AQ�#о�3%E�#���щe|��_���h��h7�R>B�T�q�E���s\��˱������K��GnC)[@��1���ߌ}�����8=�O��%|��w�U���lƫ(�06ڇw��x�+n�)��s|�C��C=��Z��pW����0S��k+���,^��}x�_�	�]C�-,�m��`���8|�����Ѫ�Ź�"6Y� 	c��Ai	��ϯ
����Z��Q�%�.�-�z�l;����<��aR��QR�X�xRzR1W�VU�؄�E��w&����0�ܐ�B�^'�'�ƹsm���ۦ��CW��]��M��7�[��⋟�>��ocn�,�^�|� '5Y�p
O��3q�D��N��ja����_�����+����4����o�}�Y���HZ���	��f��̯�D�	���C
�U�HHH`�DӀ���ɎG�����64x�WM�W3AkN����>��ǗN!�;�Z����<���:I�g
.�34�!N�]q�]��_�XR��n�RN��N�I~?�����}Q F�Bک���}�N���W��d��[��eU#b�6�DW�###�?����!6�H/_z�7��ۏѱmBh(Z���P'��*�d�6�d�P���	iZը9�$LyOE�_�2��|��Fk��b�b	��:���G]0Y��f'�k�ߚ�'��ϊt�D�Xs<�]O�5�s1�
��!�������E�����I�Qf�_�e
Qr�1|�U��G� �8���D����RO�z���ib��
��i(�-�8z븷^C`�]_o���gZQ!�xt6$��R	
�q�^o���� yӤ��ζ�-�9������c����IRb��u@h��1g���<���fSs#�E��9;�h�6�F��^�Qq����t.�������9b���ʐ�����;S#a�՞Y��_)�<��  z�����(L�4k?pfq��,x^�����k��8pr�5�	{��$��n�p}y�6�l(��������1�t2�7_��rH��*ڣw�İ���0� ^G~��L��K���/��x��,��8�>,�Mxe����Х�&O���R�fM�K�鵜~Fn>	����u��O�	�]��]�M���"6�N����֦=�Ds��=7�8=	�&�!���h,([�b���oj4���p���hx�hB��/i-�Q��"�I^c�lKf.K^"��������%d�o#�A�I������!N��ӅǛR�P z���q?!�E�<!!P��"���֧�^�-g���UA�7�T�O�$�Sz���0x�)����iZhV�NE1�	a�G�x�����	��fW��<66&�%iiL���35D}y��5�ۍ8�r	}�4­���V���|��+[�H�X
��"��2�i5M��M3UQ�ɸ���x=�����8ꋫ���*U����n�
�r���\�h����?6���P0��b�TBm\����=:�R�)n{�P������!�9s�MheY�j*@`p��G5�4C� � �m;�N�㓟�:NN3�+%� �8�::Lj\[���Ļ��/p�uWb~~����/j2˽�����7��q�9{p��8>v�W��o� �]���V�}�^�����o�K�A��G������2�E���Xʄ���i�`���Tl.��5�����W�fl�1�م�ȗVI�P�����tȵ��Pa�W0�����cfG�-w��E0�C��l��,c�ܲ1Q��3O!��̀B� @ОMw����c]+ �K��X�f/Q����/3��ų��ҙ�s���q���� \<.��O�Pw��z]�s�h?�C�ڎ��.��|��o��wރ�K�9"����^�X�y���sA��k�������]��7�n߿^�s���������9�}�疛�B�!���|��V�1M�ָ���ؐ�OOx�xk먣\aQ�q���c�F�-�9kN"C� ��TB�^j��w=��O�"�Afp	Ry@��;�G.!s&	ț�I(+�r��Q������>=��o�(SAZ��Ŗ<�u�Y����Hr�Ѹvqnuژ�"(di��D(�A$f�-�zS3�ӭ�J��kD��(�VsH$�زu�>���,�[��3�5�,R-\�K^9�_���)�U�C{$�f���oX��{ra��B?�h��DŇ{X�Qm��H|��S�f�8��*�wϴG��k��A�?�l@�t��v��[���}���#�k���
��)��Q��]C�"ːP[#te�\�j��x��ZnT�!�^(�\s���G�QQ�Ę���%L��ZL������C
�I	P��cC�QsDGp\e���YA�5B2�����Y1&��RTD7�*�q�Ձ��k.A�T7)�M"�H��A8��:|�Fsה߇��Ffl��{?�H����e�!�Gi��Ī��U��P*��<k�"�Gs��L�|3���ǻf,��H�Mז�9�u�ֽǵ��s�v.�1�u#:��'���s��@���0J��
�����=19E���1���r�h0M;�C��k%��M!x��l�{��1i��Od��h��Q��i�t��ަ/�ӏ��?�R�L�f�VH �)Áhe�=�k�G�XP���_]c�B�BIk=�U��T��2Р&�j� �f���	n�jͿ�]{�Y@s_g�gSNF�i�v.�dkT��!X��꒛�oը�����11�G�}c����<`{I��N妆��F�snM�����5~_H9l� �w6BܜI��G�l*f�䛨�׍Y(�Je'A�h;�L+��e�ד�ܴFD�i�D��$�sj�T͛{�=SrY2Z%�%�\�����0�c��cUWq��?�]��&|B����!=7,��IJ!�B��}��0��������e!�[մ�;�S''�L��-2q�4b��k(�f�C|�n1�T�}<KHɡ�+]�H��dnJ�(;����#e�W�*Rn��k�iA:I��&��&|j��
{��j���YWc���X\]Q��T���y��s��>� ��7������Cz�*�8�I������sp��4>��/c�ԂB�X��~��`Ӈfv	g����o�7<SӋ���/�C�M�r�w�û��v\��+057�}�'p�w�&.jʹ��o�$���eϸ��߷b۶m��]��m��y� ��E�d���MRe
��]Zpj�n7Pɯ�E/�o�����]Ø^�@��G�'����8�(��<�jhZ��!J_200�Ɠ�m�VC>��C=�WFKem�Z�������(G��B�$z�	������d�jo�M{q������M���1��s����zE�
#E-" ���H16G��j4����@2ԧP�mCgcz<��o�~tϣh��ݛA���3�uS�~� ^<&�zN�Z�T\|���}൯��_=<���o4��>�[���;p���_���"���w�s�/>w72a+4�0:��a�6B2Lc�p c��܀9�c�?U����ӨV(��
!*���-��bxh�2��3?@�A��=�S
䍍p���7/����"P9D��p�g��
-Y�J� ����ƌ1�Z�l@\RV��ɫ��\��e8޹�Hؤ�@4��z+�ZӍq���M���Q�ǲ�b�̓��Y"�C4	��m��%|3���_.*N��f�E3���P,6���
�5�D����,!�q���:1��O�r�d�*��2|j��U��8r
0�łS<��`�B%�P
���C�MB�ᖛp�7�!89?����1�@�A�
)+��������^衟��U�+���;�km��si��0�o�w��%��MpD'q���Fz�**91p�g�soݸ�ڞ)ϓ���G������~kt����3ar�&>�hi��hx�,~?:%y�f3�˂X�I�(&�x�]�[{D�y��ɶ���~p��k���*y�(X�����!��g�='Q�::��B�bW����9|m�ł�C�u�h�����2��_�v�G�ژ*�B��ܴ�U����O�x��+e�I,:������y��C6��n�j4��lI�cS��Tq��!����ծ���9��[�B�~��K(�֥�j�_F�b#/�6�_�Q��\��a�lz]�=�5K�w�	��C� ��ߟ�Xd�z#�MUL�g���F=/�
�r��`p�����{��G�J�'���ߗ�rYr�@!�lD�sf2'�/���5lj�Dў�C^S#3���y�{k��FԪi�4�)���r�2l�.|O�sm�"l�,4l�����`Q�I�Lī���XT��i1�=�}��
8�#�/|�3�TA!��>��D�R�Z�`"�x���S�p�~��/�;Gp�=?���|�9�v����A����{�.��ӭ+���������έ�068�gg��i��q�����b�x��f�6�x�#��/כ&=��ɶ�%�qr�X3���¿��pfp�k�l��ISWBG$�oH��6�� �1<oXtrRV���c��ʫ���o|��&l&��<N�:���)�i�h0x��J9��عm���r���qhl�(C#{�����֏��Բ&����n��}m	{�ڊ��w��k.���
>��O�3_�2u�u�9c�W�<�:��E|�_��~x�&�����l�X�{�3�go�#�ڹ�����������P�uЪw$�U��I�M�T�8#��VE-���t���{�܉��I䊫@��|;����q|�8��5�y�h����appH{(����5T�E��`����t%P��P,��Ч{A�B8!��D�Y��C�j�z�:Y���H/�hr܇�3�k�\���"��@�����˟QmV�`W�j3�x���?��1�ret���OmEo|��F����w?����X��Ȇ�I��&��5Ά���7�Z	M^��j�կ���7��K��ߢ!`R�G���wN�/�����ܳ�e���(
�H���@�B�0�o�Lrƴ]-B��1��u����K�����S)�N�.��p��?{��𥟢܈�wlB���n�>"ТΚؕ`�_���_eH�G����.n��9���67���U��p9.B�t�n��F���]��F�<�;|a���������DBE1�c:������UW�=8z��Pc�c�C�W�J0��υ�Idl�j��x�L퇄T�Z��3��"R�҉��g�'1w�J��4��O�S���z���������W���T�h�78��'�M�i-�H 7��x�M�SCptrJ����CV(��B�C��x�펏�9
��c&:j�悑�Whڵ�{����1����a�d6�W��Z��v����Ԭ9�o��e�xv0�um�z]�P�
!�lQ�~��y�+{-V��pvBf:�z��^ʮ�&t�?\��]PD�e�	�HN�������S'B���2J��D�`gsO���$.�OAJ�מ�.�n��@d��� ��2�hs�����޽�i�P�`�jC����5�6��s��"Ͼ�M�4E�TN�M�6�'����(ɷ��b��"Ŏ��cff$� 1�	�י��deo8*S$�\G��sW�Ll.F].��k��>q�_ž�`�[��� �y�šw��|�t�=�ۃ�,��΀���Q����wUlcvp��akyX�&���P��)�I6$n��d�{�s�5s����&E��<�)L��v=w6��v�=���]�&1<m��D�,�5��u���ߢ��k�'f�e����/�f�(-���B�%6֜3���k�}Vw�5��� ���F��j��UыXs�?�й��E9�����}�4lL�h�(���i#Ѯ�S��MϺ/��*�EЪ5�|��v;��V�ަe4�>��b�^6is�Wq��8��fП����
���e���8]\YC�T��j&_3���#���N�.�4��%��E���H�MH�ʺIf�cP[4��Y��Q�X2�PH}��ղlO/{ڕx�o�Y�����,N�<���E"�"�fp+����AlU�����b�
n�u����C��/���&�6�Gf:Q��A�RG���Y�l����w�W]�ӓ3��G?�;���,u�.��3��y�[��Po61��G6_��BJs�h��� ≈�ώ�[�l-/�`qqUY!3��8q�R�]А����Y�FK�N�Å��X    IDAT��)\x��xӟ�	.}�EȕV����B=�l3���"f�f��]��ڂj^7NR؈r�fn���
����{咔N��,S�M*k�9 �)�F-�T/c�����x������7�8'=������5�v��)�����P�D�I�߯�c��M�?����3L��t��Ewl��1�$�!��7��1>��;Q�s���:6Ɣ�NZ���Yˎ��zi��B��/��}��×���##˛���ϿՄ���'>�����C6<28466b]��]~����XR	�%7,�]�'�C_�Z���۷��3�R0X8la����Ձ�:�;��(r� �#�ѕG��5:�Xa@�l�����fm��<D�a�DLC�x�P,�.�Rm�X�OvE�@D�Բ�QAb�'ȴBR����&�Q`U�
��X>�n��T����Һ�O�z�ʂ�,5.��P9g�����A/���%�isN/��	f<N������J�2uQ���'j	�OM`qr
��Y�U� �UC��$L{�ژ��Y�	��$5�Q��x(q�x�4B�"�3�5q�-/�57� �P'�gQ`:��.g��P;oZ��Fq�Įh�^u�D#�u��w����eC���Zw�q\h�ʎ��5^1m�Β�̽�k.HѰ�`�=[�&n���k(D�Y�Ys�>�I������5�ހ�Wn&�@�\^�ؽ�+������oI���H�Dj��@�u��U�(i 6^;��a�5��ă�E�����c����!�*�L=l��k�4�5��W�[A�A��6G�mW�{�'��O���E��K*F�V�v�y��>��������֐'uii����>����$ȡw?Ci��B�\�):���т��8)��4Q2@��*���,���OBZ�]������]�!G5���lE��q~�Ҙ�n��D�A4E��~�sS+�Ul"F�6�� �GZ���yϊ�{�5�^�Pj�j�L\8?p����`h�c�u���`sX�ЕXٹQ���kD��s�!��5ql"�;���	�i���o3 �k(��l�)�6*���sx�	�,k����p�V��I��D���ɣ�i�H^q�ϼ�97"�k'�_0��x ���7p�� 
�|y�>�l����MS��@��t�b�PXB��&Ͼ�U/���;�`]�>��~��89qچ��6r�sl61<�/��d,.
R�QG1_���6��������TWZ�2Ӯ�8p��xR�Q�hBAmN]�Ea��WMPt��/��M|�����2'q�:�{�rP�X�MM�����7��q�UWI5~�8�8�3����_�t��s3r�ZZZZ���À��.�������OM-�iaLM$���=�b`dx�)����1<~�$�u6�Y�p�0��T����?������1>~���K����#�-��c��~��;�/�w��"�� d�J�!>���;+���9��lE�ՆD��h��G,s���#�L��"�k�>�{��)��▗݌��4f�e7:���b~�˳X�-�P�"�=8D�O�=}���
�YX�C��G*���c�A��e�PO!�*uh�)��Vkב/Pbv�X�;�6L�7�4�q�4'h�9,�������Q(��'|&�{�ϡɃ�\����Q�E�/�x'��� 2�a�$��'�����;~���a4;q�~Bq�Cq�yt#=0Q�e0J��|t�[[@3;���W���?{ݫ?|�Xz�7m6��ߪ!8t�P������}�ɿ����C]\N?����)��Us@`�h�qs��q%�X:����i��|��/��z\xΙ���Y��I^ԁV�<qx����V(��B�w�pi���4VG�����\%���D�a����W�h���ڍHG����D��+�U���ud�z�+���=Nhˢ�e~�D�<7����&�0Z�-r�թlH8�0.7]�aԘ�hMJ�u"W+��� ׯS�C���uJ��W'��5Ug�ڕ�#I�)�W�6u�4�������g��'�^+jܨ���lY,ڤ��H�8��W�i��h�D���K�c?ο�\���Jc�TPCP+�D�b=���&pm�Hu�$�����ڨ�c���w�l#���:
oc��^H��?�^���@�7�V�xV��C�7�^C#�չ%yk�E��x��I։^t<��2y/�-��8{H�7�)�
_6V|����ikD�]�K���n6庡p�FU�!7�Q�!s&��i�H�4 j'�<t�gs����h���i<XXQH-�K�7���5���<]��(xMIXظ�3��#��o�缆`ݥ��2�����,G;No�Y��⏅��*%�	'b��[�[G�Yo��#�S"VܟxI�̺�3N��$JL�5��y�����6��haͲ5F�Tf��{ͨ�25�?k��{.�:�h�	=L���$��9��^�����,�-��U��֑7Y�A��P��B���Eٳ����]Zb�B��s����Ntnm��$�vS_�}pQ���}���#�{���7rqυ�<3��� �"�u�M���l�d�#���&�uq���$7�FǬ}7��o<���_S&�i���.�Lg���D����"�%�U���::��9���D�WKuD���(�_^�px�K�������S�Gp��8~��_bfv��V0�[�Hė7���\��dZ�6FFƴW�&��v�K��?ý���r�x� ���لќ^6B"��qN��%��+m4I�ؤČ7����I�H�4JEݟ��^���	����Us��'���&N��p�%�+E9jy�F�V��ر��{��mCW"��+�P�g�HB�}�c��C�����!<��(jM������hU[��r��3��\|�98t�(���o�{��)��i�0:փw����� �XP4�em3��go��)ڕ7A�\n�6��^�Ǧ�����_���p�ؓx��������N�fO`|������[R0Y+�B �ku����j�H5˭���Ė�D�!��p��癮W�V hďr��烩��zY�N]��pD@�Q����3��a4�S�iM+��NQ6����AE�t2�����!� J#�A"8����ķ��{೟���ϡ�g&]�l�K0��A�9,���8�a��h��@%����k^y�{��5���ӷt�n.��?�VA��������>��?R��hO:&��E�)��%�$mn��f"��!z���Q�ʋ7��^���A�������@�d�r�سX����r��'�����ca���?�p�K�H4��/*��f>�:*5�����핏w�VD�ZQ�?�Zi�ɲ�Z㘨�R�CruX���m�.yv�^�(!'� ��Q�M��%ٶ��h!�#��!Uǉd-$lÂ��qW��cꞐg9߰�k!���v�qZY�#�K�
H�:�VA�d�;�VBB��z]�J��RO4�XY^�\�X@imY�!&�qB��\3Q�j��B�I�`�/�4h��O��Ʉ(����������ٗ^�P:�|�E��������������F����^qh(��r�O���r�q%b�r ~-�U_�(�C�1w�Ch�{&��z�����_���ӏg�jE�F���'7�\�d���,�:�4kAZ�I��(@�f������ӛ�y� �x*e�H�:�(q�k�l:oiצ�w��-����%׻��.,L7�q���<;�U�g��y�F#���
yM�w��umx�{t#(j �wR��h<��օC{]�Ͽ�|?�"�~�2��B�H�$�t>�94�s� ��G�s��zݼ��5�E�n��������w�^M�����f��~%s�jk�\�,�����|x}ĹvT+6C\7֜l�ܛ>��:o��/�ݠg��߮�������L"<3 �V�MC�3W��#M����F�V�ю��������gD%�v@�{�k u�9�����^6�T/{��my՜�ꔖ��PL7=����D�8I���B��Y2�M������Ĭ�s/��	�f�j{�7�6���刖�����;��('�ԕ�Ѧx��C
e�Q��4vu��0q�&&O�Yͮ![���{��,g���+t�Ju�u��b���j���^����������#XY+ȍ+�[(�F��$�̲�âʹ:�DDSh�?�
�2p�sGc���OJ�e��fr�$Q~*Ӎ[o����$����"|�A���h�qz��� hçٝ�|�lv�2���s�Į�1��+��B6��P*�F�|0�L_=>���?��_>r��g����.�m��:����½x�{ށ�.>O>�;�?��^�L/�U/cx�K����f�a���@.�G_߀	l4Y��M�SdN'����������V�����H0SY �AZY�}��}�x>����o�ڪ�� ��{1�Zx�O=���,����2��
�^q
�AO/������U��,���۷��;�����v�/�6m�*z%�� :���>�P�}Saf����-�Mp�г��E�n�&j�*U��Y��$��u�Eӂ��v��Q_qZ�b�?̽g��gy&zWN�]�{r�(��HH�%��� X����&{���k�>���$�	�P�@%P������*�:羟��nq�?���K�LwW�����p�d;�5�1䓣H`�}�Ѫ����?��N�T?�U�(i���Ŏ-e����a�$y�ct�˨�W��o����o���7��'|�}�o?|ǣO�}�`494�n*�lf1r�U��Ӥ�4��`AUD�@�e��A*]�6�cm>�M�y\x�.��c#�.
ˋ"ʱz]'$�E��/ދ��|
M�!�F��E���ÈwS�$�ԆギS��^��[��֎�b�T��'۟�:�6�6�3����:�M��]?�TBB h�+��J'X�#���+�@�@E��T;Y�$[�)i�7Zm,���i-��`0T����"�t��^�dW��%�Y5gEJ��I$�[u�.i�m7����m�l�T,�U*`��a�� I��"	St�Pi��S��a���#�!bɭM��ĦMF�Z�f�@|��ظ}3�c\�J�Z�gQ4� &���f�q~��7���U��]���Y��3!P�8���^�f�A���x0�P@��!�\�����r���ѫ����(�
��ʁ��U�!�,pS\�1��LV�A
�!K���ԉR��i_�|��g�≉W��b &�$&����Zf�e�zUyv:z��A�Թ
~��.I��+�ϫ�
�B%�]�� ��������O�WH���`Y�d����ҿ"g��!�"�qO��l%�������%�=��I�k��m����d[$Yk{wY0�^��8A�}��k��x���U6l��IL\e(U��3e���g 跃���S):3H3�W�}.21��]��X"ʮ��>^�7�k8���N,)_I�W�0��Q>c	���X\Y�SH��hT�f�';����P��S�����9	\r�I����4��{Y��O�#^�W��h�9c�.��Ʉ�)����˻��C%�D{�.���!ut�FF�i�N��A
d_�#v[��422$%����<�KD=�6�P�Er�ܧ8\��D.�Z�%A���D��}({	}�:��s��>*����u�I%%���/��v���(�Lg�׾Di\ߓ��r���C�R�!7��V���j�)��҃�[R�4��r���Y\8H��|�.�LT�ok�c%������⋅l����ާ�����⢠R,���h�[u�����-04�~��6n؀5CcXZX|gddT��<��>�~�i|�O>��o�8�t��v&�%�yƉ��W,!xf�^\y�-���0sl�Z	������x��O�m���w��x`��յz�D̺[��'��]�v	�x���yz�x���vH&�VN�*�/21	߷G�Gg�<�_>�KL�N�ވK��Vt��~�iD�4�+c~�<�Yy�p�e\�dp8?,H�!r�)��ϊ��n|B��f�"��,�X����"��Q�hR���@+֑��`yV��9�|� �bJ(�������?��L<��ު�1�K�8��Y��s��3��"X�_���HG'Шf��c�p���a��004�V7���%i�F39Ź�S١�r�	:�Z�v(3K��ť?���}�����o\[���Uu��o�����;�C���Z���a5���� X�Yx3�A��x>mV����q���'�02�ӏۂ��6��u�X?�G�ۖK.7�j��r����(b}Y�v�^�p˃ȏn���0_�`viI�ch&�K�ə�/JlV��0�V�TZ�Ɛf��O�A�<�XJ-�B��G�s��C2��9��h��*`�NSMH�tti��lT0B���!%�d����m��F��"�d��)Qz<@-!�,v�u@ǩ�gɈI0�niU���]���@�C6``s)�K�}|a~Q��H����$�QbXIv,�I���j�*�i.��Z��X���12>�u[7axb-"�A���f�rV�ظ5:1G#X�VQU�A���Pywؓ�U��W��2����WND�@ǃD>'V56A�ȃ2'*Pg�E�V���b2s���0�F�P��ʡA����i�������P�Z��F�l����dV��bm뉶*�7nT��	��CG{A��_)NY#Y�*�8Y�8,� i,�:��$�d�m1X��/��%3���J����}�1y0f��t�LM=~��\=N�+J;�k��W:|L�ga�v���ú�Wt�6��$	�"�h��X�E��}+�ւ&�L[�$,-�'TB�0U�١��۪��1�.���m�$�����=�:�C�6��B`')jJ:��J*ufԂf%Z�Xݿa�eT�mUb��WKx�L�|=y�C�h �[�h���(;`-9F�9�9	������?�n�u��Q-'H�z��֌%Nt&.��P+��a��>�e��DN��xģ�P�:���dI��=V'`~�R�	][%�A�X��"H0���t��6��BǄ-�-�^'s� �S2d�� � $({I9"�H���A5�G�Um=x�HOJ�KD�����]r��Vj�Zn"�j!�*���<�dc��)~i/��22��C�*4HF�~ m3��t)"�%`	�'F|�wV%�V�I(X*K&�{cW<�������s|A����K�D��N���_�C��R���x:���k��g0;9���Y�c)����Le0�f��u������ظe=i�X.-#։btp��mB��t���G6�3]�DϾ�2~��Ø[*"Jiv�٥aW�N�ZB�Nė���8�����������]wޏ��ڵ
6o�g?�)\���cfn߿�Z�p�-HQ!G�TS��n��p����?��T�~��1����3��5Go�WG�l2�s1?��E~dhX�&F�'I*}l��t�p�wa��2��e��P�pt�0f�g��GC��|#�#�naqs���Q�r�I'a�ĸfC&C_��U��%TkE%�V�;�eg@�DW11|�8�L���w���j�� E&Jo-�&"C[7��4�b���E1�_���u(.&�����Ov��� ��!�@��E�!��G�:&�>�F����P/�VhV�Ԑ�T���C��o{ەgo^~U�@x�J�!��7o���{�+���!��4jى�&�hKK��6�X���-�}���Kyͮ`)�Hù^w�)x���-�J� (.�M�|v^�#㛰f�Z�yߋ��ǿ����Գ��B��}�`~��f���I����fU}2djQ���d�����:�Z�:��������]!N<%�)H��!#S��щ�R��F&�QFM�XF��ly����C��P��7�٫����aupK*�/
LǿW���B��*-�gVe����'�1���@�UCU�Mk]�E<8[M��寰0;��aif�n�&F��O�ը`z�(ff��ӬchxP��n�    IDATO�#k�
��Rc���L���mܤ���m) ϒ��t���O�1[(`��H�d���*�VUm�0����,,^P�<���� c�è]nD!P�D�p��e��'�	�*�l�20U0�.�%g�#�ip-o��O��c�W��+��^5ڱ�ڸ,y��W�4[IRԪH�Z�K�G�dD��`ǎ����)���˚g�jz����|�	-�
�;����eqς�:w#S} �z[.rm���p����J�y��6p��g����`s�sLF��<�����p�=�Qu�1�*ϫ�<�n~ߠ$��F�+}-!pO��f�@�Xz�����Q7��T�P<�B�a��X�H[��9f�E�VIw�C�#u荫mI��U��K%,����h(!�F%9NШ�	������)Bx�W�=�C��x)JH1غ-2����Y���` �	ǐ��8�˦�L	e��b�%@����N0�1Q�k��!���"ޠgI�4�G�u��D\�o�ާ��^X�@Ò��uq��(W���� r�w�������&�O�_t��.���D� gw��J!�aW�L�k�8��`������y���~/
�y�3��{X�+�8DIT
U�����/�[��H�����,��{~�'ۍ6�!�1�>� �sM�St�6ވ��B�G�x\VT��}&�ɠ^("� ,@ӿɡ)G��Ɍ�M F�vX���I�A���U��(��/��q��N�(�t�>�Q�����b�Qo�:H�h�/Y�!���ۮ5��pl���ڢ�w�zM	��M�Q�177�r��3y��z��%�V&ׇd6������Hf�]Q�T���|L���2��u�������N��߾s��b��N����7�?����.ž���+��o�]�G��s��-OO�1�_~9���/"�N�����?��GZQ$�݉��Y�X��d͋g�Ը�G:�B:�����e�ٺ�9'6l�#�&��N܆J����^��C�P��U	�46<�n�$�ݻӳ�8��m�&���s:C�\U2*�(Pm�Q�WPGu�yF��A��{�p�$�-.�ס��{� �K�J$�8�H�|�Yu
bt�xMӹ�R�Hv��@����_���?��ۃV#���J��u���������ܻ���A�e<˪�-f��O]v�y���~�{��)��'7<����}���>��?�Кlbhm��버Ig;(�x ��f��,M�}Œʸ�����78a�&\��ႳOF6��D�%b��b`���#7��?}w��Wh��8i�9��d��b�l}�Iժɥy��a���T:�5k�m�.M�ծkä	����6 �33�869�V?E�_2���_���Ϛ�@:��t��N�rQU!�7E�lp�j�``U,�0=5��%Sr���UMƑVO�A���#j�S$T�J�.��� 8��$v����#���� ��c�l�j�Ę��cX\�C�/���~\x޹Ȧ�4�������C�c�v���J����Q�X�N�0�R[��+���� ��T\���RE���zK���Sh�#��e@�s�7>�n���A��{vH�N'U~9���S��4΋��t��Ѫg
�X��J�Ϊi��靗T ������K\v���E�D���)禒����52$��X� ë��-)����A�o~R&מU��R�{q~���1`�r.��:�[.T��J�U�$�P	�ɇ���*�c�Ju:���1������*�P!�L%S��~t���\�=]u�"�� �&V����k���6s�2��x���=�����.U+���a�@��-�@�C�9	k��C�^�q}*!�q!���G�&���}���dӒX��g��cɹb�K���u�QV%��� �Sg��iaN��#r����T��^W$�����>ל_��j��\�xe܋.L0�}n����sHVXmΐ�DIPi�3IJ����� q$�������}�zw2��"�I&���x�K�?�ݶ�����{	��u�+(Q�@�a{�';��j�L?�.�T"�Ԩ��F�d�?�5B-��ٜ�[��,q"j�-b�C.rnP
~���W�yĽ�R�h�k���4�3^D`�V<�֙��a�)�*	/�ϣT�#�j�/ZE{�0N�6�����E����?��ؿ�"?;�J�d�!����XP�k���ɣzFJ�#�7�<�ѤCp��R�cFMь�����h���1>kq����_Y8c���м���ݯ�o���ޠ{o ��~O�wmo��^mO�f֦����S*���!%B�I2ܴ�#�,6lڨ���[Z\����gg���Qr2��[S�Z�8�c�0�t�h,Ma�v�K_��8�S���}���;p���`�Ф
7;O>���'p�_�CS���o�u7ߌ�i�H�(jRB4�����n|��G�`w�q/���������U�H�T?�ev�X�`Aa��K/!A��중��B�Y�Q$G2���my���s�߀����+�<�D6�BeY{τ�1�|ڰv�:��sxz�3R��:�8��y&֭���("�6*�"*墒�B��
?;A7�����h�e�A����kD�1��T�艔ؼa�M��@6�D�3�d��l"�Lz �� F��!���n�w��a<��!,OV��ax`\�ކ-[�;�{b�n��x�hw�B��5�k��v7�����Ld�?���Kް�_/8�D3�x�_��Cp�CO��?���x�
�Ǔ�<�}L�$1<YG	��,S�T�@�1g����t�lС6�t"�f��l<�Mk����5��01�-�cӆuF�f_����x��$��`z���%��EI�Ku,,,�&Hh��e�sX�~�>�����˪Z���41r}����fu �_*,[��JK����k�r� �M	A� 1��*�k��^o`~i�bY�!�̱"6?G3��ԼQ�&�>Ӝ(=�j���2��{ qqA����vpG���KD��s��k����@���tǎQ�D��SN9	�� ]���R>r� ^z�E�3)��X�����0�Ŀ�ZS��)/��\�R��H�Y5�h��M��C8��S12�/�?��}
�H;N:#�kT-�k4�t�\�+�a
������,��@�**?�u����*���r��Ai�o)9� =�!�͆���F�4�>%J
���ǟ��Mp�:#��ì�		��� �ڨ�a2�RvP<i�����K��Uh��]XR��=V$I��6�4's��]��MS��rn(����)�y~_���
��ڔU��ҧ���A��%�����	�m��)����$F�5x����\�`T5�*v�C��a�F%2B�	��+�eWL:�!Q��ρa4֦�tq�?���9�Q�D)�Tp�@�{r镠^���H>3=�|W��e.�#�C%��)	��1!=��߃'||*�1+��䌴I�a<��<%�LQ�9tr�X�@Ġ�k��� ɫ��g� ���p�L��$'�y�Ġ��y����]?���]Ak�q�����ο^L�������;wY���:.4{�9�`���H�v�+����y7�� <U�[����Y
v�	�Q'@�� ��1�q� S�=v���IRn.����*�i��0���5����GN^�P5b��/7m�� �	qal_�{3 �4*M��)�P��?��;q���C�p߬�2)�!�Y���ʥ�� ���9΄�I*�m��=�m��:B��������/�����ǑLF3�]/JrJZY�7� �����G:�L�U���H�H�n����H����%�j[��fEE�NiI^<���$���}��Q����v;���A]��L��E�	r��I��v%+�0��%����Y<�"��i�}����~'���<���яq�]���\Rc������i�����c�q�Oo��tf���0������z���.�����0<2�;������'� N)��a�j��hxǮqWL%@��������j����m�������sN���q)N:}&�b��Q�/cny��E�9G��hM����
3�&g�077#��uc�رy+N9�De��*WQ�_��d�X�����͝x���ϭ@%��(V	s�-���%�ɣ2	JP%�A*�Vw ��!�"�C2я�����O���'17Y�Q�F�~�V�;x'�~*>����8���F��އ��\�lc�d2�1����������ч�i��g�z����޾�?2t�O���o����ȯ���G�鲚�E\ʎ-�����%I"Au�	��ϙ����L	"v�Y)�۬�U�a ��5i��S�hxd��a�y�͎�A�:�nLM/c~���h��9�<x�4�����e>2ڏD������r2�x�Ǵ�1�E��Ĥ�?�ܧ$�M����翉͖d`�Z�N����l�3�-������/?���1�8H����?��8�^ͤ�W|�j�np|_�Kx��X_�b��q�����
��r9mf�cb�HF09yT-��۷b��b��;�#(��739���퓓#[��_f�� �I���`� '~����>��s&6�T��2\x�8rl7��s�/��u�	ظy;��(�(#k$h?p���o5\��h�-�u8�W#��CWs
I�%R�d�I�$V�Z��(I�ZwafG����LU�N�C#j���1WQ�'(��{�U���\�ܦ�է�ɯ[��h+��*=~���åX���d�B����N��\�ۧ�A���#����}�!*:n�������a��X�̯���{&$��$x���מ�'J5������<�}���ח��z���<a�h	�(\aŏj,$3��*�̩��ĞR��\
�F�� aW��J�+������U�eZ`�O��+I^u=�����۵ԙ	��ꍦy�����`��,�x,<���v7���4WԜ|\8����΁�O�=I�3 �?7 ϒz�	qp�� ���o�T���1.*E[K+u)�L{��ɮƤ��cV0����4,��ɞ_�Uۙ���!�����e�d2���F��U�1��r���v"'+�%n^&[ܟm^Ɠ��1һ%ά��9�sV�3����B�FC/;�b��Jؽ�z"����Ɖ2�u{�(2)�|�E�̟bA.���"
�%J�O_^�G�R%�IKZ���I���T�Z�#Y�jꀼF��%�"�6�,�q��_�S���};�ڹT�*��#��� ��L`,���3�+�f�(Tbm�I2��{�7���p��7�W]�F��X�����Dt��	M�����3�����w�EV�e��T\��V)p�|~��5����N�U�q[������Т1UgBp\)�0VI�����zC	�c��1!z�oj��3���״\D���R��A�F	�{6>���c��x�ɽ��w���w�+NB�T��m��/���<�����݄o}�����׃F&:�zTK��?�ןƚ�	�����������O��)ˠK�B�T0��5	��r���ю��,[$�f�V	�0�i��B���]��P�/���}x��X(̫�G(��Р���MU|!����G��bzr�REJM'n;g�x����&�d*ړk����j�����[@8;���L8�:#�'�����^��],���/u��u$b	��Y8N!˂�ԅ�*�6<��r�?K#�Nڶg�:�n?��ϱ��W��&6m�5�߆k��S��H'�2�l
ȍ���_�~�غ}7]sC!�h~���^������y����������w�c�Hv�:�d$9�Ĕ��"m���!0�w4��&�lXD1�sE4d8A�gL�l�XE�/�A�@_�p��@���H��0��(��8vtŒ�|xܔ�V�'	�mg���HM��z�V]r\������f�dΖI*��-���f�΍X���!��̉ō[Akh���O�*Y����4e���(f$VظQ21��� 	c�fR7�h�΢o��4=@�B^� A�a�M�AFh�b���km�Ŗ���ЮK�I�*!��I�p��S�X��5�v[8U,B�n�!�`��R�(0�N��d�7���p湯�e��Nt�	�s߃x���&�^�V+�J�/�a`���W�}sZ�y"�A�W?�a�P�{�j�.J��*Wܬ���7nrzr0�|?�dp�;��+!����|���\��J��p�e���7[�H�1�ܞ4���A_%@L�i��#UQ����5g}c�k�q*P�p��%e� �piEwY�8���0Ms�_�L#�ǫ���������_��ą'�J��3`�ݡ�}dW��.�^�[�QB!�0,vR8��jo��2�VמI�3�Ù		֞Lrl��?vlR��d���!��l�m�r�)y"&�@�:?r9�v���)M�!�������1'4��F�5ּ>�T�lhPl�`��� 1&�GvA�~�W�y��{�|���w�<�Q���0���m�B�8N�x]�+�8����тe8I�v�al�`�'3��upb��R6?3���)�rY�'(J�h����r��{���CI��RQ�[�A[�R��s�X�kTp ��<�k����ҫE�>��������g���O���C�����%͗`f�y��¤�2ˁh�N��c�J���)��+&I��u�T(쌼->+%�u�v�������yv�0�Yj�Vx��	VM��a#���VD�x�o^����Mؼق7�g%�����K~tg2i�A0N�o��Z�<2�%���4d[����#|����j�/J"�D����c�]ж@<;��3ɟ�?��N�bQ�P�@�C�Ԛ�%��T�����A���o������01�r�hgd:a��VS
D��kRҒ�⢠T��x�*as�]&�MK �|D^C���R��j~,d�����]�C�̳����]�o�M+�ر_�����o>W����ǵ�݄��y�sٴ���� �o��-��?�}��������^: ���b�n�Er;ˊ�S�EKY03v-��6tny�.�]
@���O=��}
N9���4�_~��xH*A��1f����ؚe��xS��Rx:z����D$�s�8o8��B���V˅�+˨6*h�<5N5;S��z�>�n��E�|rN�������sR0�ZS�m}}����JGM㹽�Ш�1}xO�~�П�;.��{����������&�'?��p��;���ŕWݨ��Q'o����}2��#��3�:�<����C�����>�k�n�j��W��� C_��������i�T�-��(��8&/i����To&��fB`�Y�X�\�*�l���E��p�&����v�~��O=��s��h���઩��9h�j�A��_97XV�٪��X�M��������h3�U�2 �Y����j��|�B9'Y8��O�z|O��]O���saUCFt`5�/�o�*
0Ƥ�`�V39%�n'v������m�M�ݑ� W¾)����X�P��3����Mt�4b�H�I�>��I�$�% ܭ(�ը6ЮU�70`�`�����dK�b���bs h�	�#僁�a����q�v,�*825�C��b�XA�;߃e�y������3�j������������7�{�/��x%ӡI��
n"V�Le3�J�[�C��fh<���iⲊ�?����&�=���4��4��-���🈰���(�-9a ����U���lϭTd&��P{U�R�1��F��B|xP��k1��*�:	0�Fȁo� �!:�&Y���7�Z�*��߮jdFLA�c���2�ι�� e�����_O�n�>+ry��3@��y��01m�B���k���
 �-�2h��3���o4�����
�j�N�<�u8	�>#�u�u�jl��k~��~����(���!��vx?A�\E#$3|��\ŏU	��`�fXxK��|U�    IDATi��;�����ý6�U��y����K��!�G�Z������{I����I�M�@vh&?W\��u�(���'����CG0��`]���ض˳����9f^PR��7�3��4ߛk�������}�Iځ��}H/q�����b]KB��z��2�tp~���xB+8�s�.W���������g�g��#�dI{]��d���{W�C݌R����|?*,�z�:�����bX��T����G0�Ob�ݷb��Gp����༳�m�����7E/�\��bS#�C�3�ߏ�����TT���Ȃ9}4"$y�	΋/Ə����q�xe���9�M�~e3�_^�����r�U�!ZJ��Q��\*z����R��"�}��E�P�j	�Oڎ�~���߾�v�2�!�Y��p��P^L�!�	�B�O�ga�Xo�<�V�4�N���{��uH] "&&�n�/C�	<��!|�?�Oo���Z'��_���E��"��B/��
�J\P����8���ڵkp��;�LM�����(�����֝�w���ǰ{�c�<6�N'"*�6I��]�궗��:���\ ��X7��l�o8��s2f������Qk��	` ����/}��nۄ���J�KK��<���9)=mZ�g�<��t
6�]��d˅9�t��7�#.���9��{��5`�S��ڞ��T�礮����R�*�Hln��#��p`�AL�G>;��t	�?��/`��6��?��^�>�t�|�~E�?�����N�<���j�{�0���Ѿ�oś.z����*<������o�ş��]���~�����o��o^��yi�����Z4�1]q������ԄP��k������8�Gn�j�;4GAv0O	e���eX�¶��Kr$_'�Uhy6���ҟ a�]u�jO�"d���
-p�W��00�,�����xhK�B�V�d����j����9��[��7����W4�l�\~������werS���>V�m�����c��+bT��É�b���F����*&T��R>���ˊ�g�>d��ޕ�����Ԟ�S���hbt�l�q<6mފd6���yLN�"'�º?|ͯW��3�̃�-g�Y0�c�)P'�(�{tI����M�\�md< 5ށၙP�T:�"a�V�E~+��ys瞈��5�<`�qu��ϻ��IbY�j m�:c9b��$g�����k�[R`��π+�b�	=+,�:gP����fn�
�R$2 ��*�N��IԂ+o�SJ��LS�a2d�&��a F��|�?O^�'�
&�ɠ�l�*��=z�Wi�z�O���:P ���q�`0"}�2�G�;,ύ�<q��Qߞ����`��a|�*լ`�=�o߮g�
�%������p�P	�Ǉ��H�k=�5�x���0G��4�K	]���0�k�jp:&��������W5?H�x�WO-�3.��e�~vp��G1��S�ˀ��Ov&�E�t5�t�#�ϋ��v8a��4B:����ʺ/�iQl�k�>#��`Pίo�.%=!�{>����EAcx+�=j,�q�� x�O}v��}��9V\J@{�S<���'D4��H*_SRG!$Y�N�Ln��&^7��`b��4���g� ��[�1� �8�f\�l?<ѳ�ƀ>�ʩI��*O
q�Ӣ5�@��s���Iӭ�1ڗ�i'n�h�����^�UA~bTE#�G�f���R�A�֙��1i;�3�ћ������̼������Ǆ�	Α�<�̋8xtF>��U�ܒ��u�����
n�8�.y(�	B,Az�kO՚��	=��o�9����#���<��{�$��Zc�x�e�ୗ\����)�Cc��,]O4b�UQ����fj�Ȥ�:����^��f2�^�q�F��Kt)�A�A?����7;��z7��S����v�,���7��_�K\r��9`]��b��l�6��$o96��\,(8��]�54:��{����<��{��2���+!�Pb���L+>ȏDP�2ڕE���X�e-�ص��s
r�iT��;�"
�E$9��.�2ff'�~�Z�8����a�R���ff�035�v���Tg��'w<6ML��9�:�ޛ48��Q��&D��k��q��YVrًٌ���&ʸKA?�@�RǞ^ƞ�/azz�J�Xù��2��!��	��7ކ?��a癧≗��?��?bl�Z|�C��M��{Ʒ��}<��~�clٶ�x�;�Ƌ�]��p�MWa����>��~�S�~�ͯ6�׿���﮽�o��M�8\���@;݇H�n���a0�Z�!!`&�w�}�T 
��V�cIj2�@4�̈́A�O���i�!�`B�(rV i�&�x����QI���FuZu���*��V��66�TVAw�L�����iMX�*����7b|��j�L_\	G�d��^a�d�P��TL�x��˃���w�(��a��y]F.cc7���*��*=X�c�yR6��L"iUp:FJ�;�<��}T!�P�8u�41�
����B�9��I��Z�"�����e��8���������y��{��0�z���kC��/#���P�@N! 4�aB�`����-n�RU�tQ+T0�G��9��?�/g���UVTH�}�~����!yqZ�kg@���d �����DB���A��B��CH��\o{�ǲ�'<x*$��ҝN�X����&G	]�x�m��JeE:2��ł
^<�	�Q�֎���ÒA^��-vt�%^?��C�&[��ڹ>y���u��y|�~{������y��^Q-�_��Y>ļS �\܂GB8���~rέ[�^AmqyY��j#����tH�@��㶙�k���@1�&��P�lvo<`�V�PE��#�d��л���^N��z����x�����@���U�=XQ�r�m)��Q�T���ڊ�q3��$��I��Y��:��ך5Q����@�m�&b��8ӿ����1�Lk��q�y��R7>9?���Q73r�-&z�PSj3�KH���Up�DL���d)��>�|=�ǋZ�ˋ�4I��҉g�߯���qN����4�$��*8�!9�"_�{���?v�ǆw=}W��N���}?K�=��w0����"ŤnTFW�b[&F�מ�H��[��
�/=��?� �g��~��E8��5x���:�|�����q�ӳ8v�(ftJ��i�.ǖIEJŤZ�ҵ���*����r�oøIgT��{6��[�����ƙ{��͛%�̿�y�]z5v�yV2Qer���:
q��i��qg���#y�"-pkO����?�j,�\n�W�n{�nT�:yQ�s^&��*���^g�0Rö�	<��~<��e������I'm���)\z��������j -($��F&�,ͮ�91h���	,;��"��~\s�u���s��,	�N#K	�KIXk�P�:*Ouq�2�)�Y;��'n����!?҇�3�P(/ �d;�F����#r�����w`d|Lh���2�gg��g�M�����l�׭�x���X�f�dM�k�I3!���<-%��5���n����?�j�ff�H���9<��s86I�^���8�<��,N.�5g���]�~��͗`~y��z-n���~����?��lކ_��>��7���ۏx"�|�ø�7���Ǳg�4n�����޻��t|����_����'I�������8Zj�_��t?"� �0�������7���̫cx^����#8c��S��5_��b��z-��5�֒e��-�B
_�*�R�-HIF�lYB�Ā�Zɂ0�>;X��[�ePS{1���ۤ�-�6�E��;�I������A��`�[�"�Jf�&�%<��c���lF
'��zx ��o�2�UZ?�V��������F)I�Q+��fS��L���DĂ{�Vu��2����t-�� �ɓK�*��}t���Nj;��2n�U��5�Q,.�����8��T�؄!���1a;+���{ld����pK
����o�nV|:j��I�xB%�!����K�$వ�� W�z���-�-OΣ5#���l������a�R�����3������a0���2����dPE��$w�W(��B����<���(�h�����സ\T57�?�����p�feM�c�a<����	�C�����t�*�w�L������@�{����Uqޏ'l� qȑ��df)9G��H/��a���n��t$#��j���ǒs^z�����4��y֒rw�V����)Qv�a[Y���^Ʉ��*&Gf�F9P;��m۪�"���Y���Zf�C�&j�3@OƤG�&1�	��������&~�
���l��7!۷nS�{>v옞9�����cG�0�g˪��,y�^̹ R���7Y{��^/�{$-o�՝3��imH9%����'XS3(�2�M����a�Ν�2>��ӽq�VCz �kg��ƔX�&s��hm8�z�%B|>����(��NH4a2��y��>ǅc�E%n����sA
<�+� ��_C����1�+٢�ձؑI�iu0�g����g�k��[+.�
Nپo�[�0;�����Bcv
q�����4�����C
B��0��|,I�!!N<Jߟ�Y�+D���Xs��Dȁ"�N��ύ&ɹK)9��B��8aM�B7@WA�B�I�!j{~��f�l[�n���K(���May9�q�Z�F�Z^qNhT��&�IS��p$[��MI-����^��w��<+��l��ܓU�{��U�Y
�Y�{t�-�
�-K���B�֭݌Z���r�D&�u,��Ν[��8.}�&fg�P*�E�N�鳑�>F�$"%�G�џKh�]*07��X4����ಙ���=��sE�ݻ�S���;�Ʊ�G��!����%�)�b���1V�)�̵���1�r��Z3@�2*�"*�"�F���%���09uXR�#�ؼ}3F֌"���7�����4�utjd�ql[��m݂��<���2��zC��PT�N����Q�sO���ۏg��VS,C�C�Caf�����/ř;�ć>�����H�������>��� .~���|[�l��n���������p��.�G��8��M(7��~��r�ya/����w������7ڦ��^U��o���Ӿ}�m�8Zj���(�Cch������(op׊F����[F��D,x]	C���GV��T5<�4k1w06dy�3���@~�s���W���zτ�P��Th�"gW.��`�
\�X�%�
!�D����W2݉ӯë���LQ���5�|�i��A��c5Ք�k��?1�j��I�WV�o0���F8��*�g��<�Hr,���YоRZ�a>2A�gĄ�*y����ղqrC,1r�됸�-�p��"F�ҁ���L�I��[�2�{��+�.�P�聲�8�=FM>L�N�|2Ą���TmiW�RE�?��A�}b#9B�N]!:i'[��9o��;��pg2�1�+���r��ʄ�EU� ���V~�He��Ԫ���4�d �˩OWRVP�Ҧ����z$���:5|~�|��k��Y`044�f�Dɞ�%d$5�!'�8�aʪ��( �$���d9�#�=�P���dr��+��|1ErW���!�Á4V����Wt9�ه���_���ϖ�Ʉ��4���(�c"J�\	���p�YE�Z"��ő��ίf��Bq��z%F��(�
�~V�W�(����ú��@�h��2XY�2���V�`k�Ǘ�(}r�X0���'$�2����#���f��׼#F9$P��K�cغy�?4����%�#��$�y������M���θ9�XնĨ)i?�CV�Y�z)
q�\�.���-U���J���C�={��Q��I*�֬�nk���#��k`hP��~� �z�|�<��k�Q9Δt��s?�:cLhB�c�� O���"1�&`���HH"c�$�;Ns�/uH$��6:Lt�g`�U���Y����� eF3�<��l�39�b$���^���:��?���t`?y�=�#ƹFY\���:��&�'�tӖ\*YUp�U���֩�t�6dU~�KM�������E9�-�T�C�d|�<��ha�o[�ƹ`��ǎ�)av�7����3������ӺW��{�+d	W��@�}P:,.��E�޳X9X����1�9�BW[W݋t��^��/U!�{��3!t6�e׎2���tSga�<��w���|�S���s15uO=��x�t#	���\-P,��o|-�v�E�"�<��7j�r}C(Uj8c�����]R���Z��+��cS�޿� ��t��0A$�>.���*���<b��iq���F�e�f�y�N��bvq
����3��M �R/��8;��ĺ	�ݸcc���F�'(-�(UP�PD�K��I�1��c��uR%"l�
�ƣp����[й���q�r.LNOi��+�F���їD������?��v?�3v����x�oD���=�~p�5ؽ�	틯����O�)֯Ǎ�_�o�:_��O>��.x��7�<�,�|��~�	L-̡/}�/�x�'?����Io��ʿ�����߹��������E�m#�?H �f�~=�L-n�Q�:4�an�7m�ʔ99,�P��R��2z����+u�R���"#,ː(@n��`�7X�-ᢖ�%M�Ӎ􂙫�Oą�	2�v������C(��h�~�t6L��_�M�C�_L:)�!��x=[��`��N���W�=�v���d`ɱc%�+����a��$Tὅ,7���`=tu��� ��"E�@�6o�S�#A�2��`�=�d���Z�+�%8MH�䨩�G�00U�B˛�A��$�������Omp����޻W�<0ӝ����B�WǜB�`zBƃ��W��mY�ƋgŐ8S�B�u&�b��>Ǆ�V�x<��0���Ȥ��'�7�I"�6�R���&��C��aϪ�А�:r�jys��Zx�J�C�*���&� �``��C/�K��H��wa����#�����ս�ˣ�񼲓d8c��*a�p����[�:ܜԥ�B]���s8ׅ�!�f��׆w8��KX���{L�>�c�b�%Z[t 'V5$e���9jC�^�r��z�>���wW:���S��p0��U���'��9l��9���x%�:ԍ�b�7R�����޺Uά����~x�Z��I݇�uV4����w~p>;>C��S���J�/�l������2]325�������C�|%�a�c�%u�R�'kM+ y�ǯM�s�6F���N�� erأ��|O&�jE�CCBy��ٽ4x�U�C��w��ã�DI�d(�0x旺b���s�[��U��eA��\�׭Q �s\�@&��gıd���I� �>�D�(�	��u�*՞�?odd#�>lߴ�Nzq��w�w�C�:*��rD�nz�x��{�R,#lne��D�S���0��ƹ�<&���a�|�&�M(J���f��.�T���5ó������A^��T
��:;O;UPJ&����GaiiE�4jғbd��g� A��_A�+D�q8���X t�yM�Xx���ÅK,~�X���7	��BR��a��~,�&��S](J�_�h���y�F|�o��w*^~y~p�����S��_��!j��J��V��?������%���?n��O�ҾC(U;��_�q;����_�m[�┓OĶ-:Jx�Q
��o�5�^��/��1�H��MU�X��e�=���C�;wM���y��ݰ�}:��Hf��g9-�E4[5T�%A��0�q=�mX�5��KR:='j�%T���بI�~p o�Q!�X�����B�Ji�l�V��X*�8L�1dq�d?r�aD:)L�Ğ��bar�7��w��y������g��O�w�s?"�<�sv��/|�Ӓ������_܍��?o���Q=��˸e���    IDAT�gw��}���l`��@��������O����`��?^UB�g���S�����Mף�cp,�B�{-d��!���ΘJ��>��Z�$Ӧ��Y4��U_�Q�W$ض� ���η�2��7�Ʉ���	�\|ʕA�^���qm�.�hv��3�J�yJe(BHE�-�7,�*�<�	�D�W<�RO�-ͭ,�`[�]�d+y
_~����}����NXUiS&%��j�OAK�9%�`i���4Ң�M;n~�;��@�)#����CA�_�ê��vYu�S*K����~�<��(���e2ƍ�;6��w��;Yyu� 8AH<D\	�]��?�d�V�O��Ǫ9��rf�;
|nL 8^�m�T�'�3`1<n�{v�\��&V2�f��TV�?VA��4F��E�+J�>6�*�x��)�n�dp���-8�Ӊ�#1��!I.����"�,�)�$�$n�1���BC��Xg�s7p	�K�*l�V鷷:ґ_����ܞ^x�{��L�e�a������E����������P�1�,��w���0A��\�<$MҨ���hx4������a��&�UYÞ�]8�C�]�N�(9�?�Jhpo��}��;�TVY�P#(�9(6܇>�:,�1��f�%��	#ׄ�ޥ����.��;���ͫV����=�1�
\��{L8^�㰺5�����ӡڈ���H�@k�$iI���~O�ezct&\��<�m۶mul۶m�NǶ�tlw�a��}�of�ܙ{~W�U�N�]�jX��?l\]�BTƶe��M'����KGF���#��Z�}
*� f�Ks����o�Ms�?�b��%���iΒw\���@�w�)S�����'V9�-�V2�h{\�B5}�����&a�.���Wd?�u�Z��y�/w��n�{(��X��X�(�g�n%	F?��#�H��������GQ[]�[�js�C��� ,�%By��3šp�Y�Q�|���B����qN�^ɳr�<X�����W������2�7i�����`LR�1u�y,����x����s�#<��������P�N�aXA0�Rf�����E�yjy��ۨ��Oz,��=ǣ��.j�Ұ��墵�r5�H���z�b�;D�޶�c�Gy�Q:��	��$������y�4U���q�z���,��d�.��b��\�����A�t�>ܲ'f���sө�8��iR�a,����:Y^��Gw���^�������M��j���k�mWz���޽�<؉�`�+K?� 0��u˃���w9.�ya�`/=Z����|<���F���.�b9�a��U��o��-ɩ�63Z��ۢ���
8�:1]Z*�ӡ��Yf^CH���7�#W�?���Q��a��a;����|0x���������i��U�Hپ�m9�e)~S��:���)S��pI%e��	ul�V�qs���sן3W�Tr���#��,�]�]������W�����
%���>M���^Qлe�W������)����W�xv��[���/(��ɇ%N\�ւ};��MGBS0A�)�a<�؂z��ʳΌ���E^�"�P�n���t�!TS��DV�|H���Ï�ͺ̓�h����]�yX��?afj/�JM2�$v95Ra��UG���d�F��v�ۆP�F����"����e��t�73���-|VL�gS�[��-��Gk>��N��$���W1Ibv��.������r�Q��>4D5���|Q��j�h:\b� ?ݼj���i�J�� ~0���3aB��n5�j'<O~8Pm;Y��ĥ��yO=�eP�_���80c"��XQs�]7����f�tEE*�����=��E,%����\,3 �9�K�q���#��&�����i�ˣ�)�D�_$㋵�����3e�#�Ƞu�@���S&���#4��.�n3�X���X�v�(�Ii��k\�MZ��'c�*���[TV�6>��ԇ��N���P[AA�
�~�\��WV��|yDf�dZ���Qi�aE..� ������߇i�}̿������X���y���-�6��a���Ggq�.�~U"�Ës[������X�������i|���_�4T��O�r	gPB���i;���"g�Y�ff�¶i����ؤ��w��{q����r��	u��g`��""F����^s��Jz�X�`�i�+Q'!$�x#�I�M��*,�nH���UYn��0��V߮�wY,/��^�L �!�mvKª]lJ�Y�m��E$�,ٯ[�`G�Ds�L��������"�_�J �ûA�nL?�X����P]~������b�G����L����K��AU��f��D�HV(�a�ǹ�]{�a.d�Y�"+�O��;�<3�,u���Z.�rX�ٟ�m$3u� �]K�A�{}���f�Z:tsV'��Ƅh/Ѻ:�T�E�Vꇗ�-s������վ�����*c�^P�|�O?��Z8�3Y	�����݀f\��!g[�l���5����͋���O��b鼱�\(���v���r�W�X��I/w���q�������]�ȣ�Q��f�&���|Bo�{��Myb�R����������`?�2w%Z+��X��&=�l��5}⸝.��ْ�4�Ua�V�*�=/��wQ���q�OG�:���&[Y��:�*�{%�'+ŉ�����p�;�Ĕ-N7Z,'��}h��M±ɮ��.���]����x~��s"D�}ٱ.B!~��D� L���0�jX��}�{�jGK�D���E ܎<���5��=�� ��5�u�ⴚuR�+�?h�A�:w���9
�|Kw��P�W�_ê0d!��#�mӝ�X{�� ������u�m�_,ˁ�If��Pm��=��ӻ��G�����i�z�ƽ�n��Ճ�`�QG��Ͻ3%������Ԍ+�UO�'ߦ�2z��C�u�9�"'$�ՕB�f�$J�"�6-�uƝuѪ�4�k��4�ž׆�b�]���~%I�6ߚ=g�+ʔ9�eA��:�v�J3�i��}k?���*4��hL%ʞ����g&����ѓ��|qҒ#�M;.��ҳb'΃w��RSFҤђYq̤�>�L��f�ҽeɪ�8I�b�-gƝ�Dщm��CyA�e
/�B��f򭝡5j� ɞ�� 7J��R�g�q'�L��~�Ъ}+I���,��]���,zR�y#�!'a�4�3�U�~tO8F���ogc��/�<;�	��f���Z">�b���<��Rd�� MYy�a�8~�9,�1J4*k����d27��F�a���ds�+眚L��C�b� X,����f&T�l��2��9;�_&���[Oy�thPP)䛾��>�뜚�c}	��V6a�賂"S��V���lث�"�af�h1BE�Ɗg�{���9�x$.:��/A����*�����|[��zϒ�^D:N�(r;*��<F,��r<!���Ţ�@(w�e�5U��=L��P��.���}r�yƧ�����8E�<�g{�X0�Y��V�=��6����2G�"ؘchà	�R��ȩ!V����gn}|�{�?a��$���'K���hL��n0�1��K���}�?�ݪ����%�$�bw9�F~���)d(BFA�CzT�o@��;�!�=9��7L���:'�2��`��'�>�fo;<BV�b��� ͜�g|E|2dY��GA��B��P.��ui�����e��t��EuZ���Q{Y��E8���e����D�����1,3P�V	���b��q+��;�eA{�����^�bH�!�y1�;�@����3=C�K�}Ō��Cd%�'xQ��k����d_w=*�i���QMHH���Jb=�x�dB�2����̑��@*�v=RgX<PC�H��S�wk2a�x�@��YO�x�B�"�-�Մ���M�i6}��r�ïU��Y0}0S�BC�?�*Z,0�>�˝�N&�b�.v���]EB{���'�="��{�sh�s��7�,��x�ґ2��A��r�Ә�A����6��8Y���X�x�w���Ϛ�.So���#�vc�	�嶃|�G�g�~	UG{|���5��?^VyoK.����Z�%9�L���{�UY��{#J���|?__�!��)��)	_��^��4�����'C�Z��X�Z���nH.���I5��μ!�:�Ha���T۹���As��j�ӡ��-��P�U�
�qB�C�~�k�禐.��ʃK�j���l���\����~"��!FI��J;�����go��t׽+o?���44��Y���|&��9�]0����?2�����aV�:�y�>p��e5�#ƣ6�Uh6N�?���s�Ѿ��/��p9���Y��k4b������F�o���"��"�%I�RʸH+���p�@W�v�eRlYM���S�<O~������uԜ���$?R��ּ�+���"{����'�/��(O�����2m���G�E�8�����[�ƥz�Ʒb��
�������(r!�*t�
tI���4��/�q�:�R-�1�2�<Jv�٫Z5{�]7k]�0�صg�0/-��m��ZucƗ�ބ��	��tf�yǖ=:�/
�vRc�q��t�� �X�㟹��uڦI��j�2��Vz�l(���X��ڱ�L�W�)/]�)Ǚ�n�=�u�YV�ī]<�V/����,X������r�Č�<z���IO>�n~\�n;�S�i���q��
�D�jԬ�Ք�^�aӉ�쮞�˰;r�F�i�ސ�M:M�ű�Z��8����6��-*�v�I�);�?z�oZ���a㉕0�p��I˩|�?�ѭ7]�]̺F\�휫��4ؒfa�b#6�OB b���BI��BCah��2������
I�QJM���趠	�k&ӗ��wj������i_�ZW�bLb�@���w�<v�������wE�#�0��ln!��i�A��u�$��c�#�ܘ��G.�B�[S��m&������5��hlW�"���r{S$G ҥp'q�W5�Ԏr�����G��b�v�o[�f�k='Ilid���W�	�c.��<���n�7��i g��]h�{�&�7�tQ�:�`�%ލ<F iV����q�T�K�6;�S�n�h�+��h�F<�eT�\�{�M����YR��(o,n$$��m�L��8^���	��]1�Yx���S<[������?����{�}�Zh$�c��G����c�GȎ�UBt�c�2��q[w���t6��zlF��S(L�*B%|�ez�3�#�ӹ!���1�oBֹ��l� q�������j�et�F�I}zl����a8J�d��[va�wau����}H��V�̆<!`�8������y �X��Yq��0m`�'���Fh�'8����/>g]�y���U��cTt��64�M�W �or��\�z#5��O�bN
�q-z'��S��"�A��b��>�c;��`X[������0ץ.]��z�ȥt�(���Ĵ�+�[oc���$�>$���c�pV'6����pk�~���T��	aV#�ü�W��i@5aG���_C,� �t,%
�Fi5����o���(������0����N������#���ta���	����[��c>	XFc{��Fܫ�)2'�{�9,��y}hV'����G�3��N�Ukp�����!p㡽6��钳���\�򾕭/���여�M{����{0�X |��c`�|�<۬"ɝ�_{C�����V�^z����?/K�懨�Rw(_>��!"���o �ˊ;|'�Ͽ�~O��������.��KV��rCNB���>�1A��P�ȴ�g&6mMeâ�!��<L�����b���8H���ǂY��EU.t���K���+�ct��A�/��F��S�]�,�4����z��6g;$��`ɽI����/ue��=�q���C��V����9�Wȿ��8]p( ����z6����=��}�v���0Y-(G����X�/T~�u�����s���T�%?����<
�t����~߿o�����<{Tص�P$|:�yB����Z;),1-���X;t������ qJ&Y1�YuW��ڤt�2,]]B۬��uMG�!��]��e�-��j^C!���Wt�o�3ow�R���ʺ��ͤ?���Q�[�
;��`��]Xթ-s�b>��f�)��Qv�'���ӝ�lt��K��լ�Q?�����Qh���}���i�ֹ�3s�꫟9f&�աks����ͤ(��g�ʼ�TE�y��jh��N28ȆF��?P����eW�"��&_�����:R!��{���G�[��P����ﶍ�,C�6��?�>tN���!9ą�'�Ǽ	G��Y��w_��g��n䟃w䩺�$�#�+H��G��zͭ�
�.^X���n���{�En�Y���n ��/�=���u4\K
��]��Z;6���<��ֆ�ÕP7�t�/��͍�	4��gH�Cf��%�M(��n�f�S<"h�|��f�� y��6�T�U��j���	��s{��p[H���c�?�JD�Cݫ�P{�J�%1���X�a:]m��ÈK�id���=�6�& v�����L0�%������fq�x��&BC��{���_A��ұ@��V�� ��`�bЈY��(��׌$(��ER�F���-"��@�)D��[[٣�̏�Y�e��~E��:�Tx����U�Jr���}/j��������%�,a�Egz�̿!8�����s�lݦ�?k�1wN�y�t��Ï�F�I��G,RQx�}
`\K{
�.@@�� ya���!P>!np��P���m���?ɦW���N���Ģ;�=D?x�l�B�L�-P��Զ+!�����{�@����B
#���<$tx��v��`�z+��خ�n�����!J�#ô�|$�ZA�aГ��S�c���O���y���q3����ʠ���샰)��B��t�E����A�~��#l��_����;>��:�v��n���h�-�� c�xi�Q������Y�{l��S���b���v��=��/'G���s"����]���i�Tuz�, �fQPX/x�6���RK�٘���(	��-}�r��1��^�9T��F�o���>���}���B������uB
i7�}� ;������`�H-�L&1!��]���dJ��0d�3���(��dc���O?	�؄hP��1��Xw9��Nr�Q�8��b%iae��-4�O�꽁z�4���y�͢��g)���w/K�p�K&���ŉ=t���yE���]����k}\�d��F>9��\���������}��-Q`O�9l�&��_����?�uk� �0��?��l��L�>��F��tI���S+�+�EY����s��P�X�6W7�\*������;�.|9�t�3+�sNX�����nS
ٻ�뜳V�U�5�=<���(:sq���ԩ��ڀ�|�� ȕ?:[tU�to�Dd�s�L�M�Y4�vo�I��>J�J-%)��A�b]��o�ks�ᦘ���K���{����[����AfkiP��.j�AP�=��a���v!�oMtU2a����K�'H��97����p�f�׃�_��O0���s~X>` �����%��
����8i���\����C��.c�<^8C5����0z�>5%%š�3�JY��Y���p�mE3z�:��C����Ii	�c�ʦ��Iמr�R�����7�;���oA@}����8 ̈-��g��6֒q%%�)��A�\bf��塠�iǆg��×�B�k8��u�[�q�ž��樓����,
~�&�ʮx�07+h��rSQ�)��@���zD������P}�I�>G��2����V&�)������t��|���ث#�T�t�
T��܇+����d˪�LH%pz���{��h��4��Р��k�r;* ̾\`*�T����.�6\>:ȉ	0���=�f9Ԉ5���^��K1L� ��
.ڤ��� 2f��/�堜��b�a�弖Dj�q}�4ّ��;T ���68CP�+H@��8'�e�K��E姠������'��K�7��l/�Qȃ�p��G_�����UϪ�D���R�9�j���u����ԙJ7��� 6z��T TH^��~G�	޺;�N��vv�j6���X���[���@�bcT| kgi�� �iy(<e���4�2�;�(]�a+Z�>�4l�����vd���j+�����;>��n�T2>�z�̪��wY��Ϸ�*�/r�]fPX"�q�( d��Y��J���k+so���w���6OOX	�z]�'ྲྀ�0#��<�J8�<$,:xU4�r���( ����e�F�ܬ�䈇z�l?Mx�|�Tܑ��6��^�Y�yL���-�cA��8T�	�}��K'�u#�w��ܱ;��a�u���ߺC��i�zYc���+�}�G�F.A_��l�G��@�/� �H|�L2ar�3�ƭ�o���b�,���ʬ]LQ�-f�߯�'x�����|�'���;��i��<IU*��Uק����g��FJm�#\DT}���%Y�'e�����3�/F�i�c<;��7����ݎ?�_�~��o6�P��o_'� �9��=*-�ħ#�~��y�2Z�'��.��Q>Sr�,��m�1�zܺIu�,�Y?�jR�)��o_�����/��."}���P��-��k�a?p�=��rol�
��Y�iN�f�v/*�D���.�әY��7O�Q��s�K�Zsi��n�y�SS�ҩ4u�Y��f���=o����uk��a�Y��(K�l�"h0Ð�"�x��h��&S'��Xle]ӭ&X0V�M�O:`���\W�D�轖��.�pA�h�xN̨m�~�J�� U�g]��6��|ŋ�+S�|G�"A�����S]��N���\]�}-��K��ɫ��>�N����Oj*�����`���m�1Qm����8���h�	�,��I��AZ��B	�K]�Y(1����`�BdkSڞ{W�|� �A�.�YLq��yF�g� ���� �PI��fl��R�n8�+�?o�&�����e!��1lC���w���*��i�pD0eԮҍ�����:�:�A���U�ӗ	L?�\.�'�3$�o&�#
cSj�Ĉ��@.Kt"��P�n�4�͊=�W2�?�ZѩÑ>!��}P)SB���T0���X8SL`�%3*�Z!�)��r�57-����p?%@Y\5C�m<n@�1g��a�a�u�-	������8��`#����F�)��x�bCi���Z2�����w��*�l7_rΤ��0;[�KRO+p��y���c�9�6�$�����ЁL �Z'�	�S�;����q,� گ/��a(l[b@me��Ψ�Z2Vf+E5'´D Y�1Z�E�-7AqC�y�|��b[�a�1h��r���H^$�|H���
־��Ê� 12}�22d�����N����{�F_~<�D����֠�6OO��\��1��c_Qi&�5v�X���O������R��'7���|��8a���yJh���,H�Þy�	��O���%�3�j�a6��SwGg)�<�$��8-���j���a��:���Z�QL��%Z�K =��ɀ�'<�#\��0h�!���j9����?TMbq;����6^�lQ�/!^�9�DB������e��ҁ_>A�=��-I��?�W��N�nG;����ދև����"�y�[����G����w�����Y�oS>Wes�7f<�GV<��c&�.�D�Q�������C>M.i�5�|�f<��N�"��s G�w&W�̘�Ǌ�DN:mZ˩��$�ŭ��e��Y�����14�7�!�g�������d��t+�U����q'jZ'�������t+	1��G�'U�#V�u��Q�z��)8QReի���ž�TC�c�u,���e��J���^�(�,j���\(�U�*Kx��h���8o��f�-��e�ַ��b�Q�H�,�J9�F��|(���:Z~��Jv˭Ӄ�t�2ɪ�l�Y���ۢ$@�̈�eu����Y���0n%/�{���֮A�����j�?u([����:¡1��iX�[�9"»m�d[|�f""�'kW�>-���M�	E��x�Sԝ����6�)���/��=|�5�t�F(��1�}�A���G��8P�������b4�P��x�� @16eX��^�Ÿ��aA�52��njfԣ����f��Kp��1��
��ǀ5��e�B�|�׌p �K G�XL`�l�.�8��Mc�}G׮7��~�\�Aj������M��BGM����e�$K8�~���r';=C���b��u=╇Y�	g�ŊD1�����Mq_�y8|ȩT Ao��]�����9�D �f�T��*47��J���(:��+`��B�-��oD ���(���$H�/��U0���X&i�g�[r��1���!F�2B�d��6v�հs�?!y�7E�aQo׸<Z�c5p�{�{ֺ֟��|����}3����+����B)�~x/���j=��#�l�2A�m�G��ξ$���-��#�]�UH�V%A�qz�O ��(�M(���a:���J�#��W�x���Ё����n����G��Ү�h xC��u���O7s�?Sߊϸ��	�������W@ҡ�����J�lӦ������P�+��a�~�v����������hs�;^�Rq���/PA�?>��e���ɮ}����c<I��������_�/P��x=����lEd��r;��.� �GTy�j㪯ɥ;.&@SQ+��1�b�t	B0�Y����f/k0���P���ݾ5�����^�ư��;�ֽo��wf�8�diÞ�& ���ҾҼQ�P���I����ǰ1����tN�}Ϟ\��V�k�L�8�8��ުEl�R�c��f9CoF��GX�>�.ĝF9kg[�[Y�(�Mvt�v��#�@�8�j�c�pQ�������:�*mip�s�o�M��¼F\����t�6�P�,XCM��N m��6С�y�t%rh���<�6+�^a5�R6��~pF��"6z�y>;��=ـ���:�ǽU�ɮ'�Q�(J�Y�v�8$͗) w=�m{�Kp���v�O��B!4��_�/��"[;Ǐ�	�z��|�9�a"��o���:���q����\r;
����$�pS=�T�dˑ�ʸׯ7����Tb0)��`	�'I����β���'J���c�N�@��9�{!@�X5�v�[�e�1��|$�%�Bc�1 iO�R`�%�.�!T4������R5r���v݄�fi�@�w%�1�t�Γ�Y��P��Ek��$b�߶��S#��sX�+�'�l�<��~�;T�����-ũ��*	�]8C�����:�#�\�W4��e���L��̱���PM��"���}y(\�0�g�<�)x�;/"<�ꖮ�_c����ς8�L����?C��8b��Tz�G��%���~�{IG �ņ�[p�-�3,T(����eY(,#��7g�r�ݲ�p����V��H�����b˄O�����=�i��t�V��0����|B�mv���w?PUcYf�^B�}�W)��{���[w_&=�<���5?Ze�����3Os��;̡�ӽ�kOH���{
����X&}�%s��g��vc�NtӄX�謭]o�o�t�ܑe�����IF���ۦ�s�D���oI\���AV�%�	��O*�WO�1��s�i`�|9�;�V�{=�Z��(h)ע�Nc��Lt.�Y���6C�o"c�5K�Pj�L.:�<�I3�k� ��Ѥt0�R��lF
�n<9��ƣ^!t�W`8w�2̦T�|�/׊�9
�Mʁ>"<�R.W
��[;�,�4� �@x���V����[&(H�7��DOJ��{�3 0X'�O��e��!�M!�Y�,��S���Yp�E ��\��&�M� �	2 ��AR�T�U@�2j�Պ��^ȢZ��(J�����O�vk�2�{#�-�ta� F�a�/Q�p���.Ƥ�ñ���Rh��/͈)�Y�j~k/>�J���K�RE�&(�\�dy2�f!�ؑ7�T�ڀr�0�˶	�V�����#���s�?I=���C4% ���u�B�J��}b���!!�2 �9:��3v��� �dix,w��޼�7'��o	�t��*�r~_db��
�N�(��wǌ�#6=�=�N�A�}�0�1!��]�GR2�P��覭�#��{/�O9�$��Q^���\G����� ��g�܁�	,O���ܭ��U����q�b�-=�7��y`	�"$��&kBi�����R"(F�u��O���?|&�q�Ʌ���t���=���s�R�O��Y.I���wT?�u{�U�����gg�®�?7�o0�ټ|� �+�u��9���n�]�l8�%[[�����l�S9z�5I����[1rЌ�.�������n+^��kGvk��:� ���`�^��m�$٢��fK���&��dev�)m�L���9�4�j��ra�pL�t� 쥺˙rH�C�<Ny~m���7)e,*���M�,bm��J�X���.+��[e�nW2����g}�v�ܠ#1w�jYM��b�f	7$Z��l 7�\��S�'-S�D4z�r�(~-�V�2{�Ie-:/odu��ٓ�β�*��,^���i/��	.E��K<Rk��t���Cw},�S����P
����b9����^�#�^}��&[,����G�H
�
 3�Ϗ�&���Vt�i����=�ӕ��Yq���;]�\.B���҂L�#	f�4Q�/>��,�Z�р ȫ���-='q��^9!�P"@l���NI��)�=j�4��2�.& �]8k�bfk�/1�ѳz�gˉ�N ���B�Jk7ˍ���ac��i�J%דd��h)���bt��H����V�jA*He��.�1Ĭ��}C��-l ��\�����H$!W`ݯ5�xa�;�@I!�Z���A�Ym��]�7����5�E�y4D^�豕����l�ooX=����Iť�C{���6|6��'���篋��2����Y��[s���FA��b����s8'����w��)�����=UBG`?e��Řq�?� ���rl[d�mG^ Kh�2�4_m�N�{��I�����^���ꫫȺ4�-��SGJ>2Um8+��t���Wq���=�B�=��+®L�cU���br�.��yL�е�6� /!��:S	6,�[@7�y'��,��V㫪h�`f����<���-""b2H�����z�z̫��I��$s�0���W7�H#JW�����W���l�")�R�W����C�m���M���9y��)+��rᤃ�
���rE�3F^M�
�U�h�r���@laa�9B��Mnؖ��a���2��a�(�4�m����K3��{� d�e�#�X2�j!컇���)�~U���@�ɟ�<�@��䐵$т��Qj� sd��H�ͣ��Q'��s�d^���� �i�U��9��4�(��?!� �Pe&b]�X<?�ㄑ��@~ɜ�
��uX8�����t&b���(�D���'$�!�]|J����|�,�A�YJ�kǈe;��-�(|"t�M`�`S�*��&d�ٖ�&�}�9�^�l�TG��\�@mM�a�I�:��2ؿ��7����5�a@B�qO��X�J��1��qFވ���X�|�УE�?|--O�pEc�+N���ߓv�Eqm2
^h��v�+
�J�-��r��z�>�$�~Jϱ��-I�j�������Z�|���'��x���(�2�Wq��l��Ϝo��E�U��IP����N����z��e&�:���s Rue����l���H�;�r-�5����N:�==֠���%9󥮠!���0�7xJ��q�e􅶨��ڠ�����!�ꦟ�n�Y7/J�PQ�nm��=/JS��\��w�+��F�,�g9��T��ӭ�E�	�9t�(�>�9�-��L�&G�^�8<����������}�����TKm�4�m2��ܖ��f�uī��Zl�ԣ�̔�T~�k���XEc�cz�Z�aU�����&�s�}#0
/fi�5���]�[_U����Ɛd���۷N�$l�g@^]㨐�Ț3c��u����!��U9�N�s� qDz�8%��E�WB�y?ȉN���'�=�ɤ,Gi��)n���GL�����i��-�.U�eN�2|��	_����F�u��Eօ�e�!xBj"ZS+\*&��׆[�Nm�NbzT��mh���"��n�o���MG�6A����4duU���!c�������a�g�rS��8�E�g���dy�=�C �IS�Ek�% 0l\^A(�U���7�Ma��<~��dn,<O$@�4& ��\�2���=�>M�%��\^9��7�����"��g�>���'���[x�oӬ�ܟ�[��ϟ�s�e�K'��C���	:�9��v������49��Ei6+��`���/�j��6�#�����|Y�S��nssO�4�/k�m��V�/�պ둮�k��+�r�5<�Ҳ�J_%�)3�l�+��L=����(C3_@�.��d6�Y{��6�hJ-9ԍ>�"������\aq�UWZWݵ���ϥ���Ί�KA��d
3f�1�p���#sFF����f#[�N��f-������y�pR눠MO�;��Z	V�h�M�6�N��ծ[��q�m3;��|�"٢���&e�;g�;��J'Gnp���RH:e�h�����d3��li��j�	�A��1������R}�<v�Ȝ�%^�����a��	nM���$-�,S`��~19Nx���6{ь��:�1'���u��>����#9��l��� �����:ZHb��P��@қD��s����J,��� ��������������:��:�ȟ��	C!�k�%��`�,~��E��ʙAr5��u��cw�^:��8|2�c-P^�\u]�>}p,��`�{<���E��	��tc��s����4���=Et�z��<���_��߼�)n���r�glb28~v���ٵ%��Ő@b��XjC�\�������l���քO.ǜ�*�l��[��\�v�[�>I�� ����/����~h��r���u����I�Wb)Zg�}.uzH^�:�	ǜz�E���e!̟�4����KiK� k��x�E�c�����o}N�/�/u��S8��`���U �2Y����V��_^'6[�E�nj�33�|�++jqT�;y��:d�" 2aX�q#Pc_n��U�5k�<�̔A�"�Ӈ�ϠI\g&��}G"�5�ޟɉ�.K�����>W�x��aV�?�!@�&�'�-ѧ�q!��f�=��W%<6g�X �Ѡq�!�~��T����M�Ɉ�ZLJ�+C��N��5�M��a��{V[����8{��?�� 	K�=�o�^k�^Cҍ �R:�����?�_?5z[�[	�>z�)
OH�9}D�|�w������`
ݿ0��m�]�*�<��"���p��mj�bwο��ZQ���\|����%k���#�M�)K�q�z�춠x7�.K%��"�'�l�ƺ���[��j5DH�	l �V
-�(��3���Ç�����2�YԦ�ӏDo#?F���yd�������!	���ޖ�C�[MO��imY���.p{�<�/=DצV~������rޚw�{
$��%ޚL�H�&�5���a70��TcƉk��;zZmkmkןpf��r�̫m\t�S��q�j
/B����7�ѷ�^c���bL�����%?������rY��e���N�{|A�N�{�n�l%5o?�uk>ks��y��tY�_|a�?ވZ�>�u�R��Ͼ�G;ט��[���a�q��=Y���#�0�]����h���/]qH�D�)v�Vk�g3t������w��c6TѲ0~��P ����`K���ʽL�t_�T���g�#�O�kΚ�(i@�k�sԒ�r��S�~�G�&ayz{�$~}Tc��HU]mn��N��i�܉Z�^,.��M)Yu�bmC2�?��Hh�f��9�Va��NrM�D�lw>�6F��-ʽ{WM�ʀ����1��Ņ�ԞZ(�ڱms\�R������ϞWk�2W-�����,C���l��ܮ�#j���R�r�c�c�	Z���w���l3h����BH�݉q��7��*��H}���ˢ,>=�&��llDM�f��mSm�%6�,���� �!m";=,�N��䲻H���ԕK��=������k��TB���zk�=����{HA��w��P���Ï�͞�w$"V+�c,��\��!������c�q���{o�D�ԓ�_����?����#��ҁ�"�����/�V���n{s���A��:&���ct���������_�Qִ�� �y��
bu"���PK   yaX��:4�  m�  /   images/6ec16c1e-7036-4ea0-ad85-1b4c89c7aac2.png��s��Ol�v�ض��vÆ'��ƶ�6�m�A�4<�	���/ܗwg��W����P�GC&F  h�
2Z  T�u."��_<ῄ�`�	 ���ϡ2Y�I �x
EI��}��t����W�1��V�9����SMLD[zx�hi���� (������~�}��g��6�($)�3�TH��Z�k�xO�! ���9N���� ��O}>�a��?��{�{�#�>'8��d�W5��8��,j��N�@@�������J���Inf|�y�<�X/IJ�D�XXǼK�Թ�1�<��Qۄ���$����F ��[ib͡��1�#�
�/�H=E�����f��/q�y�/Mٝ��u��NT����rΎ˝ ]��'��%�'t���
���f�Ŭur��d�7���{�
tLS)K�ih�H6�@�Խ�ϝF��'g�u�A�fX�쒕��q�tzk���6��~S�'G]=~'����I���|��1��5������]Y8����^-�%�*d���L�'0��6Y��{��t��xEvO\���a5kO}OT��>�݁sL��G3|{!����Vp�)�7]l?��U�1?`4�M���M�c;�:d]S~ fjXYjV��7ٗ�K�^�]C«�K�S�!�Cfw���l��-o��q��;PLJK�A���(ݦ$/��=����6��|��`&,����_S�,�}�N,YŦ�kO�oӠN�#E�����2�Ns`���d�W{ß��� ��P��/g����
��"�N�gb�:A�Q����0 j?8=��T�(��K����7�ޑ�ԍ��g��N���=Q�`�J�,�ͥ�l���o&�xg ��W����ջ�K4���9v�Ԑ��'y������׸	Yv�������7�Ѿ�g�ݯ�+�,H}��Y�^�����1 �[�N����J.��݋|��,9��<5z�#���s�2dfC�b\T4���[Ͱ'2�9�O�Ae���N�� i�8mġ�M1���)!�����*rVz:�	�N{��flN:~��v��E)Na�4{p�����`���է�"�����;P�[!��4L��H��R��W0��	�6<�6<���mUp4%с�<���S,�Y�������.��VN�]�p��U��Gv��X�ɩ�;
�K�t'[
�h?�8r����&�P�'�����
T?�����a��B���^`,6a8���qjgⲉ�����r~�Tn&�ujg���"��+	���Ҽf�(:�.;�����yJ
Dw�탯%L�A3�{���:�*w�;��ș�9���*�Ȼ���2_3�	�@�͆�9T ��	v�G�"������v��PU�����n��SI�*Q�^�@�~� �BH
7���X��Y��2+ _M��e��NY_ AE�jqj�NG'����<�q^ֵ��D�SfU"J/�?�1�:ȥ���v�e`8dO���9��#��[�7��3wd�Di��JGs8���T�6�<}��|l��|Q���Yr����~��yETd'�S�1?���J>	PRWWoR���p�g�W��
��q>����F��ߣR~ȫ�'��eԥ����5�d!tM���
�N�&��QbOdH�����x�h��D���^T�$'Yx����A{$��saC�qk�#�	�{�y�珞��O��� �k#6s(T��$϶����J�� �|9���������9��Hh�!�c?#}i�I���zN�,�M�����J�[2D/ٯ�[�y�`�]
�&�2U��e��^���]��������\��
{Q�z-W��H,	��ּ/�U��_�U\$��q�l�j��"5���B���2�8�=L�߫�Ȱ��k]��&��}ںXS���1]�p�"x���ID\;;���J��Ԏ�f�ٸ�	>��8?�̈́},�h�{��A�+�są`**N�ɝ�3�I�V(��6�[�����y�T�y�k@4u����2u;z���k�H,5�*Ǳ�ɇ5�j�g�w1�(�Z
s;���Y�����K�z���g�����g�R�  �Qǹ���Z\�9��5u±�x�lѝ]�	��[�(2�8�!��4�Ȕ�@��y:��������6[��ޙz�9��x��� �3��	'xѲ"
�m�(Fg:bC�v��-Tr�)��R9;�7���mlˎ��.�
d��ie�4	~�`�#�Q1� IrX�h;)����6�Y(n&�.$F�+�M�~��$�G����셉���0���y2��x|<��Ǖ+ݷ�>��Rm�=S;
��'v�"u�b�G_���AQ <�;�/" �5;t� {��S_��)��ѳ��s��?��6�Ě�*������i8����X����hQ[r�d��ncm��/��XC�C�/�S�k�7�%�b�V�*���ji��$ 0��C9��g�Ut(��2"ٝԐD�d�O���-��F8�O,Ō5jOcϦĹ�7#��F���FB	P��m�v����˯���t�/h�-���w{[�]�_��A)ή���qp�S�EF�:w�X�!M�Ї�I&�h�' X��a9}����a4�-/}ΎF
wH�} �ڑ/sι�fL�9tW_���k��s	��akecxI�o����s�ſ=�oF�MŚK�+�fξn��W�H�������llU6��ϊ��[���H�O�3�X�U�xL)�43m2��-ۮH�M��+L��y��Y����?o��\�v{!Uc���c�KkK�U.I�eeD��W���;����/s�Q�*$&�sH������l�\���mYa�&�	�]�ѵk�n�a=���rk�ϋ��s���i�1��ߜfPmQ�H�l���l���2k}��ޘ��I�4�\ܿ^�������8�/
�hl�{��f}eS���0}�ptn����'�=Qbs(�#��]J]��`]^]M���<���}mD�f��8G��Ж���?U������V�#�"���ފ�)����C��97�?]�h�M����y�n"�*a�yИ�+|!�|X͹T��l�\��÷Q�}h�j��Ng�kn쉣ț�'_�H<������s�҇�ޔ���H��
@�䅈�z�)�ݛ���_e���r29�"�g�Z�Ϲ�o�ʔ��JZ=kԇldst$����	���J��Φ�X�צUw����#/`�XW�Px[Bw���B\���!���:a�c\�W���cG��	��|m�[m6%����|�C5��F���T-�r?]�Q�gFZ��NVv*��b6y��NǺ��\s��N�FlL6�խ̦Ѩ�`�[t��'���Ͷ%��Q�BT�"��������aІ� �`���sR��E�����\׶<�x�{u У�Y�u���$~��ms�S�Y��5����a��e�dl�ݞ�{X��̯.�3{^������^�n=�04�2�Vn�Z�;�)~T6 ��<(G7�D�)�d>1�� g��u+�Y�����K�gw���YT\o鱇b���ra�")ra/ :,�t˘�������+nz��eMa
p�8�����țӑXޔt�?�Jwu��8H4,����c@�ol:M�5����@�Yx&}��)�h�w�i�>[)c{��LFe��c!L�p������o��<����\�ǋYץp��}:�*Na�EP%�-�wi�4��I�ry?�������2����2��[�Q��E����b}W��54h�t�F_G�]@-T]̴��ޖ�N�XA�Nc�mv����C��m'vD�Q��2-�ڗy6�1���2I���91���Հ���,-��2Y���=!��R�Q�a=�0P�0�֜Ci�[A�2�����~��fFva�󨧠��:�NB���<�P<WF����(cuc��T,�/h�K�E��d�A�¢�rvvU�1��OϦ��F\#��c��_�� #�)s�6=���� L���z�f�ӠP�l�N���8��lo�nߦXԃ���I/)��o�l\_܎��>��}��tB��P�f���q(iY�:����쑍��scM�s!#���xv����qd2f�'�Ʉm���#�h��9Oc__�I(��3��*�4&��h�q)d�񬦎�JN��eK�J�V"kSmOp��]M�*�9��t�@���7FJ���<��Y���|#�	�Ʊg�.;������.�3�ڑBJcOݯr�:K�a�0#����( Po�?{)Tq	�~��!s�f�v�=� �kŠf�k��*�\ITh=�Y}���.qe=ϼ�/� �<vB����tl%�v�{q�ԽQvv"�C9��0��r�ɼ�v�}�>���Ո�ш�w���z�fd�Ûa��yc迊l�-�y��=	Ga7�v�$th���C���
�4�w��m�/5Q�ҥ)���f�5��"���{Ȕ��֋�'�0ce<������(,�o�sj��w+���t��v0�ٚ�;sAJ�A����Y�Y&���B��r�0�g4�2�OQF*�{[�GN�oEDN�����_8��Ӟ��l�`�o��̙g~ر�e�I��IV10x]�F��;��{L��<xU6����kV�#�����,�bα��؏k5����ж���-���zg;G�4m%+A�JrA���ƚ}�u�7���[gc������J2�����ܵY�k�gdџ=����{.(h�k�l�B��yLY�Cd�o		1��Q!D���j��<,�6��u��5�� 6�a��u��.;�D����5H�����',��_�e�p\-���l�<I-&�3n�Q��ju���3���Migi���׬�\2���   �x�ۛ1O�ʊ6���8v��I�@��`{悃�<��$�*&�|��Xcߺ��hßt-|�a5�*�~�F����3Cya���j'�ޕ>�(�4�G�	4�YL�� ��|�Հfl�_���gq=r=�4D`���_�'�$�)9|�����w2�������Ac3+����h�Ւ�C,H�𷗕�3H.|����4Rp��7�C���B \�'�#�k
�u��,�a���TS;�����Ю���VZ-N�&葎g�jgJ�66�$��g�Oɮ�

vO�~��33�KpO[��W�Dʨ�$�8��aY��08���	���a ���k)�q>��O��$���k����>�uq�'�9�hbM�~ex�Yux�B�F��Q:�<'���W^�x*�ҳ�g 	��>�O����NS��3�^e�X��x�pR]b ��Y�}�o��p�������E�=O��:"�.ԕ��_WJ�68ߗV���J�bUî�ߋ�S�E��G3�{���O*OG}G�pF�����[�����{�oR���v�%�9[�ɰz���A�(4,Ȏ[���(|���5��p�QAWoğmw�8j�@�97�4�U��mf��΁<�PCF��l��)R��~�+�!���>U�$�%�j��gxv��GZə��g���?$���L�y�iR%�ɿ�������x�٠|we��u� v������s����50B�hX��]F�R(n��<�K!�o���&=���!J��pv�X1@�݌�T�V�{��]@��x�OԾpʹ-\�㺛�a�j�i�b<h!{��ޖ�T1�S���d�m��3qK�@!�i-	�>+�������
n����/p���$,�?���'
�֐�\D���ߣ�C�`�6����2�9>i�������zQmI>
[R��Fp.=��>i���^E������)�p63r�0�x��=�ǡW;�j@7���g�S��p��Z<�#TNB+oI���j븡@w�6.�ŁAt�x�t�ܿ=�����O"l$ނ�u��{�������0�� �G����{E�Q�]��][a�s9�jL��1@�����^C�Y"-�3��<�_�!�pP)5(�X7��� �͞2̩jy��<x�mZ�0.G��!��/B25��<�9�B��Ħ�Ш����X��N嚢��.�ӊ��3:�|sE,���}��E
A(+X�g^�!�oxL�		ttK|���wi�b,3�\ �i��ֿky01�߸�\���pO�?(��qf=85������Ѫ�vj޽�P�#���<G�cP�!����Պ7(@�ڙ�l���CF�\lb�O��v!���<�Id�9���%Ԩ��"C\q$n�C��2��*.Eس�}���|����yO�ϴ[�ImuBĬ'B�C�/���z.0/\��SĔ��ǲ��iiW��2����6�ƝIHk\�54�� �����EB٤IKHP��F�U�t�x��}?���I��
+�|�|:��!>��gόJ;;*�:�>�-^�!���J�5�×�j�~a���]����3c«3U㒳�Ϟ�̃^��֚��pB�^ԁaz�s#J��t��[���N��G$[�H�[f�b��)7e��7� (Bi:p��`pCLߝZ�"w��{r=�	�/��>=�_�L�� P�8+E�K��y�fv�'�72��S{��r9=~�	����D�O�'x��
r?������ez� -���V��Z-j�qK��hJ�a�+��Nav�J�35��hn��9�=ћ�4oZRF�z�gp��R����ɳ�V� �KU�91<�xF{!8)����k;���L�#�)S��&�c@	�)����4,@�Ъƻ̊���ا�	ʎb<C�������a<C�e��Rc1KT\ ���W�}�s3k�l<����;����t�l�4�S�c�`��=��r'��2��4�w���a}�QU9z��e�n�%��1��?���x%Z{He��H���ĸ�G7����&Fk{5�E��-)�m�Qd�NO��(p�"�s��K���m��OL�0C�1�*Ed�|,��a��,B�m�QfD�� 1�x:~�kqO��I��x����� (G�j\V)\
�@��H�E�4y���j+hŇ��G?�A'�sL0���ԭLgB<��߉�|)�N����,����Öܪ���\U�_���0qƈ/�6vs5�k������Q���4��7���:.J���x��[9��7��{/�޿#��Q� ֹ�'QJ��5�<G���lLw�Zυ�|�߅ew�����%WT����Ӣpy�f Qʙ}6��Z�Ԕ��(��q�\|�D��5�"�t�!�.�S88�l�]T/��w������{9�ɮ	�Ĕ�gͶ�r�c_-?,�AYa���dA�)J�ު�"!��U_׊P��#�D�v�ƭ�jY���k�O:��ɱZ�Zg�<EO��i=3jd�������+r�Ka#=]�AhV�_�=���!j.ĞbG���c���ꢨ�%}k;0SR�oL��4$�9�

����_{����؎ �%y�D��M��%��.x[��葦�=�1�p)���+QU:r����2�v�V���{���?����ބ��N�o@��� �J�� ��1������1�^��k|�y��5h�?��od�8�Иgz:�&��>��.��'����S��s^�E��7ܔ^O��Y`~�u]J����zo�����<Sd�^���m��z�h�H�l-�͓H{��'���6�}��nU~�ߘ�\o�3^���b�>�uc��h��k��
�C!@�T��gn���ωܱ!��
�ϰ�3��^#qƫe��L,Lo��Ȋ*=�
D�^^V�?���b��>�=��Ԋ��tB0'wV������$[x��ڷ��6�֔��B�L�n�Ǹi��s�×֣������������[�)��ͶA�b�ڙ��P��s+k���.EL�Ff�(2U�q��N�0�M��$��̨B%;>!# ���	�@�hd7����k#>m(��=q]
R��aJ��◇M��Ժ5IQ����- ��p� Mm�F"�*f�8�3]Dl�'��7�S���\�	iID)�v4��ކw���BuvZ�<v)~�����){����Ǿ��a��xH@�c�Ǟ�ܗ*YKL�� y0q�q^x#]>3v^�ʪu�N��Y��-�R>:����y����5�:����a;��n3nĻ�s�%���A�_�
��g�A��lݎ���܈��0�n���?a#��b5�6&r�ˡ�Ԁ���d@�A�3fX�� f�����fW9��笞|դ�������g�-h���J�\��������۫jKy}�a8x�S�%J�i3:uđ��j�x��pE�i���qҳ��ܕ��01�CD*�6�q͎~������B��s~�+�`��)~��bWwzQ�"@��|:?>U�3-)#!�S_'Fr�i"|���z�.E���if4�D���uW�nZ�����XgzmDtp�Zd���8�� �߆9AC�D5Xv��ig,�����zk�J�?,�VW���l�#Bb�B �?�Ӭ۳�`R�ͱø	��ԡi���#�_|}�F�y�=�;"���[f��Np����⬾pp߸g9m&��FQO%�[�h��+�2�����eH-D�!�=��'���Hoa$%zg(���~��u���^f�
��&�������ع��rW�=5�$ǝk�@^*?�v��R����[�\"�G��R��OG��s�7*�/���_U�nF&{�|p�S/����(0qO��H�çY�|���ʊ�j��ìɹrF4緋:�z�Zm�R����ͣHK� Vjܲg�c��eg,fU"�'�(��|�yC��ЬsE����D4��KZ��p���di��{�����2,�@��J��_B�"���H��ϰ���|.��ʂ��-�����-!�3|.P ���o����J��WQ������M�U:�Ua|�N�X"J�)��a��ɴ̳�F�@tΔ^i��6�y�cV�����ǐ�!�R$�qM���s���[e��s�֤/�?k[�j��9�Ꟈ'�$~C�,YD$��n�>.ڙ�y���8n�^>%�搽��0Y�w��.թ8�M0f�mHzK�!�kIID� �%?ˡ�tz]Ş�[���}��SFpuw��ƺ�4k�1,g�{d�e��^|��m�eH�K�%��5�2��S�y(�.�py��hd1����*D�h�U�%�kc�-rD�Tc�9����I����#�T�!`d>����`��6��Wvf�e����=x�{7�/�]��1t]Ǜt@N�M��Ia��dx�W���reL�� \��%��c�^�O�qJ�0�#:�K&~�1�����ű����o�[��9��/�	x�F|c_��^�g@]>J�iR�����=�kZ-JC��H�n+�i1:)˔��[߀��ɇX/3��X4�r)�2�~���_B�e�IE#I|s��(��?y�N,�ʛ��uX���H����z�����{�G�減��O�������􆢂�+�䫁��݀(�	b���Dz��D�R��#ի#Q<=c*\��֨3F�2�����)�7��,��D�V���â!�mB�n]���=48K�����b��U��89����[:R�-|�3Y�}���O�cDPv7�_��
'~��[��
�H�Z�s_��;�	9v�f�Ql4w���<��tט�U�F�i�cWcO�f,e������67��6�"��jش��/\4����������n�Pe���L�I��1�?�G'�yj�B�h	�5�q��i�U���8�L�$��>���c��=HWE��c��M�O#��u��,p*�WW5�z�y+zȖք2�oP��9���
v_]�ֻ����k`�#�<��AZ3�FmZ�U}z��b|y�Nb_����'W=	���Dh����1�PO�(�Jʞ�JI���8����{6����|,���_x=�#�]P?����l�⠣!f�l;�;�^Ԇٚ��)�C�KNڣ�c~j��+�|Ҧ3Ӻq����8��V&A��?b;TfM�����|r:"�wU�mp��)x��غ*��Ue�^�p�O~�l{wi&���usJ��u���#[���M��lߖ!���d�}��fz �����%!��C��7��D�=�9�<�O͕�?jLyVu��0��o����*��ȕ�u��ǵ��S���ߕmk!)rʚP{|��_,��mhi��C�X(!n��6�B~�_����O.��;�R���P��y�A��;��_C����k_@T0Í*Σ2���r�a���u��M_�$Kt���A���.QU�.`xm�E�2��TdEu�[\���f�9o�`���Y���ɒ�%�/'��B��U�u&���iS0xAe�֗5!7R���7~,)�^� X�[+u�U�76	��%��Ӌu2�W����ҫQ}���}r$8�N��w8Kr�G�"���V]�����ӆ�K�\'�����[,�q��ºo��oc|h+R����D����m���
_�Gm�ȣ{��%�����-�7����_D�71�ft�S�Q�|2�23�&'���K�w �����ZB��"����.E��c�ݡKD�N���Wļ&���J���X�1�rL�Hc��$/�zò)&�{M�v[��ą�o��х�)9��2je}�}���sߗS������B���Y�kp!�7�Ųh��w�w$�I�Z�߬�
���q�u:^�;��z��b�{2�1 ؓ[�:�|y.8Pf-�_2&Y�Mx_Z��u9H��j�:`�D����ǂ_m�]p�9@���������4;?'���K�fh�~�'Ъ	"�����E�_�)c9���ʄ$~��P+�q����3�����ͨp�!�g#()�IcE���BJ~H��|`֕UG�����,��7�C�ELZ��_����+7�5�QD/r戁i�ٴ��G�:�'� I9������� t�J�@R_U����.͝Ni��7�K�K\�8���F��5Q�z���NB^�!nEË?���L����p��Wiэ\;���]�a�8����#(;�'��M��7���+�֕���D?�DE+�:+�6��t�����eƬ|�Uvb ��Q��C��=~�i�ڥ��������\-D��?O�S�����&6��}�by�����>�YHrq��P��%8jdņk�A�!�U��v>1�!�)��S�,.�/�m�n ��;eץ�Di%C��&S��nw���2r�����їݮ����7�~5Wΐz}��G���lU�JK��3�'ex����ψQ9�0��X��6Ϫ�h�%��� �/�σ_t(��t��"�)C��ϻ��p� �݉��;Ocj,�B��C�Ή�W��V�������`���x�ǢD�(߈�\|7���F �Y</���t�|���1\�_2�Y4_����uM���gG;�z'�?�������T�Ye\�-e��R���q�LV���������^3��2Z�i��5i�4G(҈j���e�Ä��������@5��6�+��H�����#����U�o�n�a��b͌$�T`�g�e�Hq�|�H��� ȼX�����I�Ē��.�7.o��=dG"�N�?�)��c*�8���y��H�	�VO�6��
�B/����A����ۤ���F�A��\�lI�g�ǝ�̖���z�b�n՚�$���r�&�jc������{ɷ�Ǽֿ�	��L���Da�5ޔ� �0rS�4s`|Ǳ�h"�{����8��b��ug��RC���B�����.���J���xG�{ҡО_��3'P^�?���>��H!kf�(���ARbU`�F�!�ߴDV�2����� �1��vP��*M�i�H]�6���O�~Ӷ��u����AL�S	�w�a/c%���*��5���l�2Y\F<ue��������ܙ�^`�gT�D�#��kW���j��IZsv�0�xe_����7D�4�"0cc+׋����1cIeǜ�tfz���bs�E�������$h|�4ϡ��dS��W�j��^�gp��ߖ�h�����1����4��6��?�4�����������w�����e=D��*�^��e-���(k��'$E/�~�#�?����)��>��{67G0>A3�
��/����DG�В.M94�ؽj^��D�?�=���s1xdU�z]�4$b��c�y���'���ʨ��x^�פ��l���,4t&IA;� �r�4�� �+��.i"��Wo	w�,J�j�q1��(-��3l
)C������W*��vэ�r	u��iU6�^��m�P�K�O�R8�AL��a�읡R���������˛рJWӟr�u_r�@z�����-�2]��	������T���A�g`3t����F�EЅp��]�pn�C'�ϫw��؆��S��/w*�>5�!�6�]��]Q��� Y�.,Q?>7V�TI�1��tE�����ۮ��F�����Y��P��ƶ��#N�[�ɟJ��w�`���*��R��Ϣv8�M��QѠ��|�  �:k���_<o쀖���]�G�	|�{m����O��Zy�ֿ��F�-Ml[���ph�$--[�)A�l�G��íE���p?%T�)I��_3���Mf��qj%���*EzW�Z�%��a�2C��la:��k���9�����V�|հ�J���6�g"�^�;|��0��ăn�EO��[tn�2+'��
T�܃�ƀ��juq�o ��G�}��_��NG����=�?C�@o��:aa��[����Z���I�[�<,' r��$^mM|p��q\E<�br�ά�d�u	�	ٮ
��ի��M�EG�LY��'����=�a)�7ڲ9J��Ţ��O���S���&lш��J���lߜ~GD��S���� �(�w�F_��H�'Nc�W����^��ڳ�J(>v��΢�O�^x_��l_��(�2O��U^A������c�*n PNH���f�c�9t�6khh�I�]^K��<��!�?�4]�I�3s	0���VT#n����R�5�{���2�o�wXv���]��+*�pJي"��8{gFޣ߂~@���?F�s�L�ɷ�ƀ���F��Q��p��<��0xn�|!J�Y�����v��Ԃڊ�r���厽��xL�k"Q1E�������IN���(�Ċ�>2w�&;��Dx-V٪��.���ز��B�

U��:�N?���4y��(4xN� �O����V��HDm	�[���-��
��M�Bre��!)Hj��Z���t,��HpsC��B�ߨHSuj�?]>��V��� E�4��&l#�>�Դ�\TgAj˩�{��f<�c�2�vI("�q���:D/�ƀ�}h��&�s8�}A�0$7t����f=�OAϢB�O4BAw!����L׽�)SK�8��)�vi�r�4t����q]��֑O�����,g�)�?J��ϖS�(<r��^���<j:� ٺ9�Mu~j�?�/��3w��B�w�> >��U+�Lx�'��Ra�"��!�����'�nw�p��G�S��	��bF���Z��%�K�?lO&GN���؎���e&��m-��I�颂4���Kj��+�Oj�B"t_A]G�^�+�<`4�L(�Vqg�*����\
Zu�a�����`_�6 ��Ӈ4��!�A�?^ʘ|��
�[x�b�Y]��H�J��љ�d�?V�J��)�U{�.�ͫ��ɛ�5^]K�P2m���A�s�˘��z¢��k�Xk���ڦZ�I�Ǭk�����z��UÀ�ܻ��Uw���\dXr=�$P��M��uJ'C7���fO�R
�Y���Vp2�:~=���؊<�7�n�j���������|�����a�U|��&�����W���4e��o�FU�O��,=<Ls��ߋ�"'����dE�/��f��q�<��
��M�$�~��_0��z�Xfl�ԩ�r*�6ܶ$6�cs�⁭��x1��C�=]��?!·h��ͭ��9`mvt_�q��4���A���5N%�r�;ѥڀ]�(�Vr�E�$�Z��ĵ��m��SD�T���+&��i���G1�za��j���V�k�ҕ䫕��"T'��_���<�Ha�W(�ɶ�Hx�׵��4K�ZW9�e�4�b����ۣ	���±�����,ch�_�ga�!���~�����`�v��G��n���ib��y$}��V:��Љ�8��i&/��|35)b�8������q�S��)&���n�u�h.�3b�&jY�9O����M�,mÿ�KS���F�[�J��q=�us{�,}SFJ5��ַr��v�~�K��us��<C��D�Ze^���Y"��]<��1%eg�h��:~��Ke������	���'�n?�-�xS��e+ �!��:������zt+!�D�?�<QLOK���LM�]����",)jpS?U�x($8LTw>��/u4W�����*�CO�%̀f���Sd�g����\e[�K��7�����_�ea�[+�}��`.y�����>�Kb:ဌҴ��A�"@���.w(V� ]^&���
��a��ˏ���`9��`~�B��U���^�|Q�2�W]69�#��K�h���N��]�d������ɕ�����)"���t�����H��R+g�rQ#IU���Og�F�>O�E��Ĩ:�&�7�|�X�r���e���{�'L:�qBS.�5o�9� ~�~��ɮW�@����%+�INC�d�B�Bq1����);�1�񱥓�e���Vt��i����.��h�+��' p��Y�W���mD��B���$�8�l[E���Mn�w��6P)P���ui���J���y���gJGϥHd�J��[s���s�z� �0d�mNȔ�H��`��}g�z$�Ll�� ]��}QoU1N��2a"��L��$�[�ꜛ[�GW�CrL�.
�܃/CS{h�R}�tA�����?����ܚF�;}�ې��b���D��Jaԁ�+��MrD9�r%Wfnq�dcbŔaw#��J�Xy�50��_^�Ӽ�������6�����
��@7��|]#"ܨˡ9xP�9m�F.U
m��Ή�5x����Z���(_��n�
�hVț��掙A(��I�"��2��E,LK:���ID��PQ��>$������5cZQF�	
g�q����A����
ӝn�-	)��e���?au�۷�4�.�>�_����=�&4�G`�vxb�+�AQfz�� ���Wt��Z",?�yn�䉘P�W�vl4��\���?��r�T�i���B���y��F"�bVo�LT�qP�_�d�����Z��������ّ,�Œc6.�ZSq��!�n�Lc~ª�~�W?���-�tpG~g�55�Л��mRXvVF����=7��t��`Ϟ��j�S\��܇�7S^��Z��حy)�&|h���U��D/��hP!Wb/�>�,�l���� Q(�q����9��>��aKM?���o_��*�]���̢�����H0��;:�ۼ���KP�կ�(�rʈ�a!{�������F�Pot�xH�vH[=���~�2��P�,->舯�z��W=FA��GfnL�]ow�)��W�:�Y�/�&W�&�m����I�Z��ಳY�����Ҡ��i�5��^e�����\]���Z^����+���g[jӭ4'Y�� <E)�ȋ������A��'Ɋ�5�j2?�^~��o��|��w9a��Y�"��*H>����?^�h�3CP���r� D�6��:�j��~�׺����*|Nnw�o�7��R�;Z|h�Θ�ɐs�K؂�:C�)���,q������k�\5�/�c��/q�˳OYmc�m� O���"Z�s�e!���\�ه�����´�d�K4���uV�̋�jt���-%Q���Ec��,ۊ���Mx@�?"�%�#�:5O��Uy���'N�ٟ��������^ɠIK!۱"_�r[z��mȵ90�\�S5�gV���b���ل���{������.d�;�-��[h��bf��1;�Q1F��
h�����!>?�a �B����ņ�ި�n��ƹ�:3��F#+����]t��ph92a0Pɡj}��/8�s��A_���<�Pa���Jښ�D�:AJ��	��)����	��9�q)�d}�/�� ����Ag�+����t��!�~�9P����7\Gc(��K8�Ȇ$n:��g�;.����(�K)|���G>���+��pyi��&<▘�J#���l���t70w�3��na��[���*�1�У*�.��Ŧ� e@��m<�>构�E�� b���>rrP?�	��Ĩ����´噲����pT��:��W,�$�'>		��~������f��"�W�>a� �S&^L�w?x�W���o�����
��Hf��3�!TV/�ռ
��,���Ƒ2�A�����%�������ɓ'b�>D�H>�x�C���:��更���'�^r�j��FeX�l��K�ъ��0��IQ,E���dK|�NWU�1�N�Q�T�E��iU���LD	^�[�9�Xx>Wp
���� �!�F�/����[FU�_E�&a�MZ��h���~�i})p��g�����8�+oj�ߜ<~D�?z�����Ҳ�2q6�����%3"䗠h�F �q�O�C�;�0Q�9#h��,��T�"��2g��r��c��}���`R�3	��s�:bO��qJ�R�����p�\�vV���@Msy�8�,em:(��ME�I�s3�Dë�R�I]'�1��
fT���?�i�<���S:z���ٔ�ÉI�����,{�F`�<_�՚28��pGy	�T ��RO���*���s6�a��gp0�X�hv>cZ��"ӆ�4S~�L	�#L|k���`-!i�ny� a���&�L��b�_,�]��'؇��O��Ϗ����>�~��������
C%������X��_��+����s8�� s}	Bq<dcf�v�0��� ���o����T �(�߆B(^�갗ı��j�O�d�b��9Hs��oEh����a�J!")Km�C��U�{�5m-$�oK;��M �6)-�����QX/�6�/J%oUgE^`�]�ՂB)�p]Z�) �R�3ϝ
ǒ1j��>{���#�������K�u�Bs�Wz�<KPa=��X&I
�rC)k��^$�*�-]$U?Ŕ�ȡJ� '�`�@��u"mT���ZG.ߐci�!�L��D�=���$I�*�II�f�c����N�L��%>�Qj<?2�
˵0K�1˯�.`SG��b�ҧ'�S)<�,hy��p��f6c��ā�("DTG=)Ia�B
2n�s�#H����@ +��އ@sjj�)��4A�)��5o� ��>�K��kQ0���R6Zz)�Q}�vɕQ��̔���xN�E�9^?$����P�>�)���D�GR�
u[�E�cJ�ĚR��������H9�7�1�}�hG#�>����+��B����|��fg R���9�NB���o����2���ȅ��<��"[�@;r�O��r����#͔^.�4�E2�����	l0[�/���	��xX�����;����D����Z�v˴h����W�-��X�A�rAm����T������Zm�{S�|��j���{ߥ��h�G�S���ׄmt�C�h���4�>b�D�P��Dl�0�MZ�=��r}f$~+Mj��Q]hy�
�r�4�3Jl64��dG4beo4��Ѥ&�%Y`&BH2zlK�$_���}���jl���E8*z7�+I������d��bc+�R�)O�{#1�����gk��UJ	ߏ���Z�b�5�J��mI���L-��H�I��V5F(�!,��;��٨V�"�s(T����gS��u�M�!���0�����u�k�E�ľ�)��},����g�z���ߥ~���r������������4�"��z@�M�6�g	n��?�����X$����Dv��1�4	�����<f�����:�����#��D
b�l:�ʢ�|BImP(ml�J�H+�C�Oā��l��K� �E�\4������Qq<����M��&&��U�~S+�.J�ۯ�me�9��%�V�5O��.�qj��Z��W@P������^�2�yF
��O0ONiu|Lv�fPfi��e!j5?�(�P�b�[���F�\H"��G�&�)`��PF2����R6������\�d�MZZSZ�J���T#��bN@�G� �:�a1��O����I�#���*S�v�WN���&�ڐ��o����tY+Y���K	�t��9���Y�~'��� ��{��,�� P�{�.����  Ԉ$���ɕ�tk$�C"�j�I�ܩ������ך�3:�A{�Rؑ�Z�\I�+��I3_g�Њ����§L�E8v�ۻ�������˯�/�ogiz=M���w*o����H�DCh6j��n�z+:E��:,|4(��6�XJ%�c:D�r^���=�Q��x�C;{����C�L��R�^�i_�,A9��/sP�ڦ6�)��x��7f���
a��T��a�m����� 5h*�Z!��&���� ���cj�V������3!/��u�w��N���z|��dV���E�!��JO�Ci�oT*��H�L���3IF;@�(����U�������}�0"qhF��|>�Ѻ�T���g>l�����Έt*|�A���h����푍H��Gy�Rg �D���c��b�5�&|� �k��YL̗:� ���-)`�Ե���!�(�������|Ր#e�*ۊ����GQ��=/J�-����
%?��O��:H�&I��iG}Vb��>����=e�834�*ZK$��&0 *1�m���JC(id0ָ�����8�~gZ_���I6���b��EZ���^�f�wy���1s��*sW֛�]^������>_���pE�?%����^ē@ 	��`���
�(����S�̃Ĭ̥0ރ���;��c�1�+w^��7o���qXԡ'B8F�҅I��� `�0mAr�3r<��H��2�~ ���Ѓ��6�[H�ռi5
R}��������"jz��]�"��|ۿij�͈����:�'(PW��u!�H{%&���݈y��''TLY����ckh�� *�@ LeT ��F���ް�t:�~!�!�8$�V�D3Yu���J�m#�ma�ҌBpN�J�.�r%P�
�πPg,� �n��Uw����i��G|
�jZ��%�9W�Z��4a0 i�����T��/��x�j�@���kH�����P�RN���>O���.�����-ח�� �@#R�t��_�.)�5�_Cq5����x�Mf&�gU�ر���R�va��� z��2��(���	R/-o��:&}�'��>}���f4G�,{uv�x�l6����o��;yQ�y�Ì�P�f��K0���L�#�f�v!	lD��B�(��/P$3-k�v�:G,�3�Ʊ��eko��lA)OLH�G٠<wV��/��~��J�y� 6�tE�~�:J�ܠQd���Ne!����-�6_�`p1)�"#o
��_~�V���F����S0�"���p)^�
b#&���%�2Kiq|L�z���&�����)�����6x�$^������A�;v%�ɏA-R��i�Σ�D��g|O)�Q��9����v0_8[ikM�R���<q�b���'�ԔL~"?#���J}R���*[a�����}�����i�������0���W�-���hf�9��,�YH�DɕH�@I�h��-�K"�u������W����A�;p�8iڌ֍O!���ό#�H/U�� Y3J�>����ʖ%:��1��,k4�(~���KN�2
�a��w�m��6��2��Z�^_�V_�/Vo�����٘����Qx��;2�a�I\�������i4�P*��8Z��]�~����_�J��4m#�(���dc	A���B�H���m�0)d��%�sQm��
&�*�C����4��A��������2����i/�4�(�8�VIg/�Z��p����KZ�$4!�5���f����H����.@ISp��g�:M���4�N�F��4��}@B���澬����gT��sa���Y�@x)�=���>���7��H*2�3]4����ג��IV�֡���D
�=�g ��J��R%h�\��B"�籓L���--f{��Q��;���ٷQŵG���Z\\���N�\E� �B�ʤ����)�u�47O�J��h��t�(������]Nz])2�QQ &�Z���͡���Ŗ�(�� �g��6�C��/��	��QQl������ONO������ɳ+<y'�a�Li�eE|��u���pW��E��db�:99��7!�	�l��F�	���Sd��?�B$�*j��$��Ak���|�` Қ3�hTs����̫J_&��D^��io3xk�h�ˑD~/���qy� �Ř|��P����R=v(��},��$�5������f�gԓL�Z$]��X�/�mHћ=�뭾�`Λ� U�4c*��F����1���>��gT�q��L���J����p��H&8<�}Y�0OA(H4�5�g]�N{R���SAJf�RO�pF�J���P�Xe�?p��i�aRkq���g�w�Z	ٔs9���q��"�kR�D���!R�?1���43]���j^Z��f��6��iD�|
��ZD��G
b�&)���שy�ܢO2���#2������7�|�����f���*^]��;���f���W��_=��G��j���p�X���8��hv���ݼE��K�i��*��@]���Jض�G�~!�Fd4�n��D���jZ� ��=h������!)�m(����l��^+m��J`�ֽH#�>�6l��NE��F�m�j���v�kMN�I ����VkZ�Wjza!�Lp�F
��4�a�}Y-X�T�G����D2p��GB"�Є'R����l�o���_Ң��@�/1iEZ�g@)o�I�"�|�I�����F���:���q�����]��P�\ǵ$������ ��gC$�C*ﰦ-#����4*��>k��������eG��ա���}�#)3�L/r��4��o���2d}���цpg��)b>HUT����@���Hװ�0���1T���I2�~�ɴ��B�m�&���d������� ;�l�w�����b~�@��z���zu��j^� �8��=VƂ^�ÞhX�e��.�sF��l�|�DsP�3
^B�U ���"�9�}�����W�D���-�w��79y��<�k��_P?�?M�F]�e�ZoF�X��/wA�ٶ�i~�v��D"mҒ�RA�NvɢDE�L�V����O��n��H"�
k%���E��I��~���a}�p(%�!�|�D{k]&d`���0��G�`1��Lլ����8d�0��,e�����*�xAYY������*��Az�V���E�p�hA��>�H�9"M�r>S:��D�#�Aҗ�!� ���X{k��D��K��.婭:�5?-��d�4�j2V5�=���yg�h�X�/�i���9"�<p�-�':j�R�`����U|	����/0�C�l�@�����f6���ڌ?}�;g������$��V���<�ə��aM8[j�^L�~��~��Fd���NMءCVu+�{G��լB���VI�nY�B�����+[our��fH����F�4����(`s=u�[��_�Ǒb��0����9�k<6��dFk�/�`F��kR�D�B�4�Xη�����iK�e���:���f[{Xu^v�����PjIz��J�,�q�챒І�|�Q���̓��OL��&��~5�����d�K��0*������%E��پ��,�`�v��ZB5�h\V�QP{m9 ��o;|#_#*�4�I��Xߓ��y#�l!Q�����޴$c��>#9_��D���6�*��'�%o��r3ٟ(u�����kSl�p���g�N�ˬ���0�hk�,/i0�����3F�0�bR_@(R;s�AA��:ɫP�Դ�,��8ݤ�Q�F$�&�*��H���c�q�!�~j!yfH���P��<�wXڭI�Ǉ�nG7��{�勢$�	~ �C4o�����y۴ SU��o���H�T�&��e8�v3�N��P#��eY�hm*�Z<�X�W�U���|߆F3��/��V��F7�;��fS#�	Ү �>aJ��zJ��!Ҳ�M��`��9��ښB�Ҝ������D���Wp>H�E�(/���?�g�;�K��.m��f�5��/@!h@�b��!�e\t��M�P�q�%L��0��z��4Aզ�e�ѧE�"�1���Ϗ���t�o�nT�"��WT�0������eN�gSJ�=�mr*i�S�_� �ڸ��2-� �Fk	�MV�23�ΕF�l1狉d�א{!�n Å�����z��@v��[c����9�V]�9G�m���`D� S����L��4�_"��j-j�{��I�[*+���FJg*�/}��8��NDꛎH#������4�#ߜ�o��BK����r����o���?�;��)(�uN�䙨�:�ϙ�Ҽ��`	�U�^��伉$yYh���j�a����� �`���u��h�S}E�M9ͫ�k��E�;���%�I���S�G�WB�EjLq�ٍJФ�A�M�,�>^`�	R��K$�^,��{����{U�C8�'��K��L�V<.��
�%nE]�=^c�#�'���P�`��v{���x3 �J���` ��-�B{�߿ z(�4^���]8�?d��sA���Vc�/�&l_�v�����2j� ���Y%�qkل�7F����6e*oJ��U�$��!@���"s�\6�ݥ�^�R;�Z�4r&�|��R%f�(バM횇`SZg�!�5���+�h�s�V�b4��H����t#�p<��I�[�X�m��W"u��� 5�P����T�#R��T�I��)�H�j}E-#�Y�wHi.��-�{��p�����9��)PbO�&�Ւ��Q3?�S�Ne��E�3u�r�Ύ9���f�����O��������ɢ��+�'b·��O)�lD{@�*�xkeI+5h ���ژwBn�m��z��63�� �-#DK�i���ئ�ț�>[N�����F�$�9�I��C�P���1�d��o�p�.\�&�R�j"EE�f�+*c���5�I-,�"50�jB��T'���w�Io�=X��k�}�Z}��y��n��Y��]�7uq�D��a�N�r�9���Ѥ��GBS�jo���%ju�(���s��j�ʛI4��Hn@�DzR#ܵ�jL�p���H�fHh*���=�gSz`�n^�m���n߃�#�t�&51�v����J��A���7�� ��)�sv�&Ŧ���O�:@���E�����3����ѳ��^W�(��v�.41MR�gYNhΠPKE��3�nn�BF�a���ք*7��ec��l���݊��2-��ؔ!g.I^,d�Jm�^V�f�Z�A��Ʉ<�`��q��m��#���I����vi�QL�&u�yu伤h$y��dk�%LF(H؀%�t���"�����᛬\pZj��: ��N�y����mˈǶ�����^Ɉ�������Mr^�y�{wOϊ�2 v� I��MJ�%9���J,ũJ�|J��O���o�/��R��rY�,��8vi!)��EqE	�! �>������ܳ��Dő,�xT��gz��9�s��<��d��G�Uq/���??��qp~�ќ�iF?3J;�i�R���Q��m��cBs��������k@�z6�10��)���>���?�QE6����4?#s�ٳU'�b��'DHjG���a�q묡��q��p���/���_���_�v�س=�w�����(d8�F+�<_�'^ǡ� \�}���:�iK���!�r�Y�Q���R��S�,ut����10�k­[��4�-+w�s	�H4t�O* �8����f+fURg^?~�l"���@�W�o��S��D)P�{�%%
Bt)H��O �,�ϔK���f$� ����I�TZuz*�A�5�誒s����p�pR��`>	kŕϤꐸ�5	�k��$�Y�V��$�H�d$	���&�׊e�q`L�R��]B�O��9e3=�m�O^{a��5�"��q�f��nm����U�D�v����+�)�D�I�W��,�;�,��Y1��%�	$&�����mJ��<~e�_Z\�;�7���7��Щ��^�w�����lm�xd���_�+[��l<.Sc�X�������A*���'�o� �ՙ�UFF���d�x ��u�&���]��i@�!X��8����I*����(~�zrR��}	71��\@u�f3�ƃ[H����׊��|T�����
,���n���8�e"���ڈ;>*q ���cw�9q[&t�lX��2&�XMO�J����������P5�>���*ǼmhQ�n�0��+/|���j����N�y�^R�,PC>u+I����yB I�Ԁ��A��
Va�;hxC��1�k�68m�S2FՄq�m$G�2ա�J�?����dP�R+����f�LF^�Vӄ����4���Z��`�Ң�ÐYZ8)�(�`�Ճ��<~-P���_�S��|����^�����x���2a������h]E��qY�+��p���>��z���Y�f�M����� ��@EV��������,O>rq_��~��C��![e�As�uyJHR6B�|5q��/b��y@�3�h�e��}��n�M��PQ�d3��SwӁ�`��VN��o��Lm7
�&�AdH:��[Ģut%1:���)jőp��f�U�o��0`�B�C�$�i��%�g*�����r����ޔlK�d�1��2�rO�'?/��K<dg�S��W9�ż�&o�@N�4�I�&��h*����|%�B7 9�k^:sD��~��BO̄\�P��Z��ǀ�t&�(ig�De��y�NwJK���M��eoػf��~��	�����#�q]n�Ǐ������p����I]'�Ѩ��^�
����Ʈ�,���|4�7.��b�k���[׮��=�9�i�0xٍO[؂ѢSC=��ܠM������ Q�?�A�(Ɠ֕\?8��5�������[���[��90H�l�]Y��{v���7�� J�k����5~ȧX(��B7�v{b.��[pAz�-@(TPqʓ�����0�$�,�I[$��C��I��`��y���()^0tOw¶12���>_	��Ң�
�ϛHI2�
 H��2h��X�`yNER��z˾G Ӂ�q3(J�,��%d��h�ϐ�f��ĩ��"JpԆ
��'-$Ң�%�ZU�V���4r�@S|[�f�ki�5��]�m�Owj�����(��5���
@�8����b�K�XW��p\��J�����#�7�W��i����I��Qw8��0ˉ=�1XL�F1c��S���C��r<����6~�OgL1%�,s�����>ϟ�������P��Zb���kG���勀��l�(t���Іtr0Q5� �D0NB�rm,9��L�4�)�����9e�H��@Z.,As�
���&�� (�6!T�C�qo�bˮ���Է�MN ��vJ	a)�݁��idD��P�e~�
��%)����@�di���+fISaB����7l����n�nஸ�	bfO"PS��Y'�O�n�ΘdF����&�P�N ����F{q��Ze�>!x��!�(�ř�����^ݼ������8z}s�x����������l��|1n:e�;���C��#l������"�?>�Q<�&3��r+"��a(�D��|2�Ei3�<��}�
�ZZX�E��cp�gg`��Ϡ�%�_���MS2m4��3V	��}��)<�ک��;��煂�pu�*��h�ʬ�@�!��hO"���[譶=ŗ��q~YM't�ÏQ�@�f:��Q/-���7RF���9��q�N�H���4#h��(����:AM�J��l����kH�xS9����T�4����g��\��6L���3�BU���-��K`�)�&JF4a�R�a�!w�n�$s�u���>!x��x�?�0^��'���:��|1���ޠ\͋�J]��M�o�oޗ���q1���kΜ^��4Zy>��	�[��t�Jk�N�0嬻���>�[\��#��艀�kd�c+��K�w����kW���&va.m�)8Y�Q;
�������O.�]�{��Dt�5��W���)ָ��dvb$�au���58;~�$ j'U�1��{ה��8�â��԰g6�!�����/�D{!ޖVA%�*�	Qx���S���iٌ�4Ԛ	%{|�w�A�PD�MD�S��w�b�[]3!�͂&��>Lw$��Dm;�P�i	d�AZ:l�W�`9	�uG���Ǧ�S,끢�s��i[>�6�'�{JM\t�-&��]p�c+
�Cb���ȡ;����ƍ�}�aW]�.���q����C�6��6���=E�k1!N�S��-�L�\���d�Y1?��.̞*P��ޟڊ`��#�B8���6* ��B{zͩ�D� ��𤄵( �"Ig�򒦛�,��9̔�`d�+8�x�诚����n��Ӡ���Hl�[M���b9jTƣ����!����@`_�԰a&��@��eD:#Ԥ�ĞiX�%)%�&5p�<�bcIBȮr!�o8�<�X�z�D]�%����gz�m#[1�k�,�)�tw����$�V�)L�zf�7�Մ�Dm,�`����Ш�}�+�߃��;PF���񮄴��-{r�Si��*@�@�7.��r�R��*�q���hlR�c���i��Sպe�Gj3��%�0G̭�).� �c�!�Yȯ(��|��b����9|?l^���-�C�ͺ?g�o�O��J&�sR���#wƥ�R/�����C0ERˬ�O�du	�����<H*/����yp�W�{���B� ��B����}Q�����k*d�{hbJ2���3 �)��e���,8�B7�%���C�R�Cp��zƶB�u�	����x����:"��p3��Ќ�~A&��:������,�G�7_/ѣ��w8�5���B{��+BԸ��	���- |x�2���}6��}o��ͼ[�˝EU�*�z�}WQ�6YPe�<�gO�ݦ�i]�4���:#w���AX6���of���Ft�@k�{�=�QgN��7}�;׆��A>�6m~��� Em���Vzj�����~0�go��3�~@T�@F64= �`�����Z^v������|��!@��n�����04�.Q��{�~����ot?#�S�t����h�Z��b��eG��R~3�h��� a6�����+5��-�a��D!����'��G �)J"��9����U�6TH�-L.h�$[Âw�zռ3N	����bA�8"�s������q�BC�f��rԐJC�۳��L]���>!xx���t���������!�e�aن�I�N5�KM���n��x_��y5�]����ؿ=-�7ڝvL=���.��z9�2�C;	aǡ��a��7�@a��v��A(tI���(�f*����Z�
km�Vפ)B *C��Ƨj�� ����N��,����M�\�4�DOu�KR {JcB�YPV6U|�G3��[i�Of7� n��[1��=�?i���]�(Xkng)i��ω����w tSl�)����XS���`$rX�D��1�5��(��v�(�J�@R��G�}�]�a
&�ԾI e�n;{9[�|B��۠n�1�����+*�5���;F�V5����y��*�FE�g<͕���w.������K/%;�V�m0�a8���9+�i C�bR��x�mhlR��m�q@{|�'f�����eV(m&��,���)=��u����p'��4''�.yn��MN�Y��ۙx
#IFIB8��!�A'��&�C�E���k�bP�?��	&�y�L�������fd[���dv��yr����4����3"ְe 7�ƶ&i����.$fQO%oi{��R��*� �>!xx�A�$��܊zQ�ښ���4n�]��x)�*۷�\޿�7_y�{�:����7;K61��g�-�*Z���%)$�t�\GBv�Gl��i[%ah&�ӔX4/�q��=����648�\��U�&���s�� �� M7�gY�b�)��B��)u�2��h��1��$��Bu,���#{�B�b- �n�\G�ZT���Md+��Z^�ĊN��, �e!�R]K��Pe1P�<��d��iUh^�^K�2ݲIMCwq���
\3�������r��C�	���p��ٚ��������?��'�������?}��7����o��\��1��OUB���o�t��A�s�Xr�'��L
�/�3s��l*�������01h�"�@��3-!%�I�^��B`����<9�烽{ga*��8�ա��0��|��r��5���(U��`��r#�$"+B�qNb�!Y&��O�&z��+�9ES^:E��K��≞~�9�ICjL�DJL�1j�l����6魔^���@�m���5I���J�'����'`n��!����q�@���M��_��˧������N�:���խ| �Jm�p��tcO��~A~�s�(�앢����ڤ턛�Dդ�ĭ���	�@ǺH"� ,\GA�~mh�Iޱh�?C�������X��Rr��5����)�ؤX�c��5͚A�H0��7zir�	��e

��c{�{%G����
�L2��<�"�n�3�g&��34��A&S G�L�f�H�W��(��4��UӰE��"��`K���s�oJ`���>�x��Bku��۽�6�<<�2�n��<�9��G��������Ͽ�صs��7v���V����:������`]Ȏ���$����"��u��iCZP��M`<1NǇǲD)�j���[�vq��Z��*������5���4�A��!p8Q�Mi�����k��Tf���_J�P�JyӐY��w�i�Y��2|� j�#�l�)�JD��A0V�h=$�*�x�D�z�2�*���hވ���T���4UI�%V2�Z(���ζ���~��p����]a:��A���ڵ�Q����b��;�Q�����V^�޳�wv0����WR:�ۄ�!A^�Q��%��a�D�j1Ĵ��Y��������M��r�T"U��Ike�(�&��i瀤��R��Ӡ<b-$Ƣa��2_�����QY� �	9z>��3�S�R��N�@mz�h&��ܚ�!4)���9��JRr2�@�(p`��MpU]Q��:���H���Y�ʴA��o$��ז%T%�����߽���	���.��}sUn?���\1��v�����߯�y���rq������m(r=��:7ј��F�$豔�y�FtV^'C��R�,d� :�3LZ5���M*Ix��P�bځ@��+��	oxJ�<�����c���@��7�Gw
j�@�&L"�]6��i�+���T�8�!"�6L'5� yłE�q㚤.d�;bޓ��4dMZ�*�n�mo��P�F݌Ħ�8���6�+ˀ��&UחW��&�w>!xx��خ�n�{�i�u>����Jl��.s��!I�4�vFU�P���Z	�sJq2S�D��=�A.�4MȊ�fFTN��H���a<�E�܁���=�E"(���R�צ�:�����zd�lX�#�7 ���7�a@���a�	yc[dZ7�4��������
�!BV#2.���8���jn9�kܱ(����Ѷ	�&���T�����[L#]B���\{eǷԪ���ho�<<�Q��jx�Gg��q�SP���¹��Q�<�E���4N�PCx#:	G�u��^��(	�@$N:GKφ�Ъ��aF�	D.�*�Y]���,;p��֝Q�VKۇO�O�6;4��jE�$��+v�p�[�[dˎg�������ٯ����o��Z!�??�6@���a1/���@	�6�L	�l�T� ���y���Mi�8�����iD�)���h����Ǔ�Kw�j:�<<�a�>t�?��?��}�CO���������7�t�2�*y�Zi����
�\���\|t��S"�G�u�)�5O�o�SU�p��c�hh�,��i���q+��r�(����J���NH{�D�H'$�Tm��i�˲�؂� �����u��,�z���В��^�S�`�
^��b�m��X�$���.o�*��'��������ui_��H�R�����x�����=��^��/��ͯ?�����7��7���N}�w����mX��i5�P�b\�)6I�eCi*je`b�N�����}�p���<�(B)��]�uCe	��?��|��c����Q�i��P�Fi�
YR�(M=}����M�z�������XI�	��SG��dc�Hє�z4��f�������
I���a3�S�.!��=�jV��C�2���?&/���7ţ�)��ka2hlR��/�8����]��m�O���e�]�������o�w���W���S?x~����� �i���FZJ8c�CR�W�I?�#�:�@L��g+ �dF���0���Ϧ�X!�b\U�c�I{�5�S�b4B�%/�Kt@IA�����ߏ���%�kj�h��f74��d� R��N+���l�c�%9�'�k�)�ŕ� g���(9i�Ad+�6�$�r�^����~V?IXvw/sǾ���)����O�2�����_>����W���>����g���ƅ�{���l�j�Y��&~J<��"t���x99�􍀴�A��&L7G��\t@��'Z����X��ia�'�i���kr0å^4"��P�!65v�͔@0q>�I��S
�NYt��Z!�e�a:+��-ȁ�21x��%.��Aτ�&REI][�-H"z�5�&V:"�Ab����V�B����׾ {oҾ���	���]�b���=��N|�=�����'�?�֌�qT6`�)�{�nV�\~>!�+��M��g�]O��7ݻ�3Z�h.Ơ���(p�x(����qj�ydǉ�M��@��C4tҏE�ɬ�MFRP��pӺ�h��Ш�j ��dg(��RE0i����ʹ��$I�R�׈ELյ����B���n-W��.��v
u��1�������g�O���<<�Ő��S�Ϝx��O�z��{�{�|��+?������STEز-2%D��I��iO�lq[�N��H���yN����0�fX�M�P��g��S��.��	���� �+�q%�tC�Y`s�h��p��$��V	址�@��j{]�,#T6����@�i\��qN�Ծ��=��In�����1)��%t�`Y�e�CA��ѾA^�ٷ�l�#�a�W�}z�����7�m�O.1��������cO���~��s����/<���K�ƽMha�����4x�S=8�Á�%,�ӳ`�>���? �G]E�Y���$o�@���H��-z�8k3H��&n�t� �����L���M3���G"և��"���F6�U���1�� �lRM5R](V3%}%IrZ�SQ6<Y�?7��n~ǶR�mUC��61d�1��4�O����&�he�'���e|���� �<<<&��Y����O�����/}񏮼����qA���#*%�����;Q3�G��O-U3���C�j��3S4q�t�F��rH[��:�(��R��*e+���u���$77a����j �)��ɠ�&�+��E�1̚�	����\R@-!�h�8�VVh?в����]���m��B;���wBY��0:�y�/�Dv[�׎�܎��=�v�Lo�O?���5�O&�7��g��Og_<���a�ͯ�f��8�!�,@�f$�ja�P�&��Y��(�Y���Ȉ=�+�Gk�W�"�&A��h'"R�  <w���)XE5p4WW}4܄B�S��|�}51z�BXȏv��4�W�>�����6�m�;ڱ�tUٜ�`ݼܺ1
�E�@g��{����A7����\{���X<v�Kjm~�!�	����B���jea�������[O���/��,,�&%�h�a�B�+b#��D͆3�i�L�E��/3�}���WMK^��<FPH绠1��i}CzG�����F�L1���)�Mh����%����I��Xݨ�Kf@i5��6ʉ�� ����ca��c���'ܱI w7b[��`��4o2�q���?��	�5�uMsl�(�"W���(Rξ�!�r��+���!"�K�l��(_�#i��5�÷�����y����~?_�OH|
s�ghy0v��j7x���aͷ�]����|��a��C��E`%���Go���V�Q6 ^h��(�ٔ���~Id�D��T�J>���ډ}��ZN�[=O�F\xQ(ȥ)9�6��W������˥^)��{k ��	X�>udLJ���]���ε0W/�U�`h�J�������s EQ��ToĝM�g۝�7)w����	TU�U�\�z ;�$���NҰ�){͙��u�E_=·�+�](F8#+��N�y1w�b�2��-�����MF�����B$"��C�D��H ��#]�Q�_���{2�|QR�(*�q��a�k+2w�J�״���>h��W�d� 1�xGm�.�8&��mFn8;u�)��[��jy���Ҝ:V���
l�UK��Zצ�����M����/�Y��c&�y'�W+�Ϙ��c������~H�����$f��u�IW���7Х��	D,*T�㱉�j�s�ȟ٧!-�������Zo�9���7�EU�)wx�4��ǻ�&:Ox��7"�Pz4�­�C���CL���nC����=>p�i����-��g����E��V[ =�R�U:�m������Y 8JW�-7Q�}zX����o�'����\\�Lo����Q��Ї���,�Y��I����=f���b�FIW��l-�@v�|�y�l4��'m�@�'�E�Z�o�Nu�ȅĒ�s��S�׺�O[��V5�>�=���2|����=�訠�����w_֐{���v��~���.���$
��S�Z�ka�~�9�C�c;ފ:�`�������9M\<ψS�����g�&g[�հ���>�����Q����!.R��y��b�ۗ�k��I$��1X���� �ʂ��#���m	�"r��p����5>ֽgQյj2:��#�6K�o��&5��x8�[�E�|�/��eԙ��zߨ�\t9z~����Z���|4�ћo���m癝5�=�l��m�p�J-��G4R�������y���;��<_��O^M��͝��J��2�5D��8C���{�nH����е�i�p��x}]��6�<1�ek�P�d~�X�{��� �@뱩Gy?�ׂ�mD���O��/���[�K�-+ .���|��
Ox�h�5�I��2���#ַ M��7� ���.`]�CB�p��P�I�(�T�
��o��+	ˡ��?�l��,X� ~�~�a@u�������+����6m�|����3%��eg��ԣ&7�Z��3T������SI�~?�MD|���[��{E��0����{���[�~M+�
�X���
h��^#�7PE�_y��zp1��P:��7d���� q}*�T�\W
δW� 2��Jw�˞Қ�
���$2w���|�P�Z�����x"��z��vq��τ)�ʦ?}�Z���/��!!��,�rs�z|cJ�<egIͥ�݌t�wL�����n�R�S�?� �:�G�v�}SI؊���n�|T,cXl�c��h'(�7�Tf�jg!a0*��P��M���0rv����d߽�?�cd-�[g��!��ks��x����,���$�K1�����G����y��n��]�cFĹ����ь�zͧ�L��P.�x�X�J��V�@�����a�vq|AX2F�#?����6�1�?2�j>)�E�^��	Jͫ��F��W���8�1(Pl�{YfS��f!�o�m0R �@�x��٨gcG�&��Xv���B!�%�P�X�<P>4�q[��UTge%n�US�V��hVL�T��l����]-_�T�>W��Z|sae�8MҤ�٤�i��p�D���_�p�Ot��q���<v0�C��ßBs��B�_�(��P_��ۭu��Ã�N��8��\�]��O��$�Q���ͫ�C۾���6%����p�d�F7oHeG�z�B{��7=a�`�W
�{k���m-�)��݅����_����*�Սz��3q&��N�aAˠ�e2�!����!a�榼���g-a΋Y��+��-���Z���!Wy�2��F��#`���T:a�S�w N��\�L����|�[�Z��mP�y�0���*�GYK�q�3�Ϩ�l�|�~__Wǰ�{��ҫ�lZ�w�<���=��{����>�
�!��)�z�*3Pv�C�`�{�E�TѾ%`�Z�&%���6�QXGG�޾���V���y����@�kL��G�]\�����	�����_��в�y�_a��9�Z3��� PK   ]��W�a[}�  #�  /   images/7a3ae19c-2290-4841-8048-f2fb794005d6.pngļ�WU�6JJ�4HJ���HwwIKw(!���-� �)-���͝������Zg���3�xbf���bo�񑡠��H�+BA��BAAg#�?��pOޠ������AA�@I(;��#(cM��tB�c�c]��O���(`}�F$Rg�I���@WV�~�)[Ǯ�4	Kn���g�E��M���㼶��⡴�U��ɋ���Ht'.?�8	4�\-��ү�����JO���CRp�_��0F��Gġ��u`�篾C!�&�����O eUvY��u����z1�Y}��O�@c�:����zQ�|(�
l�>A�Յ\�?7F�7�"�?������?�M@̪�G�H��Y Ӷ����v`���y������g���p_ɼ�B(�L_��,@p���ηL�ġ'ϛo���)k���O ����l�'NhPz~���o��搩���TU�g�#ɏS�74|�_�KKZFo%efV�kii���(������e&�?�=3�ӗ������u���&�B�}����h�9�LD���2oI�����wX���L�*��2��) ]*2�V��h^�"���%�Wj*�=.#C���Z��`��i~~^��Ǐ����&��3C��cҲ����}ظ�%�XX��hhhb_BCC�A^�R���'&&^�hiia�%UU뾂?��::�p*U!!�))�J��������"�zkѣ���S��,555{/ccc�


۶��DEE	�dqsk1�����g!پY/ϢB��S��{����NL��7��x�����z\������j���j�ⷀ�d��̏��))�щ����0�Hd�F:��	�n����$�4���t�4�����Tq�˵�p��|_��8�*����5$"J?YXX૩���{��� �CE^�lr�v��s��v�0rz,(�(P5���U���0ggg� 񢙼�̏�{J�II�&u�X��4�{�Jb�(��	'
c�#KX3!��-�$D9az�D5c��H��e
�̤�-s�3 ���7M�D�L?Itjl�|jJ��ӧ 6v�g}c����_�ޝj���'MMM�>�"(����A]N|.���������I��ʺ�:���p����b���_:JJP���+}BQ���Z�)�$��h��N�Y�)׿`F��B��O���Ò���+T0��Ezp��BB�|T�\��� %�GӬ1=kS)Q����0��𜙜�*�m畦~�x��7�D��p̠�z{
;q(���UUQ1�3�}J��E���͉�����!(�?���F�ܞ��||��k5jLїA��ˤ��31[/5�����bs�3��*��h��кE��hk2P1��rr�[�κ6:}����S<�/����E�)�_F���������.P�&���ೊ3��LON���۬>��rx���u�;6�	U����	����;T��A��Ϗ�'݁��������x?��\�ȍll��'m��&#�d'��K�N��M&�����|��m�M��]_Yٰ�#N���G
gMA+Gp���,!�}����)}���f������'+��� -�]\�`�R�)le����>�3lU�d2�L�H+re�K�Y.�R\\�����v2U4�bgw����n ��w^,�52�7$S+I��iP,�4������ғ����aa�w�{��O����(���y-��:�U����!�Q1���#�Ī���w���6;e\�o̔�ԙO��&$��|~l���?���qg�h��)RM.�N����렐��g�k$$�{���jV��?+��e%!��
���ǐxQ:��
���v~~N	�����~�G���q����jv!�����% ��W"5�p��^C�hDED�V�V��I%�9�fɘ��'o����s�VŬ�)����]�O�����)��uۑ�����!�I;Ǉ�3�$3�;��\�-
J��v�}𓒑S�O`� �,��*I�\�gee�@���7-�7Eu?L ��y��h�KF/9���3�t�%@/f"qV6%����Ie��m2j:��RO}:W"֩���w4h���кh~l��6כ�U��.�N����X����}�}���bDUA9��j:���;��q.�0�A���ƌA���@��X�0-���L����t��f呋�E�9km��{��ø�����t����?5���7T�����7ew�֍Cq�=Nm�#�a���@9#�2,�¸�yM�2괘���Ϳ��rD}����n_�ɢ��p�B�%uJz�Jֺ����7��`�*/�ȴB��<95U���'���6P)1!z=��d�~~p�`�- ��Bq5Z=_��$$��*^Fuܾ�(a�%hg&�p���"��D�Z�����e��%r�6�̏���j�����jc>�B���kڽ@.������d�J\Jjrtt�B$��?�2]Ld�}'�}��R�މ,�$�Q�o��B��::�|�o����Q��o3���^Er�Sv$Vg7��� ��.�Cܱ3�� �s���uj���A��Ǐ8���A�[t�� 5�*:�p�i���m�xt�Y�P�'��a���=_�������:� �O��U�\s��B���q,$(h�n�� ��czzz��X�~O��@�����ig��j�F� �3Ea�2Scƚ�6k6 ����0".�,@r����4Q�ASX���I�F��(Rss/�ߞm� z���)�|V�*,V�$��K)�y��~@�F^A��)����6�o:_�'��N�� ��a�Y͚ �(�y��������_ ���z{���!Y^C������sP^�[V�e�][���7g�=l���N����*��BD�q1����0�b/)�Qh]��N!(�zBBB���=�����o�����\��y����174�������r�wdD�y��r�򟴘��7i�^)�h�u�/��r��{#A��[b�<o�u�$�V�V9�M�h��q�)	��c��+�
��M��N�<^a�ږ���`GcF�*�� ѯ�$��H��Z�(���o�:6��U����5U�'����s��8w��e���藛oզT���)}�I��
���?�1�5�uF=�t1�$���.�L�G�lF@ꪪ�&�&P���޿T����D� ��0�ј~���ڿ��pP˟� <ׁ�����8��s��N2w�[��~�Fν���A�SK]}^�_�lF;pYe s0���0 ��wAxx�[�찰׏��Lw]]���u71������1�����u��.dڈKv�ޣ�<^�,��r��7,�,mT. Qv�Բ��z]p'3e��8y�s8QTg�Z�HF~�ы�i��w���NFFZ�n�/r[VZ�S�d�xP)�?Va�
ӳ��U�0,,�O�_�W��Z�edF������ '�0�DuE�W��̲�R���\eE ��hi�ڝ lD���j�*}Di)�¿���~`	��qp�mo���J�Ȩ������d���f�~��"<.k��A�FJKK����hHzBBB�BBC��vq����OTDk�g&6_Ֆ���8#�����5�#�U��ca�͸�'|����!�L��?��P8�x@D����p��J{��hu����"##��@k��yyY�Ѣ�S��J�`�e�Z��0�05�`7[32[�d?��"�����N����b\\܄��23�y������/�6��� H��R��x%u0���8 �0ɣ���/¦Q(o�>{�aJ|p�m�e���{�����q�t�d��y5[(�xrvv{�-��4�b8T�&yf=������g����ǚrrr^�S$7އ�~�4u={Ѥe4	�h�F���J1�J�7)9�w�ࠝ��塴���O�;�ͤ��!2�U��D��v�;E��dv@�4��y�ʊ���^��q�yyf�����%�į�Ĵ��e����YZY�}��r��I�A�d�#
�zqc}�h%�gްJ�?>ʊc���L��*�cJ|��-�2�$U ��b�����LL��b"���j ���w�� m���k����:Ym9 n�^��m����\]C#�EV6f�y>�&���o�F�b��=�R'Z������A,5�Y""��5�蝘0��W�B�z���\�9�X�VqO�*G۝d5��r�d�����H�z��������
DA��a���Mlɀ��M��1����)�������vw��t�F��S��b��h�o�b�!���b��];r�x�ȴ��Y5 �9p�V�_�g�s�( <u<E8�=3ļ]��%�[�<=�$���S�y��S�f���i��8ٗ�A��k�*Ӽ1g���`��_	��mVs�zi@�&��K	���f������8��d;���:%&&eҊ�R��Ӎ�a��&Y(I1&:������̌�9)��M�NfO��g�Eq~B�H}
���P�E�i����2��'2��>�cݡ��nY �	)姠�Kʃ�`T̺���'�����յ���z��m�_��x�j����U��c"CC'�n��cA���/�3��Xo�df
ZF	�����H��sѣз��[�E�BK)#�Xb"A���g�]�Z4������VW��_CPe;b�a�h޺:`=�|�P@�M^�*�~+�g���(�d��� �͇\a�`������7�<.S���y,��� �0��̈́{f� V�����ۙ�1Р0��IU����)]�=� ��ޓ_���1h5|2��	�Yn��-O��d�BN&���)ל��%3���!����<�w�%��`����s����(qJR�[�YC�󘰠����[����(�r���zz���t�1!j�U.�/�s�W�+>(+(D�9r�ܦ���My�C�A<�	$����$�#�=_����Vkk�rll�UR��
���Gtc�$��1�<ҁ�"���
��V���ށ -=T�o|&����$��BE��<2P?&��R�8==��|���i{;����&ۣIN�oBrr�����'5f��{{�j���b0��Oj"�"��v@�5�kԚ������=�d��6�]u�������VT�<��H
��(&DP�(�cܽ�?�E >�	�?�VY	�DA\������ai�k���m�/9��Q�)���$�/�cY��G4��N׸�m�G�ab����"I��b�aϮw�Y��8��Fj������::��*٤|�n��|�����b����b����oG�.�d��i��"^��6�@�2 bP�$���/Y�,��,b�gJ��U8��r�t���b&�e����
�7!�kғ<v�U�H�v�-.�~75-���Nf��4�x�L���C��x͍���L�Lj�P�[&���!***���[F�at�A�	�r~~���U�|�%aq�~��3���4=��h���C����<�������l�)�x���cHK��O�FCu /��]�a�yZ������`���L��Y-�᳙+W����TR�d�йҊ�$�k% 0n��$MP��ܮץ*�4ZJ$-�Aٸ�cW3��:�?$�����}�i�O��6���><v�G�;`��,�{��Cq?F���ڇ -� �D�ӯODk*�XpXw�~u{N�>�5���������o�e�D>��,nȐ@V$ �m7�
j�a4��jW�J�5�QFy�e�-f˅��-\��t|��!P�m����n�ā�E�b�(�c����qaaa��^�<��7{��E�t��)�T˦�}��3��R�d����`�^�>��2����|���V������E7����&-!��∏�:X�)���ee��������F��I4�S�| O����)���] Am�b�adll</�H����91��̶mO"��&U���Ƨ䃏�����;���N�J�źȳ��_d��@�����E`��&�����,�v����2�[9j���}�+(��=m��i����Qa��CV�®Ed�$?j5;��l���:���
�Q���s�(Gj=�J.,�ˋg������V���a�q{_�J^�GDA'����\
� 5l3�_�wNNY/��٭���g�<Y}�/t�u��*���R��A��'33st�����<��b�@7+ɀ���F��=�O�F�Ǳ�Y���Yx.���z�v6���ŀ#; ���=���/w;7Gi�}�-�.��D$^��H��Ӛ�N��L��Y׆�o1]#3�Z����s��3e֚��ڢ�"Y21�=��Zs����~Ҫ�	���R���.7���A�X����ŀ,���X����?͋ka�=cu��k}Y*���T"�6��L���7��.va a>RGEEɯY�ef�^��~c-�1�����U��@�п-eee�@��`|yg���xx��v�# �\hH�=d�!#�$�!�;-#`U�Jw�Dú��*���0��)F����ȴE�S�wwwE�l�����j[Ƽ;^�@V`�Ɣ<]�V7ʧ���Ib2�x��G���d	��Huz}��
4X
R���H�1��H�v��?�4���JrZayY��.HY"��
�[T$qfPt1�.��Ór�Ù|����?��`�bF)$��`[�5r���������s��i���\�/
°z7�<IAx�J����p��"���Ϊ�0�8ƹ�=[��U���?�w�.*�.�9��1ĥ&������7�bb?FG��`9,�c�{���樅����)� ���ba$^��\��+�����x��:FGmVFR9�'����Kcv��зЌ�RF3�;���Ɠn�U9/|I��5��}�qi�H���&�ՙ�f8��L
Jb�\��8�b���َMOO����q��?�n�	RA���q�B1DHVjx���3�J�Od�S(E��r�	�)�~a0#��3���>�c�{�һJe6� ��N.7}�J�T����k�z`pp;���<����g&��1r*����������.zn�%5x^�S��
1;";�������)���c%>���"09�@O�T�x#�����<=�ˈ�K��F�[��F�_���+K���W�//ח/�U��|�߾E��S�R��T)��V��P�")j���BZ���LN�>����,,���'8UUU���X-!85��0Z�	���#@��{�_$�H����t�����J;����4����J�!Ä�C��y�Φs�\�h�^��^�����ļ4=��#d���������+T�� 2K_��7�
�{����3�=���A���b�Ԕ2яI�_��V���QA�I^����m�k_�����&N���.����Ѿ���BL旔�$�����q��l�LPg"���*K٫������?��B�r� �z	�\��
˰�p c�����,У	����\�Ǚ���i%�f�����uN���`�ʿ?u� a����������V�G��H�����3�@[n]���r���ߵ�<T����hq@N m�	�CԊE�j4خ���u"�@[L�8)�Y�O&�}�3�8����������L;Rم�;$eo�p�ooono�G�ex�K`�5��~�����u[�2�+�%���ԍr<rIqL���,	+��|��"iAH�||�������QU�����N�ԫW�ƐU�߳ �X7l�������A8��y��&�8��7�eTڽ�~s��W�-;$#C'��!P��ذ»0����q������dj*��h����_��Ȕ��W�2dU��_�2�t��d�)�+�PA���l��� 1���ôL�v���+h�w�m������b�� �X�u�F�k���l�����qڝ%2.�c�S���3��b|QUV�s���t��su._� �s �+<��[.��z��!L	N�*��;Վ #�yx
�fO�>�f�3@<������
�v��G�d�h��`K�n�p"���v�{�N2��ٽ����Rۇ�Q�	)����
99�Ȇ��?]�Й?��:�e:=S�'}�j���p̄^w��t��� 7u���/��s����m��Y�OMCU�23%�u���O�,�o��SE���lb���i!=���NA"�Ma �̵L���$�
��?.ᒵ�N��F�����L.�]4z�J"�Sj��{4������|��V���O��}����iI�Q�P�����e	�G'�KK��_;����a8=?:���Z���7���p��$��|0V�\,t���������#�L�~�v����Jhܾ�����pY>|�������9�Z
Z/�թ|��Q�xď�UU�5��]��5�d�c�$�p���K����@R��Mfr*6�=��4�6I)C(X5���]��J�u��C.Jn�2y���Ȗ�V�� J@��4R������4�I��^<��2��4AQ?|0�F��meudY�A�D�[��P�v�/{,�+ǯ|щ��6���nR�^VM�CL>Չ��dW�2pI���GDb��`M+ש�k$3s-�8mCU��~K@���Z ��~���g�����7$���P��GK������ �2�
��f��-IȔ��BSR4�C�iU�Vvľy0�ER��`�|��WR4BBn��F���X�`=�̳�k��o\$k�jF�������S�SeUB�j8����(�h��b'���t�����M��^!@�& 1$�"�Tdy/���*v�27��e���4�
�K�٪���j�d[6��J��1�ߧ�P�g)(��:�ى@��p!��-Δ�گ���/�G�Ȏ��(K���
�{
s�b�!\���=3@! H�dy�!��l.N3:4d�E_���bh��+�����x�o�I)��/F�x�eӛ�ʱ-��26�2�v�$�!M����1�3Ó�^������V3M梢"���47 �Lh�w�y�>�˥]�|��4t����������������"�~�����@���-����2�w0<�'�$vy��h��� �����4΂ 6�utR�L6��䈄& Ĳ��8��\"�`��]�gvL��"��f��,\���q��M�	�	XhW5�Ym`ODӢ1�h�f���z�T���Zg��}�Z��*�{=�خ��K��P��,q�躺�g�����PJ��r�6$$�u��7^"!.�YX��������0�Yn0���2���7������̭K�N�u�x�m
9:�=44��S�6-��D�Y
m_-�����<�$��/��/ ��>�k<~�T�
H����%z:��	P>Q����].��v���� �=�o��=ݼ>�������h#�$T���2hpύ@br��衩���@�SO	��
	�lL�H>�n����;����ZW�i�SnU8r۝��(8tsw�����<�U���K��t�V��qt����{�a�����#�[��/�{�N����!�j^n�:�eWT�Ľ%�҂�Kč�D݉��t�u���ީ`�4�Kd�J��3�M����'�U�G����>Nr\��6�ǧ�#�f��ׯ�P2d~�����٢1��6/���m�.��q9��Цi8�c��7���>!Ea�4�2���N����2Cyy�����.dGN1���0��T��[�
4'k��l�75��+hN쌌:zz�2_ xH�i�?�^[��]�D��ZH0����	�a�^�]��E�v<Z�R�O닍⇇�J2��vlSx���b��"`�sb��W�_��e��6��y,��h��k�I�} m�	nu8�Q)�p���Ρ<	U�rK}�3i+�o&�\�x�w����Kb� ��� $|��^#�`N�@�-BBC_��C��	~������&/,))prq�����j/�+(a���_�+���)��T��:dus?�ux�hi5�ͧ��%�/�]�͑�9"B�H_)�6�'�J-��vR��_`W���	KʃJ���3-h�Z�3}�udI�Q1�.j(_�4�2�̏����"��KT�CT��kq}�d|VV��* �H333���J��T$�Մs��f�E����Z����v$-�����uM�Yg�_W�Ȟj����O���G	+���BY[�3��B-K1r�k`�EC��`_�n���$��*���:�C�ܫ�8?�큀��d�߿���EWvA�<�hcR�/�"	
@�>w ��}��].bU�)>�R40��$����(4�2�3]8o+~Нڲ�u<���-���:,d��ۗ��!��?����
h�i�M	��\��1%X[!?\�T�H����R��ܰUW�@�tQB�������'�M+)��&�
� k�D5YXXhw<�[g�^j`Q�B�a�$��R(�?���L���[����h���#n�:Y̔Η��}C@A	�)��'�������u_0��C��آ�O���_.F,�G�S��8��U�*�P�ⲋ��)�(ل�[��kL�S��i>|���,# o�N;G%����+	����O/�Z���g@퀻����a=��Qc�B���Z�2\��'`����)��JO���W!r�q� ���9)>^%�n��	_%|��FSH��u��*�v�=A9VsF$\O T)�R���%`ˇ1{X�����[d"�8������$��bC$�w�{-Ώ�s
�Љ��u9�*�X7�~)��#)�m�m�?̔i�B�^� y�#���1 d�
;t�ο�O�[�6]8u�4G��:ꖊJ���P�v}:k/�,�m� y���%~ge��p��Y>*4Iq�m�4�����8�|K%�����`�eC���t���>�T����zUj��-|U�Ό�����҅��]A���v� {SbL�?���i�l�Y�������.��� �߉
��p�[���$�r�tڠo(�d]!��&���L@"�%8
W�3+��v�����$$�d8�/��u���`]�� a[;>&�rV�A%��ї�2�8����g�y�r�!�KN���
��J�Of	��C�����s�N<@H@@@���(o\B�j�����F������55u;�c��ffF*3o�#ᢼ1�%$�~#Q�����ˌd�D�h�$\�Q�h,/�>�>���F�hZBWp���(u�'32��"�㳎�m�
Y��c�����3����BS�$�鴹�ρ�;ܛ,8Z�|����d��E7�AtT�{n'[{����)��!$f�����׬���x�.-��3H��"��n}6���W\�6�ƉA��@���2�66XncZ}����3IIIfxx�^���2���#�؊�n�cDA�	p,ena����0��b�χ��AL��a�Gd �T����AZ��2rN��� -UP�dF��"6ɽR������6���s��u����P���5H$�����j������F�3��g�BT��������h%�C�ȁFi�nmu_+Ӭ����m��}��/����n��zbGe�޷K�/��XTTT��������eV֛1�&v����y�J�h�:�r�����ӿ��01U�¡���3~���D��;a�|<Gd�x�����/���~2@;W"I�x�����W,��� c~W�����>*te�6�ܩ��P�@
I��!�����Z�-�QvJq��*��y	.�f������a�Z�v��^]�dE��-���kll����v�؃�w-��յ1��b������y��G�����=�hX��宂�n�r��������\�A��!�z<� q��yEV��T��H��ߛ�*]�*��ϝ��@�RGp�U���c�I��Z�kSC� �����\7�Y�pF�ee��hȌOM���a�A��u��1��_hh�.Ȍ;;m1,�y����������j�'S`�@,s�����_� -��������b<ڞ� 6�����e�ݳ}��h�<+y�4�^G�4}�jcS�=��pR�`}�
�&8W�1�m��z��%�� ��( ���@�����Y�@���Q�. ��Fv[[[yÃ������?�&Eޔ�ׯsh���Q��:�4�Mø�5�$&�.�Y-�����7xY� D��b6���hY���6�Q�7�&(��ciX@�P��8�+k�����8���<��͹�]�:�+�O���)���l��^G���m�Q���8��ٿhr����T�5�o�l�x�[�߾�Q�iTIh4YfWƔ��rȦ�l�u"B�B�f����@t.�"�������������Z'����8�>R���D ��zz��*:�	5K���g�Rk}7���x���W��$ɹ���jk##
n�%|)���-�1J�Ж�����.>���$JĽFC����k�����,�O���V|4폓�uu��������2(��a�%<ަ�~m����}!� )A���������9�h�ؘ�1��%��s8�;S1�ܨ���A(�y"B�111��FKL������'��@��|E>��0lF�l󒒒n�-�
y�q��������$��$Ͼ_u<W+Өuܛ�K�,fZ$���!�����\5z��B��Si��֒)� 4trvnԓ55�	3P�:��\��f���\?�<L���7	�3J|��\�*�����WGGm����%�o#!�sK��[zC�"""�aa����`8����0$��*(@X����ԋ"���v{�}�++x�Һ�.yx��K��}nRYS�A����X��h��9�N�.xZ����R��oc�9��N0��_$2��
8<����H�Ȕ�CK-��5Iĝ��ϣ466����n,���m�7�?~T[x���dH��H��e�����i����������r��xOϖL�j�����������g-�p�96�B�L^�����cp�ۼ�¥O+tm����\��!=SS��DYg�p$#�I�S:.vF5#��������tR'����B?�c���W�[F�ex�#�2].0�x��x9|��7�K�@_??/oo{k�O﹪U̞:YB||�TMmm;���%"~y�Y�n网�a�<��)��;I��I�K�#����x|2�ͧ�չ�[!Ȧ*�x�Q	}����U/��d j��{�nK�Ҁ��� ����,<Ɩ��W�o�P(��͎e��}��ɸ@�P���}� '���**.�NIM�;�����-	�M���gZN�COB���ݽo4�m���Q���[��G�j�N���x��פ�bP��Ἠ�
[i�q�.�eh�vY	bR�8>�{ �πAZ�YWs���ƱGt��)++�?\��K���KJO�
�?��X�}ߤ�7�-� \�����<�%/�iT[�T�j�p���ھ`���{������ݞS�,���� ��\�{t��B$�
GN��\�@hz��r�T}�\w`)qi*(ؙ��Tu-�]����Ȃ�����@I)� ǠƦ���
��R����F�m��!;o��0Non޳x>?����]9�u��EǾʆ�{xx(�����|�Y���,�ƭL`6����~:��W�XXq�4��]�/�PO"rǋ�'y�8���?���%\�mnl\Fr�����XHKjEa�|�<��'�W^C��b6�9����s@� ��8�vɇw�^(��&���}u۸���uX��%�y� 7R@@@Q��k�P(d�:qɆ���Jo���������H�׉Nŧ(M���:f�w~Ϯ��������B�)P1O(((�^j�������%ޜ�,ܵ�e���@��g�ihq��`I�޽�l�Y]]�%֢7a�L��ٯ߾���t�6$��*%��,�e��:�4�L*�����O��߿�cT� �[��W��R˦U*��əL����p�j�����A�v�t#@�ȉ������O��+�>"���.��4��ɕ��,oo���0�k!�������Z03�1�{���W|X�;�� \�қ�4:�m���at���K�._� K2G���m.W����ޫ?�=������k;;�Tϼ��0Y
񉈉�մ^�rq2���0�ݽXg����\﵈��3�ȑJS�2Y �4�6���8?�����)���r�a��l�_���b硠����(�K�8��6��r�ѐ�	�U����U�d��Rv�	�c�T�)v��e��qppP#���1�`�q������[!�ͽ~��?;F����A߾�&�ø�/B��[�	E�7�M?O�M���,~)�����A�@�`��:�y�o(1=�m	�H���49:6�v�ͽ� ��[ds��DKH�]��
�	�����D�"�AH����?�q%D��E�v�SUf``�1ȡqT�ZA�S~��`�.\)����7���7E�"�BV��� ��E�8n����7�Nk$����is� Sйh��Ť���W-#�d\�<��r{����?G��oD�0O$��p1P{B���m����^OlS�ҡ�wJ�V�Y�Ǌ���Á6 {W�u�l��H^I>�@������xDDO��	#�m�*�����!+J�O�U�� KW��yR��:�O�:Μ�S�w���~�22V�$�ݝ�#`OqX-lU��LKHH�_b���}��t;GX����`��/��-�ߧ�3�*?�����$.��˫�5��b�E@�wN��|N�)ǚb�`l������p�5���\�K��`
.����_���A��?������&bHԴx�>�&`��zs0���I�f@g�b$��k�Q|���o49`nn�9���^��O�u�����!!.�	��/y��X�9����n�B�	9l��PH׹i�hp~���?0P��b��x�#	��p�R�75;{�]j��4t���B����􁒒[�v,����|',��%��w�ӛ7�q���S9l2�;%�b>%)XZ�N �s$���R�~�z�(,L�DC��1��d������cC���,��sm&�{p���0�KK-ǫ�DÈy��߈<eZ�^ y��h�c-#'7K�a����	�QC�J�B,iiOE�b_B�#%%�L��2��M<�#ˊ���4�/�H^Zjj�>�tކ�u�Y�`�榦�P��a3�,4?_#��(��\���QʗFr?�
�f�������#����Pg�pp�A�(,l�9G��M���ȿ��0L��yB�E�o{U��J�6�h�����ayr�n�3�6�>�Ԅho�P��O�w3�˛���9/�UUT�$A�=f�YK��6�h�~@��s�c��5�e;{Cq+����m��_��*��wyn��"e��HR̿V�xW����<����n`ַ��z��ܠ�_��u�^a|����GQ��O0���+��{��F�x�Q:+6;�J��D:C����h����@3�,Ey8itQk�W�^UQ�e�MMb
,Fm]趹�����5kM����YM�L�RNo�G�\�ߎՁ{��͡o|�� ���z�R�v �{�֙�*ejGw *���a$ ����;N��\���S8̠�6�]�$��٧NJr�hNJ)B�t����d���<�Gs9�&�\�/d��x$����
ϲ������'l̀�Xp���h[�E��P�B� �A��,ib���>�q��*�v܃��?���?=;kbh#@�mgA9�1�4����X�=��������d(+�b&�jmn~_&�Sޙ.������� Y`���S.=�M��1����f��K��F���6���K-��_?0�I��H`n9���C�%A�$�^ٻ�E|G�Φ����Rb��Cރ���@6F��=�������[�7O��I���������d�����H9��K�*�1�)���|s��<��*&�GyM�x��/�����Gs�n��C\�����<��SY������*�a��Y-h�ޖ7�C�...�@��]U�i�Ȏ���Lfm����&����������k�f��'�����mmm�n\��MG��ǟC�����m7�G�,ϣ���:�Ka$L�ڋuV���P��J8f�y�L���^N��i�v���Xb��0;���K��a�Q$w�E��nؼυ�^y>����������=6���n^`�p2�O���>>0��\����N��11cΖk@�qY�Hy��@�� J�?@~�c�;6	��A"N0�aBwf+�(:�����rw���
��-pH?G!{c�!�Z�7�9���&�r�O������������o	*�.�:�#�%��>:��[k>���`�M�\�Iٿ#��$ r��ã���������X��vH8:::9�p�o��Ȧ�a�f|+�,�@�����G����Av�Y)(����U�$����j�&��@ti��!�sH+����L�~Q`s
8������ ^�ˆ���r>��~�Ǡ���]�m��Z�J�F��h]5?����|
�y�-���j���������qO��4>�X:��c��/�0��6��n�1�3�qZ���F��:&$^�|h��$t��ǻlK��1����&6� b��DU�f�������W�=9����rD�ڥi����Ke�ʘ_\|OȤ��]H�[Y�}cs��\��y������`������d;��5�j����SV�{�f�W�������Gђ���>m�[��Q�;��y-+��3
۝�!-����(��mfd``G��^���N���HK�jw��=!!a��3��(�R?NVZ�V�,>5�8QrX7=c�C���S��P�/,��Ne�bxo���$
Q��00�T�Գ��s�R�"��Bg�H�A`#\\]��!���o3�ז�KKK9	e�8��L}oa���-�a��W���(� � �P��J�����T ��������v�t��b�����Z6�f�ti�/�`q
�=uq��.'l�ky�����#R��Rr����x8'���:�1��Ǽ�?C���u����[*!�q?ê�D��߼��.�8\kϪ�� [YZ2T�OF�	-79��Y-nG<�:�S�8a��p9Ɵ��ljh8�������?0^?�2��m]x'��:��	e��ƝB�0`ސG �������ML��N��nV_ �= �#yyhF(�E22�W>Yd0!S�tbzV٭��!k����O�(��`N�ׁ�*�s�VC���t�s���M�%����ǧ.|G�ҭ�U��������]��Fԟy�-c��ti�)�?aE
�g$?�fJ�yA��G=�H~<�}ԘG�V��^X�b?]�"5�pxZ����Y��� YYY��H5�������`~{{�K�ׯ�+�r�dL�/��:*����tJ� !������twJwIJ7"�twww#�t���;��{�?X˵ԛ���>3{�Sr��͠*!a:���p)�D+k�b��n32��VK��O����c9!ub�S�{���+����-��wE�C�8���h����yͷo���5�����MK�U�J���|݀�P��q�5���^a<�nL{�Uq�~�ee�O��%��dݚ JlR�ՙ���[@�[�ŉ7�l���qqq��KH�@�JR����EF_hd��s�@O_ԫ��xZ��=�p�u��<2eOg�/(�5�Sf�H�r�j�zN|۩�Yd�(���Ĵ���p�Ҹ@��$NM9���8�k���������E�i9E^�N�%���S��!)Ju��V����r3����$�A��\�M��!��1A�j�R�ż��������D�C[�d���`G��J�r%@�TZ������hs��������hx�����ӳ��Me@C:���/ ������	M�$ߑ�><��?M8OӌP�C�j�o(��~k{���`������m�;v~S$Be�NԵ�)"畚�Z(�}sz�C���l1�N ��A��ķe8&
$�Imli�n0ӗ�-X�p�8
Y�T�t�W����; J�������` ���
B>-Fh�d�߯�.����	��a+��x�����pq�b�E�;�0�1I�yݎ�&���"m��>^ܐf��j3�4/��HKKK�S��Fx����u�����W#�'�)*~Э����,[r�P����9��r0�8@�{z)((��Ƴ�n��U {KpN�u�_U5@���}�,	fAM�͙ uk@��߾��vv�ۉ�[�+"�e��� 1�y�A͍}���_M�ۥ�������ohl$�����e0�B��Jc�$	A ��9�}y�����d����е���><RR\�b,��z�!)�$��R��.ヹ�����
c%z\�(b�h`bD��^n�l��ͰS�G�
���ſ�#��٢�SR������=8�H���
s��,�gG�jΩ��٤�V����	��L!��-i]P�m�����l�t����H��G���ګIxd�h� ���z���P���Xf5mI���)��Ho�yyyF�gӆ��)���JK�r;mXNsN������z��;�ҿK~��%�q�\�}8..�u/��t{@}��n�i��x�z�m�ԗ��mqC�c@	!�$!M<������<�AoV��aUݰ���t�5j�����⥺�c@h]��ò|�#D�A}�7M�V�MQY����C�����YƩ�~�¢"K�h�Khs[���y��8_
��F�oJ4!P���C\2��r����x��M����k$��^�@)��'��0���I����ޓ�̂��ǢUeb���G�:�l��
���zzk~V�o��m��@��;�O��{4�N� ωn7:��l����6����pp&L����R��>����ohh�MBJ������_�gOh#�4
����,�P�1"Rt����P8���!� �윜�$u�J���"w���� z��(}FVS��Kt_ZT�F��k$�6�D�W����|C15�-�b��300h�T�JĨ'���MP�,4�%����*�m��<p�y�R%�%�s|�Ȝ׻�����G���n�W|44�c���`{y˭�SM��` wJ��'�4��J�p�3�[I�A��k0,��-�K�C����NumMMՂ�9����)0׃��L��� ���R�=�.�� (�ʈzBS3�*?�&�fd,s���-�7"*��~;�%�S���z�n"5�B-���}d73�9ڤ��&�Tc O�^�5J4�[2�2�|����aNG�@�I������������p�e$b5��06��驩��{�wD�������8�~�K��T؇f�4Q<؇����lom=w ���,7;�ٷe- �0*:��$�50����u��fAl���Y�	��p0,�YK����T�a1��<][[[]b��
�q#O.��^+?a����;�'і�3�5��g|����N���.��\����`�2t�N��F��q��������0�b	�W�K{�5/vZ�Cc-A4�3HԘ┎dz������V1�tvvC�ٙ�ep�I��C��]xY������eJ�yur��7U����z"����x��X�%njjZa����T�|w�B&Xw��_�$T\����x�131e!#!-�y���8E����Y*
�&Б����w<W?�2uBqW[���N,&sm�H�b��@�cP��IV8�F0Y�~?n	d��F5p7�R�p)�jN�>]���9���)m��g�Gr������{D��Rv����F^��<b�T�щQ���*�$[ZZz��ǧ.�}a�5�+@�!Y�Ne?���j��5����0�ޘ
J}��!���B�ɖ3��p?��ѕ���`�t�&+"V���.��Mm�ʑ�V�������/N�Ř_��s��CI�5���|�B@Pdg�^�
��p@��_���ʫ����8���6���=Z6W.��?o�08��`5�&�u��^�� А9��[�w�U�7Ja��qr~�@E���c+������ �mGȱ�����à��w�?4GFS���C�k �� "2r�0=E�;�d��ûwJ��.� �';��6� R�Qp#���w�����%kߴ��6;��J�Z��XŲ��s�O���1ۏ�":P�hoH���)/���!|��w�I,��y�++��t8Z�x�7��hSS�٠v�W6R%�y]��v��ot��	�n�|�����݋"�c��)����R�pppx��x6Y�]﫡����#����O��A߄�k� 
C�0�]ˈ_��'V�g�t��K�� �������iG���3�����>��}�֛��%Pu�Л7I��7PY�������-A&I7������Y�����J���R����by��&���A EUeDM�o�`�*��Z<.���]��
����ᇕ�6�?���M�	}-�9��IESn�*:���k�p?��9^�U���_��:�ư��n �E�q�V��~��}�����z�M�u9����~LL-��5�bgcSʢ�-�}SA|�7CG{�z�$��q����������[Y� �j3�A��v3z�gz,� o��_�0�43{IE�I�������2̡Į;��K��q� �(b�݁WN��}ݣ*�q$SGf֬0H*(�1*,�8;k;b��7]�[��x�Hz�����?�*��'.|�g��D
�ʼ��O@�+/[���)/$-��ʄ
���qڨ�<R����ȥ��[��=6������)�ޤ��L$���=��6"���-�6 �QT��lF=(E+�G �b����تI��,r�ȼxM����ڧ��z/���z��eLٖo��L�FR��B�j�!	���.2���t�h"�NUuuB��8�����kb^�f��ߍ���{td���͍�����铰W�/_�2�tj�����g*폽S|�R^�_����,�{�# :5yO񮵵5SHP��"Ԯ/,EN�C! ��0�YͷZ�A���%?�ī���ы���1B�xc�RXX8Z�) �i��s�MT��+1KDͮf��~@e)t�l�3�>�os<.��SQR2�tҎ�Ґ�5��\JZ���Yޣ����V����ђ��7M��D ���tN�K`S~fW����%�@ғ/:����������P,��x��r��G9��>��U\�s�3�Y����z*������?C��o�)�č|OP�#4Ņ�9�?�Hg
��B����}8�?eKA3����鴵��tG�B6C��ZFF�~��̻�Y)o�,LL.i99g�%B1'�B`V��*����+Cm�ĺ9���B��ٜ��ʢ�0��Y� GJt��p	�w�~��'i���H������{x��#�n�S�9��̀46�̢�$������0��7��B�0�U�h���)#-m_"󎅊�O	��@Ōep�G�h}#�>�w_[]�.�&w�)C��A���O��C!>5zТͻWlb��	{�< ��5�%���[j{u~������-�M`���R%78z-v�ohAR���u�
>}]�,�al���)e�LL&ۯ�K���ʠ�c|h����<�]b���.l����O����q9u � �V�x �6�6~�|;�n&oҭ0��&񵡴xrg&a�Q+Q�ir޳;�\��p���yu�Ae4C(o�P�1���r��������T����D�}JY�Q��-N��TrF�JK�	C0I=�0�'�p�|�-OpQ8���$�@��B8".�-�8+�aւ�gz#	FC��t�ac��� !��S����,&&Vq{�N��
�ڨN�	�T��_�-���"?/*Ԫl���>팭��ƻ?�)���{%T����B�
|Ndl�9 ��O�j�R;�g��t �fcxq�/� �Z�i��2dm�+�����tdLX��z�ی�MX�4��.�6'�2ꖇf����3�X�wv		�P�揌�H���H<>>�IHH8��(x�o3I����n��9'P�1���yV��謞^D��M,�������8����,z-�ssu���l)Kw���ϳ���k�����=�; ��I:C���������9��l;��ש�����Z�ᡡ������a��c����4^(�}M�"�\�T60�x^ǃ�o�q~~�r{�S�(�\_��k�[c9�C&"�g#UL����# >PW ��{	�� �H�/=?~L����XxPS��|>� U��2�k`y�o7�a�_�K���:v�!:4�����EȾag��|��:�����ri!�꼄�~ojjj_KO��I�2����AAA�`;^ф���㡦�[[{�oiiA�X�'�fF�f$�
�4*5���(6��L�F����Y�����I�k�b��!�ׯ����x��`�2��tl���6V��Z\��#�~OJG�"n�]���>����]�*�Ka�R<#=� ���q\B�p���P�'z����|Ŭ�t�GZv�����GV`&���>h�V@"�b(",ۏJXD�C��U��j,���*��ll*^�9�ss�'�d���y�+����?<<�hw��#���#++[�b��տb4F�CVV�*��ͷ���S@ئfd�܊*'Ly���5S)���2	&]�h�&���Z+��DN7��e`�ݟY��J�Gi	�jz��n�/P�'���D��2z)�dadT8�e�����~��#?ߌv��C�Pa����LD%G͛1�����W�4����D�6R��I[��,V��HE��-�8�&���V `҄���xΨTT[��_t�C%-	11b;��s#�9v獶#�B��N�s,1E�p\�_�IIۉ������)�m�B��ە�?�46ޚs����1���4�q:����;1N��_
7����L9���c)$XHx:�k����E���{��>���Ѫ!����=��ͨ��5H��X�H1�چ�E�>�&�Û��D�n����
[�����5=�`����?|?�ċ��&h�%"%�%�4��}
y&UX"9�.��}���u{��I�˵�g>YY�_��[�����g��]����s�D>)C��t���<���`�}��/u���߾��*�!�����8J� �<j6����-�X�FR��u��p��v�`�����U-�35ot`���ɩ
q����~�����tt��A��E�7x�g��ik�o.�de�2X8:Z��l;5B]U<�tt	��/y��Yt1�hߦ�,V�vW���3���fx#��備���#;G�@����?�ȍ-�B�8�ځ��/b#_e��#��ݸ!��vUw9X�Kcc<D� ^��v�]����qNN���}a �0��t>��t�>C�#��R���S�ao���TjMz��:��������v��f�jړ����{���	YB�j ����`��f��{�G�e}D	��EO��"W��O�o	���^���_K�M�����[�aE�}�T �v@}�Pg���_ky�����Ng2Ԋ��r{��yɐ�ZRc�z��9�%���%~�Z%%���������D��짘]9L8����m��o��{@py�.6�S��1� .�ߦe<l��T��0��L#����tYf�o �)*++���!	Y��<;�K�;c������RȷO�$��a���w�(((eI=_I:ѐ#�'9_~��̒�V/��͈1G�{{����0qZr2�џ�!`�0�jO���S(MI\f#���I�2�)���L�>@�R���g92"�1�g,~���^,�����㣜L`��ܲ��{�D&RR�2��D�t��k܋�N�=??�:=�!�DJ��w�ۉ�:�Q mweb^�x^��b�����^
M@�i����2���`�QQQ���> ��r�0�H��	���~�M/���&�����䝝�4E�m�	�G��D����ry����%�p���ˎ��Q":�yKD�:���!A��Pf���S�j���x���2�o99g��[��<��U�u���Kg�ix�T�(��%��$�66����W�܌�u�-�z��/�?��Vt���?���>tՌ������U<��]���$�"�j�bk2�ll��N	�{�����z��=���=_��釾�a����,�:1!�! �ִ��{���ꪪ�ʙ�WN����*��ɒf�:�̨���|�O�O�vNVrrr"IIH�gArbܛ+[���j�@/5J���gapp��vS"A���E��;�����ُ]&��^���͹}�I���+��Ύ�0����h�i�Iw`?G;w2=���v�������4�`�;�au���~C*��Z�ZI���v0w�kd�+�-�S�P(�ѤõX�T�Dh~'ų�X���QC I=�nNH!���������A-'�{���9����O�>��0o�ES���tI�1���O�G�|�������o�2�;������ �ʞ�{^�^�bP��놊�wg��J�p�I/���*�ps�=�t%�g�s���,k#X�P���`b�50SM��H��"!�Go���@�|��埀j� !�5W��A�\��5��H�()֏U&�����yſ9�}��K��'94�'� Ԭ�o��+����ݥ�24�TAY�U�Hj���4������U���d��̬F�E�x��B��Eo�5���h=����i˵�Ǌ&���H����A["$%m�Y[޺���s!2ѱ�-VSb���Ҭ��"HHi���$��|��3Y!�eU��惜�8Ue���ą��ϟ;�H�+1
i{;��v`�H�&&_xxxb��]�'����z�#���_��p(SI�,uĘ�G�eb���兙���GZ�׬��В��W���5 ��̟��\ϟ��)�|"~24q�b�D2U*�h�b`�ZZ/��Mӣ&&&~`bb�q*ɖj�$���A�W��`�R��]ؑ�80
ɜ=��?��޾ͬ���-���ݛѨ��& ,�N�\D{�����59<�E�~	�w��X` F�״��K��x����Kל������o:�Z�h��3O�������a˱���u|$.���@��
���>e�ЈU������d���xߞ���M��/�~����.���la!u�)��%1__���2����Rc'XֆT��o�z��l+��*�o%$��(=�n������F��y�/.>���|�'G��?4�P�Z��0<^R:��Z[[+����Ӭ�N\\\����.�#��A,3�$�)�{����n�D�N��@����obAS��M�5$�:�/_����V.���%6]�9����Q-��ѯ_��NNN"{�<܈�5��Ƴ�Ȧ����L�M�"lO;��Ćҿ�> �|.�U��?�<�%{�<���~����pr&�k���`�Oo޼�����)z_��9[���\>[^��]mE�����{��3��;++�� ���{���ۧO�/		w�Ns���>k��\]��H��W^)���2>�Ɵ�0�����^ܖ^��jdd$�r��S��tGdZZV�^�ТR�����M3ȁ<n'kB��bn�裮?C����]��T_�����?u�ߗmH�� ���4<�������`I���5Usp� >�A���D�A8 -����h	p�uf���qdu⽰����\����ѯ��0��3b+*��`�^���j�$'�!��߫����LG�O|˄fĬ'Ult�#� %�ؽ�s�h� >�����O��b��6����"O����d�a�,lmI<.�d�o��f��ЫLѮ�>s�#E§��
n�Q#�i=E�^iv+7��[u�,�E{eDJ�ٿ��c�JD+�=���Grz�KZ|�VR�_���QGGǺT�*��\�**b�y��W�m���x�/%�QS_�R�eBZs�y��}Xz�kL�9I����"3��k	�XD��v�M��{3�u����-0Jq`�w�H���M���p�1Y���~�B��yd��贈�8�Y�E1"폤(�Ih�!yht���5��h���*��t	�S�,�5�d���jp��WS�)!��|_���AM�LX��~��������9z~^^�U�Ί���e�_>�"���j���#=��ķ�pҬg057�v;\`�!�I��~�P�z^�a�]&Fi(����}d�.|e88�R!A����2혯��Ô���) ]�9{���b�����f%ם?��q�`2=�on�U-�P��x����:������js�֭_��s�O[r-�{ߐ M���׃�Y�W�]!����}������0�>�}�B�����)����V�M�S�\��衜h��)%�m�u��D�����$�*�8\�]2��E��{�aB�*��nl��c"2+���	��\�YP�"�M����w7-�G����O����סQ����E��!�f����y�M4�@�|n�~�{i��N5���<��]��2ã���ظ����Q�J9��D�ЫprU�K��U���,ii!1���$!�Xip�x�>���;V����U��� %^��Qu/��?��޾V����g���?m�.s0�X������
��}����Ʋ˫+�5��7�+��V}j�E�IPQ^>""�͐��w[[[�P��&�.^|�fB1��icK��NX�2�l?f�T`+��Q�>XG����2���0�F�������ǌ��3�f����H�҂��D�������t������� C�v[oGq�(@� �0��0�j��r	���11�)�m��$�($�@jë˔� ;�E����pmEE���K����݀�_x��c�b�c1� "�"\$\�$̶b��)��-�|y��&����_����U�[�|X�SCN��G�84bO6*Ò��6�4xm"G��1aγIl�鞾�>z��G"#ח28-ߧ����.T�2S�_����q�����LqH۫�C�"���}�T���SE��,�e�[~=�{��םo��S{И�@L�-**����4S_�#�_�4�P$�b�7�������㽇�J�L�y��NH	{��:K�7S
6������T�D
��ܚV~�++ު��-�����m���σO�������qu����J �k]�ਙs��;[�jUw�k��a���֟US{���U833���4��������Z}6�1j���Y����43�,tt���¾k+��L�7�\"�f�܎u���貊
-�
�y�Ŵ-����������<)������6�vȬ6u}/V�6
��4~�o`�!_��aaJ�9�l�55+���F?(]4\�j�*C��/U#r��E4�v{�-�J��f�E�}(���Dǭ����������P�.�/�?XzOd��5���x��np���N�<�4�j��DG��5�4Β�qu7�Eߪ�8m�.G� ��x%x_x��a$�(���f/��g�FuQK�uB����b�JG+�}J~8�R��w�����W�@5;��;/���	������t�P�K���;���> �y�~qe��P@�m�9NU��\��Ȅl�	�t���W���v���P���ʜѭ�_�*ߕ��M����2L�����4߿/���>�@�Y�����Q#��V�'K�d=PV���+�	8�N8��+)(��(��bfM��%;+G KI��@KK+@&�>q=]�L9�K�������}�����@l�|�$����WR�W��ʁe�D�*�Էo4��Z��L�����"�?߸�]�9�w}2��\��R}�$�y����4�(䐞F=�"|ĕK\\��`*!�O�44�M!!}���C�p�({����W��%�}]�/�`b��K~��`i��z13[�HJ2A�𚦦�>uK��ȁ��`��)�����ǡ����z�z��5F	�z0�� Yb�JG+��.L���*6y�F �kV�\�^Wm�� :�I��oK��=ŗj[���A��I� ��嶍���ÕVd^�,744L���v��q����WU��#`�#�,U������/j(]\�s!f����ܓ9^k�'�j�D����T���S	HK���P�}�XM��0�66����$�uif�O��U�B�'���]\\8>'Emc���������b��=GY9�tx�
�6���2���=ډ_�fHKM�|�A����--�) ��~�^H�=��'�A_gX"��j>���i$���ߧ_�K�+p$KU��EE{Y�I�'4X ��ϛ{[z���
	�����G���}/Y�� �<�,b�����M(�)��x��0p�����LLu)II\�!��J�����Wʴ��҂��=ag𚵡�w��\)��/_#T�Nc/�>fqZN�544H��sy�+{ȵ����U�3��L�;�+�j�?�������B!p�G�o&�,`���8Z%###c $���k�G����r|/�����7Na����z����=7��Vh?�̦�{a�dG�,����MCA�)��a�T3hs{���Y�LBU)����Z�RfLeee��� �Md����Ε������mT�R@�e�	{k����Ջ?����I��U@�(���ٳǡ���^�w5�WS�%Δ�_�;���`ccS��z�p:��}�0W�e���O����*��P�)z���K���0z��	<�6m&��ճ��{�q�%�����T���_�a�ţ���a�����D�׵6�v��i#�Q5C�F4?��m000��

b̹qh�n�{;(���/�ͮ/[��VjՆ���'�2aVUU5q�ShK�y@�j	���?��*[W��=t��<�泦�8��w���՟b�E���lnn�Ad�\lS8bmn �KX�MiQ�V�4�k��DK�3���fuh��{:��B�;����65�Ȗ-ߧ��f�_��_jp?��^ޞÛ�.fptwuq�m4%"�����U���q��k���B�e!^����ZD���L&[1���̤��I�r��=���Z	+jj�,���*6��K��#����	����N��^+b��}Aq�!VB8�:7��e�P������8���Kb⓱��=YY�� B8T��,Df�2:999U��4�{piqSS�Tfdh� ������򬐓���50(0P]V�?��45i�����XY�z������uϘcz��I��W1�.TutV��zY+)%#�j�ԻC0DB?�������3N��r�v�
����b���A��ʘhk,S�����=5�����ֹ��< ��۽��4���1�:�]�Ɲi��)T�,,J~�<V���Z2��£��zki��z���~+-�id��b�5 (���ņR%�&0�/ɁFU��2�g$��v����L���O��X5��Z�z�������p�ǞP��3�0����_���@����l�����
;��-��|,�v6�𫋋�ى��½�9���S�����^4�W�h�?u� UK!tL��rC��#�U껮�x�Cs��Z,z�A�o�Z�>�X�eq��`S�R�x,���RBes(�f	���wy7x �&� ����쭥������fO6���L��u@�R $�q�����n2 ��C-�����g��;\���%��2m�p,yƟ�˞��G�
�� �f ʳ[�L�
��5?EY�0!HV��@��|���҉z+6�����***�(z7��]ز`r�����6:#�И7eT/ÖYPPPH
�8^�.+^���e�ڮ�7)��U__�KKK����Z�H]כ\JR
?Q������rCDFֶ��L��}#�))��KQ����=?9���ÇD<��
�@2��	u�5���B��x�����e`�����V�-�TZ�!��G㵼������ã�$�܍n ��7���=�P)w��R�{��h]bb��t0�P�"'~��x�0����|y:�譹�qք���f��*�@�k�1
95$I#���W/_6Z,V��e��%�UW�f�9A�����t��byބ�RJ�ڠ�1ˑ��\LՕ�o�Pq�;�J~�ũ�Y��k	5\4C�zc�ynAa���+<���N�Ҧ|qc_��ʚxl��(�CJ�w�����yQ�^�rC�y~�����4ʦ���}Z^�?>_NiTT^||��M�/I,j��45&���mml��fl�4�}�q�NLJZ����cҪ2��uF�U_^\,�.4ൗ?8���䖀�nO��������� F]�ӧ���`@kF�Of��r@�^�d�e�`&R�B��.l�F%;V\P�vt�njpD����DNw+th+��ތ��Lt��3� ����~��f��K�!�\�߿'TY�{򻌾a����r����KnKK=�qI�<��?'�G}J��+�}�9-&z�uܧ M���GUSS���YS�$�G���
�.빬�f7e*mRgr1��7����7���"�K�ڴ��):B��1�$���k͜��NF/oq�����%��^ ����7�1���:��O;J���yX�Ev�MW�aaa�UFep�P��KO�<#c���1��[=��u�'k��&��I���rU %�ۣ����4��דя%���!��8;_�32��R������贸W^Ν>��Xo��;��Ƭ)�D�������)��-������F罩(�j��H���wO(^���H�~q�2���azIH�u(�y��1� �UϺ����/롫X�ޗ/_��7W����c+���h!��@�g5�S���Yi��MT�C�\���������#G����).����US9� "\����D���o�y��H�KSJ��V1�r��" )���J���켍�6uوKQ�������Gҹh�笪E����kW��=�7��+�tG�U��'�P�5���4rs��p��l,XB���UN����
���o������-?`���Y�%�CW�>^�
"�������$�����}z��s���vuv!�4����<
�%�G�k��In��̴�E�7f�0xu햑P_84������kX	���ْS����it�BB>�Zb����z�k^�D�x��g��>3�+P2��a�RR�qq��2��=Z����1_�#�e �e�y�x�(��C]� Ogr��D���._@#�hhh�>�����T�x��M=2�����	c�Q7,�/�@�|�&��Nye)�G~�3���E��ŋ?#C?��������jsq�KQ�=��Y���"���h�]�E:���vٟ�	x����u�ꧫ�k�8H�y�\@j�ne0{n�|�T�ye���SO���ɾx�%.����o�:GZ3{{�Oɢ��=aF4l�4鹎��}�1UU���H��vw���V���|"�j�X2���A�|%�;63㬠��e=�C�Zۛ����{��+��tq{{� ��[��ぱ�9nvv��_E�X͌���C����d	y��*(d���tzf H|3;	��1d�]�
nT��M����@D��y����%Q�p5�oz�.��{����϶�h��K�	�����w��]�hA�N�"h|�(r��7�/��H%���x܀h��mr��|q��]��f�߁8�QZ��g����Tq����X�WV'�Q��%����������A����
���7�e������Wʕ����S]U�����Mg7��ݻ\\�*�����h$�sq���8߼��
Wͫted��t�٢d-�hh~�ooo���*x�Іd�|,��S�c�-��j��U[�pβRS�(�L���O�����j����L��~raA����(�w�G���S�	 �YXZbѭ��K�̂j*6�&���׭.�e�����m��#��K.U�԰;$��#����>Y6�L�g''4��1Tf�l7�Z X/�U�#c~9X�.�T��ԈH��d��;Q�ft����
����,�P��N���Е�>k\t����Of6Ҷ��D�o��.�+�g
�L�_�I�� ]R8��bFGE�v�r�}�U, ��>V'��E����4�?99		)�;�}1&�N>�� Ch'�7MΙ8Y��<��/,�rzyD�ͬV�q�ˁ:����f/:3�4����Ժ@����J�sx�x�^���C���}Ū���9B�Z .?@>-G�;!䅎�s��a�ip(��0�EA /�ol�p��	_cn��Ŏ���x����ǹ�Y*T�~��$<���P��z2:,=;{_���Zk��Fbbb>�(8�TV&U����p,��aL��9�D55S�@,���{?,��LF��HXO��-{��<-G��~�k��v��r�L�x+"t�o�.w�
M���xzjJ1�I���hTG�(��Jx&�l?��2�0u3�Kutu�D�o�IRFy�����/[��/,Q+QG�.��m ����+�Y��S��j����ee�9ܜ�bїY��^�w}�(�΄�INS�����o�^�݉�o94���f�����ۛ�lƎ�^6�(K�ˆ�Q�f��b5Qc2%�u��2��МIa�ߏ�_�vAJPtC�u� "�o�o�Ѹ�jD�`��P��������cjVI�j��RF��Nk������y^U�tb��ǹ�?�g�k\�i�c5�(��H?�%$��`b��UWGƫ�gg�ػ��g��ׯ'/�7����i89g���̾o	�6~���9j;Y�۝���6���(�K��{f�{�()����?��$(f@�Z�QBn:ͮ�0د�ѐ�ŵ����:���z�ǋ�M�CU6+�$��9�
���Z��|}����\r�MG ��@�[jd�=V����2��y5B����t0�z'�3�����!��������F��m�S46�Ŭ�T�4ƅb�mr�{�
��c����JDDDf���%��EJ�`�ɂ�0��<ö��`�6��0+���PcB��<K7���4�:u��E�۟4��5���`�Ǿ��@''�ëĹΞﺲ�&��r��--ꀞ<���r�Ѷs�������]b+#�k��C h󕒊
*>��u`#�f���켔v�+��d�?�z����I����D��cL}��C�U6ߧ��?���q�o#��KC��&M����annա�?��\c���7 B�x-��@�g�d�6��OetI�3�GCNޱ8;�B�}��ņ)%,&ؠ��^��3:Jk�l�sʐu�`x�Wa�z/�=c�T�Ƙ���ZZ��T�v޹��N܁L""����I6���T��E��Kx�ѻWw�bAH�P���rp-�BW^뭝�(�ݙ�c__j�2hM�`6f�#�'�#�)�#i����ʚ�-���9Bn�z��v���H�<��t��-�
-��d�ލ��H � ���<�l��������˅]�?���m��$�||� �/"��Bg������m@6��ȥ����tZehgy���A��U1A'��K5ݥ�1�ذ�8����L5/^� ���	�D�'M٩n���p�1Ύ=@F��f��o:S��cdll^g��hZF�@��\o�㇩��J\D�M������&�v^�r�ƅLR� !�;W0n	�Ǖ���BK+�����a�7gS�6�_y�؝�j�RSS3����.\��z�EzZ��kz�۬`��C�Fp��W�������L� m����s)/$
�����u"�tC��|T�������5-m:t����~;�,ZO�}�Z540*���3EuV�*�1�}�e���ϟ����� ����H܅�M������ �`t1��z�ƓEޏW�LL#��3E�V�2�E��y����� d����mt Jv|?3��|{��I��?:��@����T��N��yfO�/BV2��
�Jl�Z<&s�"�n�¯)�f`��P������No/v��!'�-Ց�Jg?�����t�T�z/�"BH䋦��d�����|Ŧ�,�I|�>n���߿�����B����2������b?+�Ȅ9��neM����W��H��Uy�\O\RT�����?y�����-���w}��)KT	�`�΀���d� �"���ߏ��|q=��T\9�=�4���H�<Y���\
Ț���\E�Ȩ{(�S� VV�O�d��Q��t�����iP$l�G��01Id�v0��E�eIY6�-V����x��퀥Xnu&f^�)>>�H�3�33L����Z����,/��Q������o��l��qd�����4㣦6�e4��!�s�߱��srrHIH(�%�n3݋�FE�����Rr�mR$\a�;�+�f�dl�k �Q��J�f�p��6b�1��K"��׀`Y6�S���(�'��o'+/�pr��|��fϰ�9��!JL@�"�;�)4�o�P�M��/tH�ts�[Iqǥ������ϙ��|�Å���a��(��j��5���7C21�,ϫ�c��[&���)U\��[ys�aqn�~�LMy6٭6�L(��׽�-^�.���ٗ��:P�@�}�P����Y�\�D�����*DD��+�[��wP'_� �P�~�9V��t���o������>��Gm��ϟ?�9�~e��=�ц��*���iy팑��#b|ѽ{�|?~)e�Z�5��Ū���m���x||̒@�,���/��͒�homM� l>jC�MG8�����ó��������R!�0)#,�l��~o�����l�i����wm�j�cȲʴ�TL��$�m��G$d���<�g���;�:)�Kq��������c�B�bgJ4N�.`��.���g���"�%���	eBC#�x�����߻G
��Z::`�)���ՙ`���*4������_{��O������Q��2�NƱ���-�GJ���efdY!D!{D��u}������������9�}]��|^���|��/9�0|��/7\�X_�����ݟ��v@i����y��ԲL���Ĩ�U�$\��%���)�n"�~��oUM����"�\��7qE&�E���,q?��j(�-kr!j" �ڐ#�I ��sg�d���ͣ��]YY��n/���?uo�d�[�C�@�C'�b&���8[�A��(�L��2;+�zȱScc� ��1���}�2:�������doB؊���ӵ�M:y�%#޻�)����G;�v�Vx�)^ipLqW5�a���p���J�φ���&�t��a�wvu��X8�4�E�G��5����?�,��Bv�`N���w]�
�'�9Lc;�8k%hz�����Z׋�(����fSW#�_��;:����5����������U��mRRJ�u~i��꫷q%�I@ְ�}�Zz�M�dbb2����D�ǚ���8�z�j��ӣ�+�Z�"ndTt����BBuE�G��9q��2�ܓx�����+���9`���F8�o�<���ʮ����F���\˙]�i1f�U388�pzv����[#�x��3�`A��0�I`�����o+~��E��8 �fg�9DEE�P�o!d��AX	~��]�߽AȔ��,v�"a�FMh��A�}�Q�O��6m��>!2���o�Q\��4���S �i�x㶠Ovb"/�b��|��A9�tqF�������q�͚��ux��9�����_l�Fl7i�2jР���W��f�=v^C񆻜�7"�����X$�%�9�S9����O����0Y���&�-�,D�:�&ʍ2��F?�!9N�<�.(¾����(��g�0P�H6�3���F��/��]�[i/�q$~-�5z�-'688���Jr3s��0�y�ƨ[�n���ܹc�V��������v�c�vt���.EG���ې�'�]]�]�� �nV^�yk\�?=�l�2��e���A�<�"s���T��d����	�;թ���g+_1�B��sP���O*N{�>���8����8��{)�7�;��\m_\�5�b�3��� ì��w�i[��]�&��ƨ��_og@��i�ĶV:���n^A�nׂ�Ǻۢ����rV���+�f�)ᘔ,��.ئ����B���b�1Ma��]J"�	uz��ll�==�9---������u����332�a}jn%�m��W�r���ےSR����������]֕��a/���<�EuV�H���ζ������F�$��V[t�������9�W3�w_�򐷶�r���0�.�+���rQDHX:���􀃣��Ц{��b��8�^$tt΢nK���"0 �h��*��Fm�g[x����H�m�i��c@�3�v@@����<a�(���	��M�u"�w/c����t�g���nJ?oN���*��3�E��o����3רV��7��Z��s�ZOμ��Y9��o��W���&,,,8 SL:�d�a/u^��]\||>A~~�Nkc6|b4�
�s�uLL*�_&��й�\G�o@���w��BH+z��E��k�@�sFf�#����� AWF�z�NT�~Ї~߆xt���M������ޑ׉sơ�5�h����d�E��X��Q`=�1�D�E��.i�xP�X������'�>��oc|��9�ǏgRd�+�S��v1K@�O�=b5UU��Q������ۿ��`KP`����b�I�<@o=a=	l�Hr�bS�� 4\�P�b0]',<��4V���o��iI�)ڭ���:xi�e|4���8^	�%�_amfVu՟�q��]�0�pl0�a����YJZ��>}��UhW���^8��[{u???�����9R~V��`����w?Ya���o}t�@I���G��w5�x���>�9���}a�l�"� �߰����Lc3�ն�q���'�O�&ʦ$@�^�5�C�w4��q*0#���-U]��♧��'��Ǵ�j���CT���S�r
g$��Ǟ��<�M�z��Iok�m\k(�a���u����A�ƈ�����j�rm$/ޗ�Av)��L�)�!f���R�:X�F�D���O�K���@T�eea��=���2dF���JJ+j��CH�!@�~���G����3__�L�2b��*�1�Hh$����ӛ�so��h����_i���@Ki��t@ �A��#O5A�ɷ/8�8vf��`O-����y.mT�����@-Z �i���#�D�X�ޱ<!+5�G����*zG(���"�('�n����9�OxsHHH��T&���E:�<Yy�%��������a�#-컂8��Bd恹������I���y�=ª�ԧ/g�]�>��Z� ���1L!�PM�V���^,VM�_x�ᢆUM�������4�%%�54��(��t��Ba�ɚ�������ӣ��x�/\$������,(�B���,]�!]J�d�A��D�D?��iMMM��V T1b(SV_��c����ֵ[o߾U���XyE%�G#w�E�#��'.�a���p_߈�IQ>Jz�\���_~g���C��鯥�K����^+�܃B\��$��xTR���0jK��iu�����#�-���D�%İ��������ũ�����'+o_<.����]y)uK�==H����xy���Y|7k�+��\G�����g�m#}�j�#jƀa�S]]��38�/u�9�<�E�
��d-a>����k��X'�̡#r��>&
�3����q�6���H4H�R�$�IV�
�M�E�2! ᥳ}�$����7<�h���ײ;�88P�*�&X�S	����VJ��'�����;�?X����fF5Z���ib-b���B-�b�c�kk�I���"��]�� �<�vy~Bl�kA����n�9 /g3!!�`�4f�d�S�U��[�E��q�y,�'WHJJ��.`"~�D/��ƨ/3p�_:HnE���aar��1hL��&PP��¸y���{�]Y��ٙR|ch���Ш��N����Q}yy��R��aӓ��#z?�}QTr���_����j���{a��W�7Ҥ\�B�K���:�TTv����8>,��bB��������$p����#�y���� �3IiiOG�-{|"1p���G�4NUH�: ���rm�"���w�*U#�Ӕ��邲��e�>���ʻ.�AL$���q�x�<��o�wz�~��KQ�h}������˗C;��J#�`Q��zdq�47:;;���[5�$�xvA��D�*/�-�(˸ͥh�[t�WUU�������]��h��w<�n6%��Y��®���`��9���ft��(���	�EA1������ե%�'�o8[`�t�b���C#�0Y�gf�~m�s���J����m�g�W�)aF���B��BS�@��Bo������$Ȓ�r�ړG��������y���Ys���'?�C)a^ᄳ���Ktc�����W[8]T��a����v{$$$L���D��ӲsB�L��w��$^Z�Nd��ρ�	\t(,�P����x�=#Y���]���eu'b�"��V3�Ȭ,��@L��r|~��T:VD������բ��=
oLb"r�B���W���6}^��%���K�r[^���P{�b+��˾f��q�4��2���333�b���O��0kbd lE��wL/���"к�Q:�;��s���[ ���<JR��0�p�g-58vj�L����
:�uJ�0G!�2lo;9?���(f��KK�^�s�?� ����QQ�8 ����q�v���H��F�K���Z�|�̌���T��P��=�j������QQ�	S���Ղ2h2$����th������O%{�5�U_��{z~BuBҌ�PTU �:h�h��������k@���|���Wp%��3��d�{g��4�����*�jj�P� 5�:N:��/�*�^��� �u��fBc�~����֤�$�7�c�e�z0Cs�ކRg���7�FG��פֿ��%#q(�ȑ�V����L��JV?K��f��
����[����݉�X�����4�?//)9e���dۭz���{��A��ȁӴ�牎���=qt�iC[k��������>�C�ɜ������ʬK�� 6T�����Jb�8�+�[�����ypf��HSpJGF^�;S�r$�a����m ����� ��ɳ(��#��?��J0I5��lx��;
�\�YF�c����ׯ_��O������ Y�m�v�w��<�k^s|�܏��>50H��F���U��C#��B�4>F�t��ؚ��§��WS;�韡-#`���U�qtp��	�y	�r�"�?�x���}S�'���/{-tu� 8��=�vD8;XA�>F�9�RcJUHII���y�1��E~�cו���ȾNo����.۞ӱ�B0�5��r�l�@�F�c�]w����68�8�w�����$����_XX ������x�3�[�z�E��(*�!',��S-�gz�]�
��.�-����+�pdv��c�������d�gg����D�~�N�ۄʣ�11�f���TwUK�52�B��j -Iܾu��`g=]���×B��7�s#?��P�`*|�^����D������?�Mr���.�w��RUU=BM!9���J1V=[U�x2����jO��.����./+<�^�����7�^��2����� �ccG��!gm]��9<�O)�aa���4?�蹔�������~�=��qpx%_6�A��1�	Ǆ~� ih�t�������{#�`������V�D*���M������F�`x���}F ��x�cU-}���r���LE^WU����x�=�u��g&��e{Rn�@����ʻ��v�j�k�A�^&��X�1mk���9uS{h~!�_\E-t�D`G;×C�0|�Z>}��$���N�6�2C+�ԗ�u��A�bZ��g�������mY�'�&�Eaf C�`���r�G<44tp}[bϡ�\/�v۟+M����ov֗�:�C��`���1�}��YY��8D<��?�΍���R�����]$��V�DO��ynN���4���Ȉ�~�]x7B����Ezj�.jz�9ް����R���mr���;�`b*�l��W1��]���%�V�w7�-���@�ʑ&trr򣠠�|��`b��17�59y���t-�����{�K�\u3�j�!+k.aww�ٸ��o�E0�;UvT�e;H�]�|�ųD���|�dF�5�z�i_��TLj�l����������wΎ?� .���@q��	%����f"E���$8�Y/�/؝5��M��758	l���Ӵ�|$�6�� ��)�X�>|�+ՠ�����/馎�N�+W��[�hw��f>��o�\Y\����J���o\LT���r��#��0�/�i,$~k�j��[�@S]8;BFN�;�@M�D���T�3<�vi��1+������iq׳�X��rY��xY��yBBB���p�Rc۱� /�25p����dud{�+]Y7�r��� ˞�pr^��DM��XάDB�s�K���9?��c;�È$,
t���]�M�>�䙇��.�찈P�Ǹ_ǋ������]��az�p�I,%G*�'���7i�0������pxy U�r����~�
Lz�b5y�]-ww`�<�śL�\F�Q����J�[������f.�^���S=Mtln�U�� ��^���0w����t΢y!��d���,��ǃTv��h`���?�;Z���Ц���1@�*�����2��iF7r:9��mN�G�pS=}���ޞ�� ~����Ya�q �;sr���r��!f��w�ظ��5$Ŭ�MN
߽w��'��._���u�N��>�m�����'iq��ʻ�p�����u�c��0 � ko[���1lt+H��U��A��H!�����t� 6�g=Z^^~���l/�s�݁��)?-�:��v͂�!+/_���/�@�1t�.�.t҃�(��������dO�d�����ߢ���]|cq��	`̔�ZZf�
��}^p�*�\�G$a /D_��W	�Ot1����ё�2�=K�~������q���Ҁ�߯�5B�QChԍ��-�	�&:;W ���"a%T�w8q�v�yoI���+���Y"""�?~�khks�4b#$&�G�����3U��y�H	�uk��*����oO���脷-��R����ә��}
��q��7�%CN��+�w �3vt0,���LΦz^ћ�v�]b='ߝ����FjP�ԛ�jנ��$u L#�xRd�L����R� �~M���#цP�`l8!��D+���З�(���tx�uBn���{AV��Lz5S;$c�kbbb����MYN=�
RzTG������>�.�� j���e���ӺYȑ��� �e������ŭ&s�]|��Y�6�Ny2BVފ�v!i����W��UZ*���24��eu(�������N[x|�[��K�Ǫt���8��_7NOO���+[�FL�;��y/ۄ��.vG����F���R�SP��V���J�X�_�SU�1�|�����,��4�Mi��F=dDXb�F���W7 ?< �EO�g���v���>:��*���+8��"���[������e(�"���Z�Up�'m�ڕl4L���P�����������u{���_9�ƈ$�͖��JC���8(��R�a{F�CR˾��&Ov�������$�Ӡ���v�}Z��o�z1 �-iikۀ ;��/���>HG�s�Lׇm��J���c���G�ߣ Q��'���P�"0����K��4�E=&��v��E�.0i[g�����\u���;<p��O���!U55,����ދ@��c�,s[�����Μ�o�y�4y�q�=�F�XTO9�؞���P�n�q*#��̶f>e(�!u=��vyjO�r�kݮa�g��M֨$�s�!�~hV��Ił�_��_��0�Ekp7EFF�!"&&���w4����H���[;C�!���U�З�U=�E�L)��%���\ �����JC��0h����q����ͤ�Y���t`�@�W}��1�q^އ����	w��kO��=�9��ݴ��Fm�C�n �f�T�ܚ���퇵���2��i��lllD���������U�1��<��8�zll��)�j!in�p�u}��Ƅ$�����At [���zز����=SS�ڊ
'�,��R����d�"�O������RV��U���}�|��^-�`h��n��>9=�Z��iG�bk2��U����!��}RSS��o��6�_�e�"�Io���.G���7��E(���o \\k�����z�����#�Pd��Bj��ohHIk���67���t�ֵm�69���--I���G��R����_���=��,��Ļq��/���9��I:?��h%��A�23D1H�Qh4}�I?�Ӑ�'g0
��:�;����*�L����8k�H�B:��4���k�����Q^�����`�R<��nbX-3�Q�Ԏ
��`g��OH K�r�w�޽;~��J���F���|��B%YA��5+O:0@����Ȳ���?�6y$R��e��6����z.'�����OK�[�G�l1�S�@��������lד�C�_?W ����6���;�������R��!���8��ĉ��x;����&IH�IEE5��767�wF�z���4TӇbdd5�]x��~��,��S�Ғ6���v�����KI��%���׿&b�Ea��E|���@�#K")8�{��ރ�.{���<�@� *���n�V�*�FN�h"�+��f���G�A.����b�����6�lp=lkR�=�� ��,�e����2���D3O�����`x�;�囼��X��imj¡�0���vW�L�鐮5/ X«���*vz��ڶ��ۿ���X��kZ����K�Tn�wX�M��"K��`k��=ce-�y�h��fB 2?$0�~��׮��p�����W--��ҟ�����Ȝ%Eyu3���8�Z�h�ӂ�6����n�h"W��a%�<����MЩ��#�Q�J����\ �նA
��^2���xj^��ǂ��WPRz�}uy��n߮��;�X�~��b��l��S]]]��?+Ӆ�M�D���i�Xm�|���ł�2�������|Sa�n���o��\ߎ�X�� /���P� �s�����_]U5��`M3���<�a��&��{�@�C+��%cj=�����n����K��"̻�6�^��_1������! PL�ڔ�h�(bǵ��>_γ�|*߽�k���-oB�=�vO���aߢ����ְ���"�{�#x��ٳ�H��7n�ֶif�V�[X|�7>��p�Ϛڰէ��v��|r˝����:�$QK(/C@H�5u� ݓblU_*�&���;X��i�N�o�%��.�~��6u���*�|�m�~�{z0���T��Jw��Q|�=�̱8�Fϫ�ZZZ�uuu� Q�**.~�ત�A�UޓS{a>/���/z{~��=-^�Q@�%���n;�Of���`J�Jban��D���>)�ڌX�1��3z���:��Kn9��znE��k;55%@br� _��s[�^�1��
�
ܯ�2��F|A����j�]A����ƈ���uu������->+��8��q-_+��E�%�u��VM��i������ꑋ�Jޏ���	QxC�]D�8�KV�Á[y�qW�V�w��%rt�dy�a��a����f���|�+���&�8ޱN�"Hayf��F*�d�����J}TdduTLL';��l�PoFj�R��,�sWuR�`��� �����C#�w��]�#�Aw���b��p���Ʒ?�&��I�_��5�����=�9j;����֭~q�&.J��i�����]c�5>~t�\�r-��$3E���D�Kx~���q&�/��"IY��|�2�${�B�ޘ���ԟ2����t�ይ>8�����a��?g�;-]�@���,T�ŁN �)�r���-)�k�zFŅ(��4	j�}Kk5��A��?�@���0�\�ˢ�I,�5DЖ�� A�����[�9?���S�l_�߶����O+�� ��.`���z��><І��������Smpve�����w� ���|iLB:�݅�8X���^3��Pe���2���*dr,$V\%�������?S���b���	�֓A�@n/���;/�������bMMM'!���G���'��-3���r�W��؞�'J���� gщy�76�-��^C.�ޥ�R#Z�N�	��#l��[�%�<G�����}n�T �]D'BR����9�kiHe�8��r�#ZȐr����D����=繖���De/k�� g�zH��B��y��i��^3=244,��0�1[�N��x��p �8������,�M�@ ��������#X�����y�&�;"�}�X�Ϗ]{�)y�@�l��t$Y���d�쁭�a
�Vl������i�kr�*�
�:u��������c�t��Yp$��ٶILb�V�����"�P/� �J�0ip��(�D޷�
(�޻54J��/0��f�R�?PZ����2~_+�,z-���\��8����j%�ⓓ�O�/{�R���N�\�/�H�//-�Bu�UNNN����p]]	3vMo��۰h�\�Z���-����R�lpn���(��DÉ�R�4/+�vU]� ��W�����YE��v��YK��_x@3�72:{g�$s�V���E��?>���θ��B���������e�@Ōk�F>^�(
e�H�a���Ȉ'�&Mx?#B ��#o�&� ͢W�����X��.QVgaH�e�kLъ�]Ę����7x�AZ�����\Lo��^<�y����'�t`-��o�=��|ҲU��v�
N"������� s���~�>84�GKG������`�����X&���ધf����KKK�j���p^�I\���(1Ǫ�n0qC����LLL|P'��ϟ��D_�\�$Qܕ���ž���o�o���4�X�<�J��)`,��������[z�b?FG�ރ�?o����8�a]�ɓe7ף)D�c-�܃�m�n �`���j/��9����ł��y�xwAz X�������s���
�ӶY�)��2��ո�|6Cޫ���xSvMd�z�ʽT,n��*����X�A8(kwc�TO�h_G_�����A�S ]�F<��M���
7$��Bշ�lG�de���:��WM��q��gڹ��a�I��J�Rj�k���o�����wa��DAI���oCw ((HΟPRR2�$#+JP��d��� .����D�eKj}$*er|S�j���b�F��°���x5��O��*7�}N��\N0Ei�B���u1�}�O./+;�S��H����Lj�n�j��2�@��:!��S�ș���v��Jc�%�~-�o�}�<d4y�E�y��S���Zg>�������eg�+1m����
���ˆ��-e���e���a-`��X*WhT0l">K���Q�Oô�rs띀�S��[_ �����i]�����\�=U��ו��g�� {v[u���o-��3X�l��~
���vF���+�0�c��`l��^�Kw����ʇ0Rs:q��hEe��b����.2� c��o̼�H7+?f���X���G�4�99��*?ʍ�6��6/�u��y-<�B�᪲`�F2���`�|rN�0��(8���QO+�x��Vd]յ��T �������*���zA��z��<�z$��g�=mpj��R��זa	��	�o&n��|�ĺ�l�a#�l�B�G��u?��Hv}�_����>����a��z��K��_^w�]Zܓk��g��"�0��I?��Vl� v��Ԋ_���1l �!��2�{Dg��_��^)�u���`��ґ�Il��G�nMEbccC!�]��K9�V�����Ur��f 0�z��sl���\9s����wQ٫�&Yo�nȈ{?��ct���D�7�>h��޻mt��vڮ����|]z�g�	0P��T�{��D�hH:�u�� � �s=))�����aH�(�->b�k�z>M�^��N1�-	1�ۗ��U1���`��fn�1b�Fy#���=8G�А���Qccc&H0�L�\c}���"��3m-N��PR�����k�9�ߞ�R�>��qe���cR�CwJ=��y��yPn�%c�,�Ŏ�7��-�̷
͹l�;K��b���R�(�L���E�z*�~�	�+^g�^?�)t��L|uJ!�>|���{��rz�Od��6�� ��_��|2������?g �S�W7�r],00p�a-��r������ہ�}N�~a��T҈���<�S������0��k��	�A�۟�J�u�ֺwsK��D�/�dm[-�"�T�9�U�7PW>����8>%����c̻p�Otմ��ɍ@B���M:���o� 4:��ɝ�F�(�<�ʨ{�#���=88X"����աL�E�o�����ۯVF�� ,�vW��=�A0Qop�=U���gm��~��CJ�z�m�r|477����s�̤�ه�#��E롭�]����of4�I�ڐu�ꉏɖi���j�/T����}�8�G��
��
8:��x��:��X�$����v���0'�Os?�f���<`D����N�d��S������������7��CaR�}�yNJY�6cw�ԠT��W�G8�%*������{���A��C웵���-=���ݱ��� 	��;����M��M��_'�$�#*ә�W�lBFu����W�gg�op(�2�ɋ�����d�T{"{�� �?��Z3oG�Ԫy���g�������8A�<����s�c~~^"������Zmε�&���"�.f�.3�l�O&��/[,_�<�Y[[k������b�E�wۛ4��=�j��F�ޖM��w��m�N-[[�z��'�G��?�^U���� b|��s�PHH�GO��5�%$JOwT!��?\�$Emz���44b|��>P����i�a�K"7iJ�؝W���Z�������!��*�F�����vuC�-d�%�����>�B=�M�%r"t�(��h7Q�4}������1���w!A�^>>-�T1M?~����Ew�'�/��MiMy�i���e^2�]����������S��R�b"_H"�haA���QDS��1v�7�r�*�#���;������$��M ��9�K��l
*�Ig�,ɯ�DȈH���o1��
�2�}O]���&���}csg�r��sN�N��nA�
��iee����w��Y�����y��$2d��ӷo���-#u�������S�hտn�;��]*+w��K��8�u&Ն1�3(y���/JG�u J.ojV�]����,��	S;j �FhI�b�^w�P��t&{�A�n
g�A��Iy���prpH8��Y^���Xʱ�����SCϬ�GQs�w���'x%A��Y���+�Ί�%A��A� ���2���I"��y߬h�-�ft ������}y�=aк{6����$7yy��P���75�x��h�XB�F��ga��Q�����A�T�ު�@�� k�@�ݶ��V�Os�Ϭ�_��)���]���N��@~Ƣ��)����I?�00����^�����ĈnM�H�8��	4��Qۯ��n�r>>�?/E��
T677�Qż?|v��zݷ,��_���#��x2m�Reט'�y�N�W�٫���._=�,�0�L���8�sjx�6����n���⪡�N`��K^��+���j����9�����z���_�ױ	�b$����.�>wr�̞<�9�����e����7�!{�z{��{/<])Ըn<���今6,�7�w�O�*f_��_��zF����g9�$������:Q��p $��c���m���� �ͽk��y�|([_��m�IP�ﶨ�Xw��R+<���n�߃��Ҧ���f
�s�F�: ��^^�,�~������̽L�;~����n���}V��ۇ���T�3�^ZZ�~���<��vaUg���I���M-ڸU�FO���{&o���u�De�'�oȢ;����ٿxQ�����ݕ���idm--���}�͒4Ņ����XT����2w*��������d������
�TZٛ���vNu��&>���@
5����Tc��dVm�+��5;9�V?�p7���Y0�v�y�S�˲�� ��&�~�8I�������&���ޠ���u4Z W���]���¥�m�/M�7�G1;3���;D_�N��ll�"���@�H���s������������8��if����1�KQVM�B�,�PK   �cW�����8 �I /   images/7e277f05-db62-4931-8fb6-9134226ee38d.png���7����D�D��D��	�k�{�u�!D�-z�h���3��� �`�2�6��w���'\�~�΃s�s�{���k�=U�GL����(�Ք������H����/���!qQR�SWR����rtqw��*������#|MDN���N�X�M���#*�(j���d��z-r�
�Տ#�,��!@P)�zO���\N������-rI���"����{�ȥw���
���j�St����?����-��KV�� �O�w?�Prd��:��z;y?�f/}�!�4&"�%%i,�%'_5cdx��9`H'(x�&(�.�J���h���c�����Y9>'�d{kꮞ���d$,�x H!';	�ї�}Գ"�`�Q��l�h�h�hF��yyU�=<|<<ueE� �#�S��I�z���uut����C��<����ԋ'�{�@#b��Z�p��Qq����B�s���\�UhW����+1���s�����G\�DE`/k''sB'�Bέp-F;���������?������?�?�DW�{�H����?q�Q���E�������@z�"��iuu~�Ԕqf��!�G�C�f�¨��"G�*ٍ�@  d&
��� ��:V^^���5�c���$d)��4���Ǯ���(�Kuh�ּ��s�1�l����}���l�^GM��X�媄v��� w�u����A��c�W6IB�`l�
����됭����@��!D���C��_�� ʹ w����heeX�16.Kd�`���ް���p�����Y����/\�l���D���oR-�v�����n�UO���*��X�#vܭ�(� \ɥ�b��X_�/�ǃ��ސ����wm�'��
%�� Pc�kD��K�Z8�L�{�xK���TA�Yhy8Eq}qSr�vX�Ⱥ&}y���M<���o�����=����$�V����@08���Jw�a�-g)D�Ep� �J$e{|������к�yբ� /;�M'�@�ATx�$��J�Ww�(���:X��T����+ޑr��xa-R��4t^#s������F�ӆ���>%}�mMkP�p�|w}�ݟ�ӯ�|H���U"�
��iQPa(����sQlvaW�u�� #���U��11�iDêۊy����L�]����ς�w�j���U;���:{�U�nA. ED�@7�쓌���?�NR#]�=�_����-bKB��WD�2���2�-�Sx��ۻ�*Ȯ {�1�k�nHׇ��W�v9
o�f61�聙K��e �bn�nvxX=�æ|Uy\���_�MҭH@ DD�3byx�O�hBT���C#{U�S|����̋����f��ZL������{ҋ�s�DE���������:U�"X����04��M`.i�Z��|�_Sb{A/��i\{8s��QM��:åCJ��T��I���x~�2(��l�E��'E��������ದ:�4U�y���ޱ#����BK���1��1�,{%�?H�k�#;�b���p�	g��x~A�T񢡓Z����ݹȻI� m^�lsa\[�-ιN@ԩx�{Qƀ.>X5��_2sⓟ���MU�6޼���c ���e?�	��z��O�g$����f^�s�C��R~��28E����B�����=��;Lt�G�>��M�l��;�uI`0B�����/�W�~S���$�)���5X>�����!J�%d��]��K��!��ՈV82=`�ז� �\�^UѪl���ۻfw��wtd'�2&�R㐽�1Z��3v��U���
@�n���]p���>�������j�&���F����Ǧ���O�>�������TJD˯�[�6*)�O���'QV֍�27�д�)QR(������݀-��8�s�1s؉Xq�9	�j9 ���#�ww�b�8�	�_l"؞�4.�~��d���Zt�X�����:�&�����Q?�>b�u�bV#`8kl��KR�q���Z|�֒~���f��=������!�3�'-�ӡC)��D<jo�����ǵ�0�������[Ug��7�;|��w��L����c�a�dd�܏E܇{9�9�Y��}B��7fF�z�YY�O�y��Ԟл���U)d`��O=L�:��Y��b���G�L��xN�K�������)������ӹ5�n��V����30�i�����2����J�%�J�Y$�rjq����z����ɳm����9ttt�}��x�i/x��KE֣{aR����3���r���h�*Xު�M��&uE@�V�iD\�HѾ.�܁Qfc}��.��O`)k����n�I-t��p@�pE�xW��)�Y|[X����ѭ,�ꔨk0߷�>$$t8���	�����m:����Ί��IA��?�"��3��h��ٶ�&�^-��k�����AS^�s{�������]�9H{����s��gӅ~�����W��[
�[Z��[I��;�h����#�]�m�Ϗ�Ԙ$v���Cs�T�^��gh��-��͟�R%�$��&	���i3�9�d��_l�:GH��6���Ȁw7���ݯ3���˷ĝ�����+p³�⫿&���S@Ѝ�H����M��$yЏ���v�1�����wM 0X��j��ʁk2�y�t�����D���	����h[�b?W�n�QNPZ�2�c���L�L]�R[8ͦW��Fd�4���6��^t"�xt��[ݘ���~��1�*���7C4�N�e����Vx�n��4{�ܩ���*�Q�(#�Θ� �t�߯k�z7��c:p�v|���u�e�ӛ3����˲^���
Q��AW�e�@~
"��	��Q�Y^����m�ER�Q�S�(������.������[�ыO=���7]H��吊�I�n��y��a6+��J�lٺ;�eZpCfS���X\NR2dg������P�B�Lh��㪫֚���R>}68�����#��~�t�U飘���.��0,VV�%�o��5�X��6ʂ�t���yd:w��s`����v�^r\�`��VQ�ƴJP��;�_`s�X���fyF����ׂ��6���C�Km��:�����۷���}�#����ǒ��G�YM����r^�<�I<&�oþn���4Y▏��r�|�����l~�\��"[Ĥ���.>0F��I�έ��p[�j=|Jl�l���g^��j�"�-+�Tm�Ŷ
�� ������TQr�e�����kH�+�-�[�����=A������H���g%s\q����8���[����\�v����Wx_��C0F���(���_U~QKQz�|S$&f���N����ܥY�5�ǻ����Ԍm���f#7���t�����K�����~�&�
^�]���ZY� /ɀ����
V�h��B:bguj��L�A�>���Ƀ&���_�ߍ�)U=�11���Z��%���)K`����I'g۹�w�]/���V2� ��
,�v3L|�d�G{U�S�p��8�����U9ܹ�9�Q)㌪��D�R�L��@b90�"ڹ�(�GV�y�_x�l�۹k�#(���8�㵃3��W�l�P���MS�^��7�<D����ijsz^o�L,��!����>�L�kh��S�x�0�2ROE���V��l���@�%�%��G~s%q�D����p���1�قD�t�V��(3�ɛ��_�<e����!7e�I�Sq�=�c��K����`)����d�g����҉��g8f+��Y�LqLK��%�))���U��� �"���[=?m���q������e��a씏ceמ��8V���T7�Y����#��?�3>NX�>��l���D�$qg�S���Ͱ�R`xܣ	�Ds����A���-�E�7j=�h,�����U׉*ї�C�]k�	���U88�gtz%ojZ��GY�U>\:2H,2�0�y:�+���H�`�������)Y����Ta��3af��	��%��������kau�<u7��K��R�`�,��94�8��xD�p�\6�-�۠��2�l����f��p���n�B��šE����e��Ĳ���&D�p��w�Ȫ&#A���t�p���p( :t�x�M���������¨�t�g1!H��f ��v4&�0��:pE����:Gi��[i��2��Kխ+T%o�6��ʒwm��t�~m~;*�ټy3�QY;���O��Ή%ڤDl-S�|BT#��c�SV=�&Ͻ��H D��������Q	�B{�+k�Kă����M�G��SP4�Y��+�U���Y�dj���hRR��� ����՝0}�����P�
m�����eP���DC~k�WPv�|��Hϓ��]G�/�@�%�ȯj��q��?�EO�,nv�j��K���㮈��#w-r�o����q=,�P����������Tf��eI�-
����;R��6�F�ƙ�޶�,�����\`�����	�s#��%F>��j���
�ඞdٻ�e�w�m������5q�{T!�" �X�����s�v�*tc��6b�m<{0���/����1X�y�_f|�7�Z���:�&S���*g$���_<rCe���n]PQV���VfT����'7ݫO�{mݭ^�g˪�y� CEіӣ�-�J�WU�)��� �ŎQ�Vw���c�q��c��F���#,̝Gs���F��#���tQ�P��GW1��"�`��9(�3Yq���2n���u	���]�� .zto8JΝ������O������=J������^ƒ�ÏW�7l�F�٫jT�H1U�[������Zu建��~T���V �݋H	�WbX�B�شa=^R�˙{βj�y�KE�]�pi�����{XC�S�V_T1n.���#~o�$հ؅D"��q��u�$)I�).NVM��fV�Ds���r%6��q�✧i|��Dkgn�Ov�%�r����zx������$�O�<<2��q7��`1������:剹C��J�LC�b�b2��]���:�1	��"���7���u����ɐ��Z�9���
=W➖dvK����0��x�Xrr�p�c����Sǲ�qYYH�7��p�
����5�n��3:m�Uh"�S�T��h��C�M3I7�9r��,�`�Z�UNEҹH�1�]��������K�_UPB5՚w��n||�Vڷ���e�?u�hXᆮE������P:�Ϗ�%���d۾%��
��,u4��$_W)0�O`�u}�G��p}��$��s��Q��T���x�X8�/Ç囖&��?�����׭�N�4Yb4�K�q	�N�"M(=&�����E���ݶ������WT�����E���؊��A�I����L	nB-�)�~����Fx���Z)0m���R�؊i��K�zc-�6�>�~f@�5zHՅ���Te��0�ٸr<���^��^Qq>
�N=��h�զ�ǉ�p)!��z�(@NI~��Q���Ru��t�Z۬l��}&:�P�a�7<d+�t� �Q�E��Z�A��SX�un[j��6B?�"�'"��s��:sw�������0�w��I)����������,�	�wD7U�||!\��I�'}%���g{0���}-(��MDH������������t��I�$�e�á A `_׭�,��=������UT䠑��͙m��+6r� #��*�0�t(�=|�.`���$�:< �>n�3*r]�.�?
˓���u=�@<�1�bd�ʿ���D�L:��6�́�*��d;�<h{�=��]~w?���]��l�w��34���X2���(���f��W{�@&CY-p���b�`A���*��_񚬟�_�>��g�VG�	ӓk-�i��c���eG�ꠙ�9�!��2���N�
yR�z����?'��>�̹_��po���נ��]]�㼭Ǎ��8�
�H�9��� �8 ?�uL��`�>�,��,VQyMt�a�����kx�i��ql������*����@��̄���a�x����݈����C �M����.$4��K#[,���|������U�(���2�}��r`�F��(Μ�n�3��y�\7Wo��5��mv-w�)!�Qk�R�5�G�ݚ�����@59�+�r�������=��C�LN߇C%xjʅ�8�)�?�M�Gǲ�G$���Q���:��,�*+�q�I��iC��[;?�z.�K�?\"������d��n{�o���m��q��8ŠW�0$��P�����Z�*|M-SW�����9�?D�/$��V>g�G��9���J��0/}���,�9��ϠS����b��Z�mH��}2��Cz�Y��?�G��U^p���e��3�[���=36<7��?���K���c0/�F�5-�V�$��ԙ�r�(7��;"��;�G��N�s�`�2<v�A�o�޶fWm����Ѿ>�#��qsj]�������ě��׏��[SL͹2)~�nEGg�7��s��
\��0)z�S�R;j!��A<Y��!��4�X���B";�n���](x�m<9�/<J�>J]�����.,"���&�Zm��/�%2���EG�K�W�$���9!�"4ز��
vѷ�Ȥ��|%$�����n��)藧�vM��<�#t�Q[.��V�]M��˳J��>5��O[0�~_�*��o���M�=�m���/��n���h���\�J:��~P��PԟtS��B=](�$.��+<~.�>>0��Ì���r
ڃg[�L��34�:��У��e����4|�]�!���~��Nxd�%���L�G-O�O
x�=Wgɥ�M��s���a?+ʈ���ĺv�&�!{A�=�,-�+煮B���	���Ŷݯ�_wc'+�o��R�~�fݒA�$���� �����/z���d�[ЃXh��0BL	m��H�hk��|��w�];23Cn�@�P��o"�:)�:!��,��`���V8<��P�'?;�y��<88�d_
�%��W�o��[M!.�qS�Ǣ0J�����to��4�	�2I8��<)kY���+B
�%6�3fk�w�WO.�_��p��߯�;c�_Xל�r����ʪ3������Z�çw�`超>";��6j�ʵ34�F�si"0��nAA�+���v���ʜh���\��>����Ϥ4����^�\�~K��y��``��p�������PƋ���btt����l�E��r�,嗝 ��i{/���R�ԃ��O
Mp�I��5�y޳'�#T)�"g�n�uv�5�)��a��C�?7�Ƌm�y̄�'�T`E ��H���w GlX��슩f[}�桦�4�dڷ"����&ߙ�E�C���DB�ښ�+A�_��V��AD�VR�� x���Q�Fs?����$��*:�
��z��s�Z{�E��Xu4���� <u�&W5�!�g�GӴdd~�nۇTlK����}ź�,�.gҙloyV�lr:��Y�Q�h�ά�ö�x�G7x{ ^V���9�����#'(�ތ����J*a��\��C�>)"����X}��h�b~:��������*�Ֆ�	pfh}�`��Ώ�ˠ�1X��v�A�n��*���N�a����>����[%睽��4�*Q�;��y����=�1��yDس
�$0񩛠��VEIzI$,���$���C�MIVv���G��Sw����&/���Fܕ��/��'��3�͗$k�Qȱ7���aO����s´��P��t_��K��fu���E5k��-�sKu��dX��t���)���f|_��V��$��ۣ˱�og�uՊÌ��V�{�k7G�va��E�w����篘!ѐo%�)��0�8������x���m\�%�)�b2]�{�%t���������{�������l��ߍ��6N������Ko���������\����v0���K�;��2�<���ߜf@-�2����u)�XT��{�*�}��k1���b���#��73<l��i�t�{B�Ɗ��B_�HJɀ����NE:vs�Cr>S��bYS�_1��2����Rƛ$w�2VL�2��G����>�к��.:�s1�����x9k���%�#�S�Y�� ���GG�s�dQ��ȣPT�:%�LYL{oɎI��U��1�yTZ�@�Atc3�G�-��9E�Zw����Kd�wkJ���UY��4F�O]sK�ר�ef���ο�-���-�%p�RY�얮��Mu��\�\lJ��p����P�bhFh����cK-d׌�6������+=�e*ߑ꿣��֚_�����v 4&�����|�5�{��'P�7���E�@@k��d����߳F�	/aӋ�Z�%�a�,�<��_rF���;��������
v:��.��f<l!#T�N�(�M�T�Z��f�q 
���e쳠�c��h8q��p;����"�����s��`�*R�'_�s���?JP�x���d������[\
@�$�����4E=�M- ��9������kU�]�M�V��
��v�@��Gu#^�b����]���|
��>}��af?���
��g��"^=֨:|4�kY[@]@ǭ����<ld��HPz�ό��zh�b����+�[;�?� M��gm�`񇸸)�S���DL]z��f�����x��x��U#��R����R�j?�2�3�8����h��4��Hn���<����^��Ͳ�P�p3�.�޴�X���3kA&��FdD����2�P3_T���R�E�<����/q��<��O�n|�%cwc�DQ)4�`�O��i'Q�ҦTX6���^\�3�;
&�B��47Gy�n��^3A�	��*��)��ݦ�o�x���&g���.��3���y��}^��R�33�0���aŔ��7�ݶ������r8�R5�jױD�6��X���je�W�y+�2��b(+l,��~/�!��!�&�)����oB`��[�g��Ȁv�M"U |�%����șX�$���~�}������6��lB�b{��Ŗ��Z~�0���}��ު��U��	Ct�w�z$ c��e'���*��B�n{R�z�R�]���I]-�"�j�7�S�#�BNt��H_`>�A6�8yR���8���t��;9X9h��+�|�q�/�4u�M��~��mf�ȣtF���k>�>�,�LeM���_���灶%/�� �����(O�
�tqS��5�R��$�>��n�c4<��N�����O���G�Ց��e�-�Ԣ7���E��������F��7hvu�o*L���(9ϖ�\F����{�e[Ϝ
�N�C�{{j�T���-)1_)�ٲ�j���n�߽[��G�@h���(���,�t�Z��������������ce��q��8�	�S�z�**k� @��Eg�"��-��/澝nRw:�-$zr$s3��ӓ���ύ�.Pz��Z��爫�R��o��l;�R@ݿ��:[
�d=�z *��`Rm02m��	Z%w�����T�paw��m�h}Gر>7����ۋ8�h�/N���J��"�g?ُW�x�_oQ�ݨ���@�o=����~V��l���6��QB�nZZ�ku���ab Z�^{�t_@�*��Cy�>ޏ�k��Y:�+g����M��f��,ox�h��c�?��	�O�����|B����II��q������OH�ꑲ�_����ǹY)�F��CD����aGt闅� ��*3c�������o�-�DA�>���.c-�$VD��Ry���
��[ټY.��Z�^�Ye������{�b��B*V6�*K-?:���C�먟sq�>���̺v�l�ev5��M��g��裃wT;�GH�(�5/���TV߀2~�A��J%/��Um�(!h����XY^
�n'ܦ8V�D�t�N��4V���e����O���_RF���G�_aj%g�	#�fs�V�pψ���_MV}�F�3��?Z.��g�4�?|5j�,Ș�Q���'�;*Ry�[1v������v;�}L�f�[3�B�K%�GSt�~X�K+1��6N��:#J�KT�������(sUF�3���F��� ��y�qO<}D#-bF�Υg$/�³K��9�v�#;Y�����?èF3�u�~'�r;ו;}N9��� P ����T9��{�*�yF�[�2�9��+Hw��k�V8�p��QXd�m�^sIv
�4�����_�|f橅!W�-�;1�@�X4����Ʒ�"���"��<�]"T��/�ßM�T�}�"*���:Tώ���.S#m� �zt��e,S���*��vX>wL��{�iכ�f"Gh��V�PCEGl����3#�Q��[��^��~T��c�6�x��i�֩z����PYy��D��3���A%�(J���?�V�˖% �a�}S롁;jX�M��;e0N#�L��`gKQ�@�����!#�W�:�і�Nl�[~�8�M��x���ϝ4	8�{�:]��rsڿW�v�R�.�,s- ��5�%�&
�ssZW�u�
w�_-f�� _J����'-̠��T���A�o@��'O���kS6E�%�ȗ�2�=6Ui�kW$:��% ����L�o
,A|^]��,������C2-�<�T�k��dV{Yd��Ɣ��u�go�&Ӓׇ�_���4��`��.�LJ���i~�*n�[�����t� @�Re���?��wݸ*��i�T-��ws"9�9]h?Y�L��-��C7�	/:��[�����sw:WO��u�vt����p��T�ѻ`��g0y�����b�Ƚ���ȩ�dU(�{vX��h�#���(z$��0ןe�9�Ӵ^�t�D�����}}�<�֚=(��/���I�����Ȇ*��	�&ٻ�F�:O�o��\��Yq��Mܨ��>0-��:�N�a�9t���%{9�U�0�W��O�bsV?YU��Y�j��HA�"��}檂�^��4�
q��QBF�m��&	�͕,�Q�.�#`�����J���2�O�̧~�-��ȁ��T=��5���W$�D�ب��A�`~7�8���5�\gd�X��%�����<(��=*a��y�P�
+�)c19�c��J�WN'	1	A�fj��[E���u�Qn�>w�;fS��n�$��Q�坧�'=��z��ք/`������%[~��}�:q)�r�D��Z��6�N�XR��tPw�G���3:�m��d.h.��g��
���2��!OR(cf�uw�*��\���c��1��d:)�Z�a� ���W<1_��9f�*(��q�J�<���/�/�W��$�$��yZ���ο1e'���Z��6;%�2#q:���:�n�ɂ\�`p	Cn7������,����ãl�JO�2��=���łF�m�{D�T?^Q=�*�Z���!Y����rD�w;0J�<��<G��pYaR#�{qq7�G�7��~�o�w6p��5mËb�q�1�0��a+�zI�Yv������LGE���P�{ySԳ~����j��Y���j�K�f���-��=��U�(Dt(�^ߞb������i0���uk���ڴƩC�v���H�Mᅗ'4}?�x�u9V�;W.ʟ���`��Ӈ����"�a���K���8��X��v!���Z�eۿ]b��^?�"�	 ��B�^�̅�Ҧ�ž뚈3uq�}Yj ��J �!�Ȏ�Eg f�.�w���<H߰2��	���P�h����YJ=qx]ӂ��m�ڂv�4��+ڪTIU	6`����&[�T���u�ؕt1n�ě{f����5�No����Fc������A�i�ݧ �'��j��^�9���9I�+ƝR}v�4Bb/%@�^�!���f�KK� ����Ft�c��"y������D�>}���Z"�����Fv�V���JO��F��������44����W�F=���	��-�X g�e�<�$E�o�7��y�m�<Ga5��!�vz���wL C1XM����n�Fc�o�KZxѣ[�y6k�-P31g��r�}d�ek��r�#�5X�i$)���EuTW��nMZ���$�}�L�{��W��DD~�PP���r�!7���/*����L���0�!���M7�%ѥ���O�.콢��a,��ѬǛ���b��%����N�kx�5y����1n2��Z�w�>��İ?�b�C�8���i��,Xٖ�=������O	�H�*q5U�z�萌�-!��\��or2d���t+5��s��\H�.&R���ӆ����,&���M����l���NK������t;G�w���V�C������Wv�"#{_C��ֆ�f�G��n��X�陔�l8�����]��8�0�axE�,/ǁ�V��X��n�6�Zʨ��8F��\ �nW��������Wę�Bn�2$�r^$�e����j,ؒP\q%u[�#�q���*<&-������W��VVf�Ul�#.�m���"k���yR�Ѓ�݁@P��Z����#�}J7%�a"'�O-���[�X�a"5����}�F֑��c����1g�o� Β���N�Kըl�]]%�'�"���A�H��sr\!�f4Q�u �	���;�K�18�ݖs�����V7qΧ>�K#�r� � ���0���ag��y�cʖ��[��Ul��\Q�iP{��L�#x�xMv�= �e�F̘�R���O������ve#��mJ�.p3GMR�q�<4d�(��C�͂�<�Z������ t��<z�����������~��O�r����?����i�C�m'���j0}��A0��d�Ǚ8>��A$�Zͱ�@屰��4��n-F>�ޖ��%�(��2K �O����8�w\�MZ{��T�8��D�(�1�������6}$ ���=S�������Ji�+���8Լ)"LWv��U��l�"%��Sf,e�{me>�3�h�����M9Q�X�ȭ4�G�?�5l{���������S��_c��ԇ��H��|
zBl�Rc�x�q�Y���P��mE���1՜��*�4>;���4���iM|�MCIlz��D!Rz4��Fh/�/�����f�mʭ�/x�!�ȏ�w��zCt������E��]�̫��˞7��n?�A������V`Q����9Y���0�T���6H�}��K�=��8�6�����J��L�m��|z9�9Cj���{V�͓W��������\�z�X�tt�.�z_����
�R���k^̰�X��3$K^6�X�C���*ο�t��ʿ�*�:3��35_=p�Q�L H�ŗ�X�ҷE�ח����7&g�A"��A�-IΪ3�eB(��'�-����+�\0����� s��"���Z�ͣ�N7���s�Ǌ5]��(<�{��_���{欁��P0�O������J��^G6Ǚ?�ƥ��T���K����o�������I���W.�"!��P	b�2��zr�-I�f���8_�s�d��K���a�"�`�G�vM��͔�J� ��r:6M��*����̪�S9zuf�7;0�W�B�񹏭�žvD�ؒԄ�%ߛh��A(�R��=�-t�3[¥[1ڸ�����vb;ʌ|]:9-��K�n���"�1��[��� ?ѺDQ��h���\7%�����DČ*{��>�x6�3;��*�!6Bu�[ufZ�d�w��߮��7�m5��T��m����T������pܨ�5O��?K!�B�y�b 葽����x���4��@�V(����.LoK8Yl�p�Ö>	ƿ^/d�n�e�z�lD��b��=9��"���u ��74�Oa(F~}�66����nL��9D�� Y�4��g�}h$�����@��-+�e�x�P.���!��^��^�x��������=�A�U��{yX��ja5Y�w"�f+[�E�bu�}:�b��V��/%VY��\����^΂�;giq���ҕ\hΑͦPv����g������GG��?3čH��r�*��MS�٫����@�5��_n)RF?5H�t���t@$��5l��v���o�`'���]�yJ�C�19[�/-�;^�M�x`�C�l2Lwf�R+��eA$�͛�`Z�g��/|@}�����C���a���f�"�y3
�Tna�g�y�����؊���'��:6vվth�y����wH��ۗp�����dj^�m�XJ��BB�rF�:m�S���#�F{0}���q���<�a �/Gϐ�&��dA<�xA�����&�8�D�t�+���5�����ՙ�B�ON��'@s���v�O~��g�xEx�����]��w_�P{Gϑ9#W�i��w��؏�I}ø�I�%q&9��FL��𰝲��E�n�/�g�аPU\>n���6����[���W9��&��#6�����7����r�;�����e۬�}�@���\H��+�k�puW��4�!����i��ߗ���R+)Qf\<����,��Pa|�����@{՟c��k�t�oۈ��v���4b���G�ɣ�:S�L����V�����
���+���r^m*��&7r�zCc�	s?C[[0�a9��$��P��vE�l�6��]���k܄M�j7Ý���e��iKͺ�?R�B��̒�����j^�`�a�Q!���t`�����e��[����l�9�|�����KO����D|�r�><Oe*�j�4ry��B�h���������wm������m�Gͼ1a-���E-ñ0�������]ˎȴ�(�>Z��Z�5��]m�u���}��]��qh��|�k�?&]��g����(��孓��p�C�Mn�.�?���TYWq��&�r��g�
I[�r]~�G���ɽǷ��=u
�!F�0k5äL��#��<��*.Gq�"�2�1l��V�O �<sZs�*a��0����'�(+��Z��/�#6����7~Te��Y�#�N��S%�^ra���Q�N�i�nBL; �j��U~�)��ث�n2Ҵ�e�]����I�=��$2�|M�W�90n��xD�p�C�J4�L����"%h/���"�?p�u1�{����J�;��(���<e��ϒ�b�m(���S�7�XЪm�^��ur`<(���(T~T�֘vDp�I7��.A�hx�˖�p��X��ۢ�,�T3�Կ�������3����v�9��8��^�y��t��%r��/!���t�{]<;h�]j�Q�jo ��t�R�z�4��xlh�1_��36����ԗ�>���8��ATv=c�
呿P?ۊ�&���Z|M�S�9:KcY�o��|�!�ĿRņz��+s���d����Z���g�?M��7�@���b9���]��$�䑌�)���x�{��%>�$j[�f�Ϝt�7���X+W�O�m3�x"Q���9u�p�|�$<�������-a�'���D��~r��on�4.tʫi���JOBZ����-]�N�� �&D��^�9`)[�� HB�~����%7��n��V!*U@�������l�"yz�~?��*���}mE�
�̺a��8��f[ha�q�6�$Oi�d��A&��`�w,�v����.^�d���w�Л�o��"�n�dҼ�nf6�K�#R�pS�����r����S*�"�@�Հ�4�3���� `�7��$$���)@�|hl��J�:��uGa;����-���z6�n���{���;��	�g�*�'�c�b���	T��Z�S&�:�?d%Tlj�'�'�?�	���.n?��e7��H��HWLĳ%��6#��#�-i��#dʆ��|����Ky3���q�(!�,wb���["ۋn��ٗN=f8A�G��Ǉ����<��յ��?��;mf/�,ī��f�yD;J.NV�3P�Up���)�Z+	h��kE�x�K%-DЗ��.��ڥ|b�����Bc�4�Ҏ��:uiY=����n�\��tZ$�ʽ�4s<��k"8;r�&ة�k1��gX�KD�{�d�#�@b�hG싴�GiE3�C��b<�e��{��vbŃ3 ����6v�eU!�w��T��,�Q�J��_Dɋg�QJ�A�i%��n��Y����C�G�Ԏ 'Zb�7��_���Zl׍
�Gɦ`��oa("������v9�6?˔!���é�$#w�39!�#kǾݪ:a�)�B���{����(,�u�L�[aQ2�����+�҉=��|,�K�-r��@�򡼢�T�J��Ik��z�����խ�O�K���L���	��#F[J�yP!_u)�s���t��d북X����B�n_��%�����QG_㾺s�d�����x��^46�k�+o=��N������>^�,�5��.�s�wk�>��;Ъm����ܮo�w����a�m���܆���t��S�Կ�l4j��D�� �3��Z\Bw�q/� �q�j|
�J"KV��_�$��H)ND�sXkrc�r},��e$#�I���d�|����t��_�H���6F�~�ʆG���:��Ag̯J4��w{�갂R@X;��x�3k��Do�0�a�$rrwf���TG�$���pU�F:H�#.9�P�!c�o��C55�ź�A�=
yj�2R���	�á�lȒ�,
	��
���.�=N��&�a<r8�ƾ�-�D.E{�S��#���"gL����3{%���7���sYY~���U�ׁ�1q�!����־�H� �*�8��׼�3�@��f������1��N�Ző��a�J�s&����Aj?��nr��v;���dpV�������������?�2�i=d�/W�M��H����04ѓu�B։#_��9m��;Hl�6��=��;WΥ�6����CQ��Ork��ŵ�8>hk]\��t�� �"|�3������k��HL=��`,߫����@�=�&�!�*�������ԤA:s��@?<p�ZZ��b���V�Ps���8��k0�WY4���DqXca�Z)#�8e/}��~X�P,.�%ޤ5�:�Zdy?���iY Q<�#i��� �Hb��5_(�F.��Y��pJL�Q蕴�F%׋��۝��r){�NK[Y]B�g>���n[�:#���#���i��U�bOP?����6�0�ylQ:'��_���u��<�پ�IP������D� j��y#����A2#�!/+k+���v�}�^������F�H�ݥ���Y�Y����`q� ��h�a�R�G��ym��m�F;����ae����׬5Z��4֘Av=�i��j`p�ϰ�v�������>����r�¿�h��b���'e0�F��Ӟ�	�F{����![KD^���&��"T�)FD#8{�� ��]�Z΅���A1RU(�l+*�"O��/��C�p�-���I;���y�bwm��<!!���P�qX3�;�Z�+rOP�Fk�M��R$51�4��KSB;(k!���u���jzȲ#�hS�'�/�Lr�m����o��D���m:�PT�~� �{��d���'�*��b,�-��X׀d7������FMׁ�5��Q��:��IY��ނ�5	���} �LK�{���;�%�U3��RWd�}׿���{spO�K�����;�	�o�]��q�7{1���1��w�fSvI�^Ľw��Sn�_���i��3d��5e���âs�i��Ak�|�{H��'�p]3>�����B�6��p�zz��L��+d�S��V���`@�[�v�8��0��3�5�h�t#ǏN���0�c#=��#�*>׈�C`}�ѓ�2a��A��j���2{me1�ߺ��o�F�!�i�=<���D�:�q�bh�t|,���2-u�Ř�1����DH�k��"���<�G���*�H	�T.� �9�ٍC��A��{������Y���=(�Z�d:���>^gz�s��[i�܎����i(PD}l�:}�wX�d��DcoXsچ٤=��`�L���JD�A+��w"�gA��wR��l���V*�X�y�h�D;�L�*�0��)L�P�� ����������j��7��/��/�g�y&F;6�ܮt���P&�]~���|��X𖦙7�m�����|x�: ~��>�����U
����a��=�U�e��@2�|�
{������������޷�n�{a�Clo����l؇�ch�u�d�4�F�UcP1�\|� o������eh�!&���q�����B��en�`XC�m�uy�{�+�n��FT�Β�����q�S���8!@�v�2*�;�*X�$6F�zlL��(�u����*��樓#�b*�1JoB���V��1���3�Y�o#'1���Z,l���y��-r�U���:YÙsj�0U"�0k��;�ZD�*p�F��	�>J�UƯ��.eX�#�7��� 4�?�4O:rd:�H�7/P�9�F�)9���L�z���p�HW:}����E�Xt��N�9��kF�B��`�?V9��Q�,��&N�'��4����^�LC�v�*Ñ��_��/�O�3�O���q�Ȳ"@U	�tr�`�^�C����V��_1�U5GԩۗF�k��KvԽ��+U��s
-��v'@ bv�zM�GK@#�g�ڿ}�n��m]����7�Ҿ��,��}��5����6���Y22�
�[x�.�rU��L��}�H���?��_x?����dz���r�Y�=88N����u�������8�<m-i�jGP��G��4��D
�z��:R�(�.��zwѭ�歬X]^ A���K�S~���l���Ɏq D2#��Rr��6����u�{��a��68�6-�lo�]zPy�<Z����_���[�PP��.�~U����5���8[�f�H����oP/����T��1���H�`���Ƣ�L�	��$�\A}�Z�u�ǏF �C]x�L�yl�A>1bc��,:濓�����s��#�/R�.n{I!+#�@�^�M��6\K6�d��	/~e��*#q	=K���<y.M;K�Y��M�BpS3���p�BW����u�k�jinɮF1�e!�4��0[���bZv��Ĉ`�����hL5|*������ג���5��æIr�ݝ0�YI�gC]e6��ǉVZ}a=В.��BC��ȝ�l'�sP�K?hI������㭿Śb|rݭ�(r�O�v���|����a���}�V9��&���R�����"B���.?��]#5��ܽ�h�2��m#�p��W�飇L��Ž��_�������H@>Rm5��p�T���g+Zm�0����g=�=>��O���F�W�S���>F�F��
�����)֎e��z�)�xT��xy����Y�����Bʦ�����{���j)e�G��0�D��8{C��uf�����	�:k=q��*�D) �V"B�}�W�e����Eh\u:�:�|��(�H�.ryj���<�%\L�M���ӆ����Wn��M^���60r��M�Q:��Rѵ@�f$Ԓ
Y\�F�O}Li���2Dc������Bx~�SO<���s�k<�H������`44iGZհV9G�+y�4ٗ���5�^ƿ�s��X��$��'[9�k_}�=⇰<z����Ƒ#��̊J8a��P8f���Վ��my��|��S���,ci�4� �5�0�$�4����һL*m������A�ך{6��%�{�^�:�"�e������1�O��'�`%��0��;Ic���({k8ݴ���2K�g]�{M�,�M�6��*��s��w�kw+��R����mZ�A'��vr�1x@8-����Fv!:?|�h(T_�(&H#n'�1_]�w��Y��~P������&^�<GŰ����L_�����ݜ~=���k��Ȼ٫^��>��_#�����k�p�&�u�� ��� D*d�,��6�P�E�� �t�p��=�	�D�}1�ƙ�*I/�#��J(S�q��[�S2����IjQ1��9=���mfjU����ZH�G������%��V^ј�Ly�>�ܝ>	ѫO~��6NQ�c..�&j�9�����h��S32~�c���H�Qˆ��_T8�R����t�D��Q`l�\%��Ijɀ�6z�'?���ٓȏ�
�s�F�a��1�D+��`��.����$�iIl";B
=�cjl"�2=��G�$.�1"�'��={�p&�p�&���SO�5���B����5\���9��0�>d�Au�x.:\�U׏<�i����~�\?��zm5��]2.�f�'�]f?l2P��^�9�T����%���&7us^OQ�מ��%�{�n�жc�s�9�l�}��O�"�U-����p=��W�\50~[聳���7߾@�E	��ވS������aM�]3�
B[c�n�\��,����u��F�t��9:;6\�x�������BT���u�|�,)	ۦx�\����+d�4Kj9W�|�5t�9s�ph�%&z�no�� ��hF4B��W��j��(�ZON�3�7?:F�w��&cYޕ��]-�?�;�!Z��c֝�|�m�S�����-&I��g�A2�s}h��z����c���_�+�kv3���4�b�<(˄��r@�I9��#�W��-7���n��(,<s��6�x�v8rκ�#��Ní�57..��������aS�]Zc���4�t���^?G J�P�Bv]1��m.�Ѿ��P;�)�i�=�0�����މ�U�k��F#����A'���r�:KN$!7�]c�6��7��e����t-ZT�K�Z_���f'�Y�J��"]�`��rՀU�gʩ���6M�S��74*0_��D�T+���L(j�Ө��ʯiޣQEEL
C/l�F2��Q�@N�����g�>�R�r�	�k�MY0Pg���ց��y�|:�j�xs����9�dz��<��Us:2��� l����cL.�XGV�(Z&B|��~׮^O7��m�nȊV�7=����8��#���#�-]7�̲���my%,���p�����х%��2�Z�l�E����?#9=`�;"b#4�q[d�̓�%e�``�ճܷ����VX[cT�X(\I�N's-�{�$ʶ�@l�>E�����H�� KBS<Vd��'):��x�.[bۮ>��s���,@�����l�a�=#�pr6@��6��[+i�4�H��"tP�`뫊�\o#�L2j&X��v�R��5c������3��c����y�&�q��ƽ��������'���#fI�M$����ν[u1?`�U#g�Qi38�H�\ϠqV8�)�R/%\�a�_�t3֓���˷9��1(��fv�s�Mf��������4OՍ�|�+Y}h���a��>��H��q��ǆF��̵�@ i���Ƨ�� ]0�p?ѷ'@��3���w�d�$o��w���㘂h�"PQg�6��is���7��'�V�"�o_Xڏ;��=
��2%Cϰ����9z��6望�l���}�x� I�����M�0�5`,:�0����G�h("� �#R��W;���ª89�5��k���F�t�y���k�����v2�%i���c�#�E�Ion���o��F_*N�pސ�$6��GEi4�Pe�I�஀�U̹~���
�"|�"ցPA���F�eT��&��Nh�󭩰����<U1I���k����+G>l��1"�!�Ah��3T������#Ҝo�F)���5�׌|�xί���]��Y��L�)���1��?�vԻ�����?Fi�@��k�E�.dv�5���B`���n\� �� J�Z�ar�ݣ�D>���A��e��J?8w5����'�M����%IED�iinàg87�F�s�Yx!� ����e��\��f��Fᐽb�v��Qb��|t
�5P��o�萩��̅�;g��<d)��K��\
4�6��������t��a��{��`�9;�1�_�9j�
$`gTg��yYOSd'��pڤ<��d�S'���s�ɧ�I���/�skw��6B^z����uѵ�[il����Z�a۲"�&N\�~U2�p�2IN�F%7��D/e��a�2����Z|G��k��N�ߓ��� /�G��mz]ܽ�T�wpO)�l�s�S�%��6�.Q�#'�e�o�KYQ
֞OC�{R�<l��
@D�0��2������6tZ$�"����X!�ա�dTGG���G���i��0���ΜI_��g贇C��{湧�c�!�nl����? 	��1��L���p2n��%���7=�м?ԣ;9 	����pDM��F�a����5 v��أ�8H=�	GF����.�=x(#tTQ��F�H���Z�8Vmh>��`�s���E#�*aia�!��m�cg�^�i2?=^�aD���i6�qX���րE#:�Qz��� $��G':����˷�׿�z�ޤ��{�<���TV�(6��i�5��yT���}ˌ��f�gE�6�KXӃ7�}؃��R�/�g�pŶ��������S+�9�p-sӀ!
� �"���=�=f'��hH�C����rc�B��$��pf)����Y����`�O�v5��������)G�$�xd�IH������:μZ� C�C�}x�Q�mH]o��vz�̉�Eg���;���}i������IJK��s�E��������t����9������wQd��%?),��{�ҙ����}!�RZ4r"�`�d8|jլ��î�ʩQ���e���>ؾ�T3Q.fT�� �`��9s�V?D�,��yP!�pv������]cɚΕ�fT����0����͙R���&g���wlߥ��%�c��^����l�Me��t���6����:���0L�������%�y����AŪ4S�Ϣh�N���W��J ]GN�f��.�������q!�m�[6E;pH��pga��	� �v{��!j�m�*Q�J�����l�:�$����G��%�e�D@B�6V�*��u(���rt��2��P�9�E�s{�����
l���B��׸�<�ΐ2tB��``����Th�OV7��5�#Z祃{'�E�%ŷ��$�h�5�N^��#@��.I����I�q6"�E[lo�z��	�n�Y��H���/s.�t��&i�������~k{�{�EE�,�vg�3�z�å��*bwY�et�@S<��R���hx��
D=�s;L`-�LqP���ٗI'4�U����#�|���Ci��*5��욮ctZ�RpS�u;m���X�h��U<MH`Dæ�lbЈno,K�4�(�!��/>h�牑\[��l���H���'{�����l�2#VPEW(^7�[0ZϾ�*;�"@�
U70�ۢ�ݑ�1fP�i.�����L���eC��)7ZW��x�x��Ml�4���AT�Yo�c��u�}����䕛�E1B�јf4�?�)sL�2}-j��Q�C�}�`�s�;m
8_�����y��ak�K�D�1��r��T�M��.��C������ʤ�8������ہ��A�~�"��q������V:s�%yi��*s�F	U������q��x����=�n���Di;�y�iQ����Y/��y���ʓ���yN+{�̸���P.�G^_�#Í9L�'#����
G�(H�pX��A3-"T��T�F�F£\�Q��>7c INb��#^�gee-MO��L#d����il���Ji4Wxn#*E</��䕄����N�"Z9�"2t+��e�+�>	�Z�yf�&r��@��>��1�lNC
�B��M{HhD%��{I,��3������53���#�5ʸ���r�c�k8_:%�u�6��!�@2?�y<on٦6:��̇���^J4���-׳�sdu���<���e<�la\�H� _�������d�P�O��z4'�����;�j��N��UJՆ���?q4��
�pi5-ݽ͑� �1&z����W�ɞ������}��q�4)T-�[Tc4p����%ZP70���A�:�����{���X�K�ܑ�tˤ���;w6��!m�:S!AD%���#�"vA��"�9�oCi�����D��cGA`���ϴ��VN�O�qe�V;-�Ay<��;���8Ԓ@�C�i�g�׈�T�[�6q���z�F�a����z�dsI*
C]�$��0�f�.�<r���D�ce:�l����w��c��<T�3~W�ij�kier_3��Dd�D���O��	ej��0G5�\#/�0��f� Gu)���X����>4Cx��G�G���ɹIy��������&��0���ڄ��������yY�6��X�j�������\�K?��/FY�5�+��	
������NT#���F����vUY�޹��Ǵ4��8�-�=_Fb�#�	KQj��zp��$*=p`�k�E$�a�����x��m�����-�A�`�<�񭓗4��S5�I� �C���{�^��4]_�����0��6� �MD��D����fD}�s��8�l��ߡ�����?�Cc�uW^C����n��K\ĉ�r�3�'��Ux2�%��o�D�Bڹ�N9sxaKxx<J�p�h�90 Q�OI<rtf�E�D�qޞ]N'���P<>"׼nco��j�e�t6�9P)�8O��*:���lT]hy-�NB(������ ��:�tU�]_>8#��k�nqw�����ge�9��N�;;��D�pҴ�:���EŇ�9�3�v��QG8xVa�Z�j��HS�����a��5H�-.SB@YC���1 X܇�?�!��Gȣc�<'�85�7D��Z׌��P��n�Lgy6���i��ڕk�2�,�ir�����{w���r�����NZ��[Q�"���땕�?�����!@���5 0-x�*�@P��	Q�:|��_�Vk�d˼s�v����0���.�\l�����T�p ��W�;�1��N*"�R� ������cf��O0��Dԡ/��v�11>Q��f�>���Ҡo՚S+k�}���Pe>[�:����E���W���<��M����E�� �R��2����4F�]B�F1�eآ���:�'?V-0A~�K��~�r��cQ��F��<+c�h�,��xz(����z���� �1���gLc
>�٬ȣ>5�3+>7��4l#��"3� Äa)gkWRV��dd��ђ@���� ff� u�B�6�`�E !�����x.5R
UO�/޻�n_}7��W��g?����O��v2}��oQ|/��Fq���k6��!ˍTl�5d��d�l�ns4���j��Lc��U��:�_�>s�ʟ����R7M��!5�;g?�z�sw�<���n/���z���cG�D���������g��:a�:c����,�����w_���qޜ�L9�{�������uS;Z���-�q��N���"<��:>�^��aP��!����2��!}�L`���#ߊ�&�1�w�k���Cc#�},�X8;""���!N���iແkmX4�5�u�N4a�����=�\�=£�I��W��/�V>�(�㒕���l�,�,�ܴ�W-���o�H'FGP�y/��y�Z8g}�U�@T��۔DYjjgƣsm��{���p���M�����1M5��&4�u"v�!�YG�ΐ竓�S��HX��rÒ@�n�U�"�q�B�K���T�7�*�p8�y�%��xpY�W���V"�π��A�h1K$z��7"E׽;Iڃ��g|��M�f���z�x����B�{�W13����uοwO�|���Z���YF^c���ZD����ʜ�t ��ܗ�oB��@�8��6��x��� ߵ�49s�F��&0�>� ��r��t�pO���/�1F�6^��V�S!�`� ���U���^�E`�3��u��UR7nܦ��IFE?���ƑK�鋿NE@�n���
�O�г
��l�Z{7��h}��*��"�1B���������i�=3l�P�h�����٫G��F*c��OE_'B�y-G��{*+RD�����°�$�ap�F�J�]�s��"����%�P�C�Y��J����w�8 cK|��kƤB�4'����PUŧ�'ndc�Bͬ�l"��W�2����0��0鉟�%�P��:��Ɂ]��9/C8<�(5�<�͐��e`���t�&Ց���XJ����ip����o��^yxv-�D8�L2�k�A.P��KG�Q�\��	���;�>��Td���(Q�:��.��&G�1���0w+�L�D�t��Vׁǝ e����t:u�4Uw�ŋ�D/���n��(��W^K�o�u ���<�z�p�vD��.�I�y���������7��T�g��M�WDvP4X"&���4_4!	�g�@\M�խ���H���d_���?|gT�ʡʁ��L{�o�GtS7�E�G$d�^",���<'�N4�tE8�2�Y���nd�=�jF�:WU���%o
F�����-�6��u'T��� �q(�W� ���ذ)�JB����r�lJ�CPӱ��� ���?Fh�h8�.?��;0���Hf%C�c��(��-�c���6���~��q����Q��q��NE�\�X-+S���`��gu��vj4R�����?tD3���U�岭�Q������<��h���e�w�r��b^`�3p6Xۛ��
i�N�΅k�j��2={�b:}��p��JY��	j�-_�;P-�2�7���|$��?�qy^O�@jE6�=�x�̧?Ǆ��N�$[M*,�\á�"�_�߅顙=S�8�߽A�d� EG<�.��K�M���w�T��e�$7�\�y�	�E�e,�;|"��`lh'w-� >����3K���s;P7�p	�w�r���4;a���֜Ħ"���e�v�W��2�7�'з90�ۀ�H	�0�6PZ?���2�yh����'G�t�q�T�OdN��\��pј���HD�gE/f���B�Fj�9�f��Y�u6�D�*���|��<|�s�|_ޚ�<y'B̥j�F��[j4Qh�~�ƌ���W���ε���+��x�6��dss^������W""������|�F����r�<ec��2�r�&hD��Sa�rͮe;Aze�rǝq�ч�{���pŉUF� N-��Dd�c$Ja�5)��'	%6ҕˌ�\%R��O���0lٽL�z񥏧��f�r�N��ݻw��!�Q�}����/>��Iw��vo>r��D������P��W�i�L}��U��G>Ɍ@�h��Y���k�5�ޚ=�(it�'�(nC�l^��������:f#���u Q��%�L����Rh����C�� ;C�ֹ�0���!�n�Q�hp��k[�1����f���qz18��P2_�H�Lsl��$�q�T��t;$Q잰�i��z���16��Q������2()" ���;_�-�����PQ����r��ƻ�f �vߣ)�XP� �)A�/�>�P殐޾�e��s�9F�ꑺ?�kK�jh�U)6ar"��tg�w��*�>��-P	D��Y.�7!����~L��xw����2�)�En
dD�E����M��5�����G�NS�D�����2��!�/�#�lTQ���$|��ie�&�C�_z����c�bބ��0�i6��̮���jS�۱o��UP��n83��4G4�����"���.����	��ҊAU4�a�K�K9�1;<x �qW��'~p������t6H��疧�A��F�
�v	(n�~�>C4��{�h�5�3���O>1�6�0����,6F�v_�m[N3<��]Bl9�Ȇ��w�;Ct�ikhT��1�Y]�hv»Dȯ6���!�����3th��䓶����.CP�[ιE�|��ʨ�e�@����M�#�H��U��aM�e� KY0��[�<`�Z�k>U6N(#�6
6��,�l&��u�G��er����b��_��g��?����_���v��Ѳ���D��Y2�-RX�����r%�\t�:�HL$��m������0�x���k_��2��K/�B6"���]��KW�����/�,$N���|��?������s��HkcT2�+�o�1�h�A�U�ٹ�l��v������Y��A85�U�#Fá�v	#��B8�9��ע�ݵ�@���|�6(�=��a�c($He�^6�ʓ&�
Ľ����W�N�9K*�eR�9z��viM8����,�N�Y��EW8/��т�˳���]�@�۷ɑ����4�\����M�x��-�'��낌���ӏ��4��9�Eo,L�W�}���D��0����
Χ��\���J[�F�{�y8﹄Ní�|uh�f��}),���;�k�qɎR�ו��8�D�[�������cф�M��ӿ	�2���=�0�PD�T+Ɂ�}�7_	o:��ϟ��� ��L�{���Y��3S{�ۙ1��\��Y�
�4�2�=q�i&��K�CJ���GON���Tk�ԏyu���S��[3���f]mw��9����ѧa�ċ ��VV�MiT8��h���􄜪}9tu5��:Ģ3�����Ԓygg�P$�2������t6H��F}ܤ����k�Gwc�O��"0�d-Y�[��O��"��2�@���4�-�9��ذ˛,��y�Uf(3pbַzYO}��J��d��s�ػ*�0�����z#`{LK�臬e����ݦiR� 筍kb؃\����aȵz��:^쇵�ٻ�=����\ë����T������$�қ��ɺ$�lB�L��y=D,�E��=`�
0�P�o���0�:Zk����~����_�b:ql4�i�n��6�Vl���ϳ�m�mY~�W�"�4���#�U6(O�h�X�@�2�����"7Qȶ������'oÌ�9��$=�[o��Ļ�8Y����4��޻7�/����p���V?��v��|ϳj��1�v�4-�9j���r<�%^][��	�<���]p'Jk�P��)�#1��\7�C8�]n�5�|�����G�0�!F.3P��_��)�����X��Ըw9��K���Ɏ�.��9=�����,k�伾�\�C�y���k�F�J�^g�]�Z��c��@%�zzV��0�T�M�<~&��C��!)����ŉ�tn�������[�[B'/F�nai%���u1��ʍ]�<�;ߑGzg��(kW4��k�+k�����~uv�����{��Rr|v�:�=����9����=)�#"j��g]��Ą�]rZ��C������M�F���ˑ> =Y]�?��~p��$A��I.d�p?G�K��ɱ�z�E��p�o��m󩋗.��t��>�&��:��>.18
��ʭ�����tk�;-m���q6��p^�^��?���U�r��??<'��QD�'�5,s�DuFAW6�(X�9<�C6ػR��MY�\�Cg�iY�����V��>�2{�19�i�R<ٻ4sp|��Z�M;+���G��'���7G	T���E��h�ej�/ߴ�f.l75��ҏ��;����t�Qgݔil.Ru�3ી��?TJ�f-��ّ�|�e�ֵIx�φBD����������+?÷*x�K�O��^{���`n��L4}�r��=��a�|cg�L+�s���7�{�aU<X;"u�1A��P�en�&�_�q�@�{_�e��o�GϜrZ�'��2���߇���:���,cN�H|η;�L�u����2����y�
&��'��[�&r]���	�kR�E��#i�p�V�D,{g�#ojd48t,���7碳�5�ѶW�h!fF�|�sDj簬нg:.&#>�,F��	�"��4���I�2J�\mt2��I�C5�6��Z�Q����dα�h&�M��X����S�\�����f+=\>ټ���;����g�_�ŝ�ee���z^wQ{�gu�N;)�g{�K�����r���H?���x�Qq���3!-��Ȋ������T�A�y��q���i���k��GO�����#�P��IH�7��&2#]NH����85�i��`�����D?6�/�k=������?ŋ���={\��ľuUgc��OŦ�t��D�r����&E�6���k�:!��9,":\:���&�lQ�z�>]���>���?����>�� :fvpB\=�;����56['U�5�ҝF�f�����Ϝ�����{w���M'{~s{�4�z`mb�X��D��ٻ�!�{�2W"�o%�m���z&��6��,�>��,;��fC.k�\n��? 	��M�]Cc�#w�]1��'�79����������`s���收1��)���̍��&��f���X��FGzcl�~���=�}�B�R+��w����!�$�{�!�����t�1Wg��a,z�3��?S��:q#+!<��8K�s�����@�R���3R#�؊�� M�+c"[+�l`E[�V=�5���T��F���� �&hD���I�K���u�6�PQyn:FA�˻�B�C�D�1#���LqdO&�hu���O2����+�捛(��8vXm~�FL��1-�<f����{+�:��lUBz?��P�Y��q���覂�=y.�1��ү��6��L(���2�d�0#}��ߌ�Q]��1����_IS�i,���|,o��۟��s�xuh~2�(ݩ$���	_n0cz�p�ZW�t�f6:}���;0���if��P�w�IT��ghN�Y<__�aCVL��c��F3��߸�c$(���^���]�| �Q�����i��K6�����T�����։��= 2�eS���$�t1�0�E8r<�� v'��p��3��!��XG:9�>��Z���Cц�3"c��
���s���ۘ*�x�l�+bd�����L��ؓ|I�t�'�<qB��8�N������s�n���X#�+GS������3b^�Us0��é��J����t͹��ۙ�^��G~>����G+�TF].J��8��V��bg�J����{|��{-�"q�}��{�ôpLf�Fҧ^�T:|`"���I���-�ۋT�D���)e:4���f��H,�~U��Y��"2 y�<�O����Z���]�[Qgz���Nz�:��X�5�������&��p�\{q�Y_��e��,���C�)�����]�����}��m�q�R�5q�>�1�y`]���hM,o��i�v�KP"�JH:����#4r޿o<���!".�쥜i��;W�����~�r��O�gm��K��`�6$	�[ϋ�Р�r�c���<
CtL65�Ad�hc���J!+QרFШk�����5����6`��CDm��ҏ�"��M�Yn�P�PC�j�m��o��A��QJt�&)G"G�hU��%b�,�p��Y�Dğ�ѱ:�����[EL��}�t6�+�92��\�ӷziqy�s�)��
Ghv>xv�3�ȵ�e�����ێq��,�'Tm�lx>��%t��[����9t ���+�����y��O~���ԯ|>�ݻ����{"Ǎ�F�o
����ƫ߂���p����ә��/�QX�'��?�X���t&à_�|9=��Ir��!�����7^M��(������I��W��P	�*Z��o{)1��M\Ѹu���b:4��f�|&Y�)��l��U��@YG����s`6;}<�#B�p��53�Ϟ�wa�ߠ��GN�C��e^m�J��wa緅o-A�p�1��L)��}?d5�*ျ��`ɔ��=���k�uj�,�&�R�:��b D�goL*���d_E~�g��7%�ѫpD�;��09*��!C���mfv�D
��N�4���al~�@��\q����{wn�A0��:m�E�Z� �9��TX���No�:T@��}��p_�#|Z�7�m��de��LTg�GԠC�!�Z�2�zP�&�f'��s���m�'0�q�8���}���Z�m�H�X�y��^��1�N���m?;�9��?ݳ�P�L(з�(�Xq-y�w����0��Ыݴ)��� �)'����U��|�)cOW����8��2cA��䧲��ԘV�!��I�vA^�^�� �{���OA�%X�4)�?0�Ϟ�Cg��k�=[��Y��*OGz�D�s��0�2�F��L?G��3��o~��Z+Ѡarr8��C��8�@�[q	4�&��Y���J�c��ˀ������$W�ln��jt� �$�h�%2i��r><r�U4jS����bw��&6� u�B��WG1Iޱ)���<�>�m
�r�6��k�kr ˊظ���&�`����&kH��*oXfm�� @��2+����Y��C�xB|�-�3���mn>kZI*��S����];9�0X� ���rL:c�D�#�[y��U<:�q^9Z��q����ϾU���Vz3�:�����0n/<�4p$9��A�/�6���4�$�ur�+���(�S�O��|�s�}HE�%���Nљ����~?Z���N{��SG�q�'�Z�;W���K���0�l��&��ߌ)V���8���o���H\����܁JI�P�x��L:s� }��F�߫�&]���a�v�k�_aJ��Y�_��K�yr�v���u{?MEΤ�Qg�w�{@��K���l�B"d
�k��/��Ȥ6��8ՃY^9v�f�/��lKk�0O��X���<R�=*�����Ǡ�3O��9R뼯S��Z��{���=��$��lr�<Q�E��;�p��M�����c���2���7�E���4���>,�ÈY{�kū^.yz��B��l���^z�����
.3q6�KQ�k�ܸ�O��T�ߓ��>���@A��F��+?�?z����S�D�b���CSp�@u2�C��o$�.m�Jdx#Cަ l%\��q����g�����O���p|T؆~S�h��q�
t(;k>���A��d7���"&[h�����p|NJ�p�C���Q����v<���.H�}���A�� �"4��>�2��$�IY�8��+���� ��$��?�<d�}(�i�n.�)t,��45�(�"�F�KݩZ���^D�P����؎,ʦ��5j,~��"���%Ym�F�vt
�3:y���vvw#s6hg8�Nm��WU��Ҍ�A] i�ƏA0��e�Npo���L��L�"����
�L�k�����AP�",��D�]X�hacx��NBVO��a(Ҽ��R֥�|D�����a���_ߧ���)�M���#}0D���،�H#>��i�� ��A�
�(���5
��Un(���s�թ]h"����W��M�<���*�����L�Pɏm�$��q"�P��nnC�i��#L��3��;�Ӯw��>h�׾�=zso ����󏦓����cy�����g���b�H�	s+KK��|�f/"���Z��� i?�;�u0�#�r��W��g�{6=��@���}#�\�s?vx?���� ��6M>�H�MO��{�ݨ��_�?�������/xe��ԘQ����p�z���`׆�l0��Y���R�~+�'�����m���E?!��`��,�Zc񆬄s���C�p���h��u�|Y�{�jq�ϻk���������GX�t.�b_��N�cD�sG��ßX_�5�#��8`�m��y?��FV���g!�7P����'"�
�p��3��*t����NA6��{���do!z*DE���ڬ+&)
=�&�fY�����N8s�Zg�9L���@T��@�X��<u�C�����y�=W��q��94������Wq��d���%�T�x�ڝ��#��B@)���@��0��I	��s��� @<R�`�S+ {p�Y�SZz�n�̫�T&�6���i�;��6��,�#�S�"�-��9Ň*Bg�t�q~����(w��B���Sȶ�̃�@�كD�ܓ��ai��Ju��R��*�@);[y��l�hroV�yb�~���i�~���;�����IT6�aQjt���p�V�"���bx�z���*#�MSe�X��f��˦��2Y�1}���],��� 5�[{�
Kj}�پ�l�N�p���(�ql_iu]��\�΂�D p��'��gTFA$s�n��+�ȳ�v�!��%�5���W���FF��[�*�_����N��d{�L��Z�P���!!eeyTϗ�m��}�J�v�oM`&��(.��W��{��Eo�6{�e�Ca}�Ԟ�t���t����vz�߇��wd%t�Q��o�}�$�� !a|ǐ�� i�`�m�Fi�O�����\�.��;���o�St|���(�Y��I���`��"=�'=M[کt�� ���hR;<`�܈>ܤ��?{�aK��Q�{>G�x��QYb��̞�J�����H^�|�9�p�ǿ���Ty��A`�A��џ��'�3��ȸVｋ�{�b���q��/��1�'[�p����+ rƳ���ka�#*��8h�v��1x>O̟�$���;?�?�Э���ڳ�K7漚=VnD�<�u�p�@؋b'kP���_�l���N�<�`H�:Ƭ�d2�t��edM�6��и��&c�DT�a�M��+ȸ����<�,��'ݻ���@����iehYÕ}��0�#�u�0�Fy�~:b�0�{Z�/�
�Kmܷ����-]mP��Ŭ�v]E�
?Y��bTW���:7:�2�Ȉ'F�ʠ ����Ed�z��h�@⦑���ׅ�
n���Y������F�F&"���A{ L�0ǲA+�#����	�I������l>��-�Q�ލB����z��P�A�����������.�b��0�@mc�3�-��F]M#0\�y���U���ı�t�:}��! ��?�n�74'HT9{��J���MI{��r���è2�'V*��yؖ�mn,��$��ڦ��D�3�14�Qà�����
ύ =�����#J�hݺжd4Ks`#c�������U(�g����^%,�%�ĭay^@��d�K�3���/�Ґ�R���<:P�:����az��U�9�o_yI�S�E[�BۍzY��k�s���pUA����5��Q\���M�=Ӥ"��[�d�hY:$2��ޤ��n�=���qj#�O۝.�OP�+3���|� �|���xX�Tl"� T�M��2�m�ק�YYZ�8><��.��FI4��K?�Ŵ�z��7K�9�f�&0���w����:��:p.�Ƀ7@	��A������.�� Ֆ�q�w�Thݟ��3��9r�X�ε�i�i:oi�HX2�萐�3�g<�lbd�7�����XVs@��F��.{��Y"as���b�U�W�W�OAZ������5t]v����,�L�|u���gr����8����p�>q}{�#�C�Ĭ:�Y��.,͑�ѐ��aw����9ɭr��"h3�Bגh��x�و�o�uep��67Wu�kF幚!� �!;��8�p�u��^	�<"|��93�!S>�?�1z��
�6�n|����[ A����:e��?�� ��P����kbf3����~by��L��nz�����HW�K#za�@.4��o�uw��]�/�reN�z#��ѾF��z��H������{=�9��-���!Cfɽ�F3�2�n����K�%؆#B������
3h���1Ɔh� �Q&.��_�AgJ������[;��l�L����H��z��b�W[�v��"�i��o��7���{�`'��cG`$o�ӏ�:3Z����E|u�'}�{�h�@4)�4c�a�l��B�@bð�O�ׂ����U����	�L��RU�X҃��:#!s˧��*}�."9qg�)�~�J8	#�*j�e��ǎr ��]�_�#�%��������oGF���ɪ�)�b4��(����jF��䒤�$���i�x�|�ǳ�@&�6���^fԢ c4�iёМ���ܣ����x"�;���w��=LO?�D�Y��V�ַ�G�c8��t�*���{�v��I��p�.Uw��%��{�4��q۠]h�Wei���~�f+��F�Ʌ߾7����8x��>~:�o2Z�֯2�㷿�C8��z�J�}���6h�{c1Dk�:��L�:7zV ���xf�B�]:KDB��KD�A��ܹ� ��]��n`�/�܇.08f��?i��=w!���!����?��QO�"<ʄ�/|�Ӯ `��i�|��<��c�,���w.�7'�=�]C�a��t"!��@'Ѕ�m��c�/�oF���a�"ES��X�F|� �[��p'��������Wk9���a%w��S����v�NI�����=&�]�p��q=���'(C�q6��~;��Dݠ��:N��a�����u�a\�_εߛ�S89w0����-G�}�w`���ՙt]C���-|-�/��:�׍6E�D�L4pny��o�r	�:�NST�A�����H�]&8����gi�t�5�7-�W"�蟜	�r�D�D�b/���Yg�z��U4����U��Pz���u�H@��Zv<"?����E�p�E,�Y<�u(�ևS��R�Mw�+!�	�_����[��ro*:F[[��ܐ*ΩVԃ��2�(�����#�p�U�����?��KQ�:w�,��h:vd����z.�����p|b�N�m�k������ŵt�v3ݞw�'��
1�x�6f�[��t��jqv�I"��� ǵ#l.�\wn����&������(':�<e��=Bl��Xv�<Wgoս*^�\�ZMC��
'��n����8�0�UC�N���6eG��@���%k�&�5c�9UZYA���x�+�ʫ�%��r^�a������6�Չ�܌6�0���y�w\T�11���?�����NG]��O?�^z�t�|�v,.��?�����D[�ҋ�?��;{�'�>!�w��q:�Nw�F�ۿ�?ŀ����C'�.d�y�][�"����0��?=�R�09�3�.��}�t���4��Yy"���� z���-������\��XZhn/p�}�{��$Ұyɱc����x$���^Т���D��S���]8�~p1��Ǳ�nݙ֧���������i�=�y��U&�-��}��P�|�4�i�ɹv�l-M$bB	���O3&lU���Up�En%�M�$���ôLV�n9��Ʈ�3�����F�ZaP:uВ�������\�w�F�:�fFJ��v�15C��ԑH�}p�F8k5��6?vvfo�!3�Ն;`^>�Y�A�זIk�����5�{\���:|�0��~��Aw��{�@$tIuݺ����aC��R�$�^�)B5Gr���1�3�s�D�r�&&��K�p\���w�)��vA�Vl��J����L�	GOlRn���hiIe-�5\�����wx������N���%ջ�$��L��_$g\/YSŏr
��C��.%��|��@"E�gb���W���U�Om�	8,V3�07�Rb������2��f{x��;#8�V�1�yǘ����1���l�������(]��uX�F���PZܐ���������nݣԫmH�gK�-��<WV�y��l�a��#h�S��ˑ�Ng��Cx��|������9��r ��ψZ�Q�-�'�.s}f,lK]�n���*��Mf-��I�B��Zd=���������/�,�GVN��*+��̤��=tx�묈|�oGO�
��$�Y.g-�O��c�c�B鴄��X*M��lb��A� bt�0�w2��z#?z,r�����ӝ[7ҋ�=��"ߋ����-����W�h������O��D���>BW�u�rHJ��p����W��jL_3��2վ��_��U��%���4E���%�t:)!���#F�j�̢�eV����`�׼8܎��uo+��W~/�w�c.��GOГz��=��J?Bx"a@����1��;����?�"���߭��t�&��t��.��$�i��t�@&L�Ds�Y�f#V=B�C�x�DǱ��;
���}�U���Q�r�*�F�� V[�b��*���3h�+��oTgh���1H��Y���eHf�|�޽;��7���3U�׮�� ��A�(�1D�"��1��=H���q�c��G�uF���8��i)sǞY��Ξ'(�;������G&v~h���y0~@=�g;L�
G�ja�m̺0��w�s�ߛ���,�
H����ӧ`��`��.=�#���e�~�x;-o����!����Mp.2��9׏NN<�I^S�f=�s�BNdl����JF=*g2����#=�w� ���49oT/z#��E1x�T\|&�r��nҒd<��b�����ԛ;c�����9��(#ٻG?9�ç��ZIo]&g[3�:��܏��Kts/]��L�r=ͭ�E<�-r������<{��wQ��˟��s��V��2���g<jy�.�朢	K�7��7Dd�r��_1�H���{������N��6ca��=�P���G�֫u�&.�rbSDUYɆ�ז�]�����\^�P����|c�ge��ZF<�S��C �\ͣ�����x�U�2clC�B����su䄉�Ǧ���(�A��w`:}��X��W_al�Uƕ>�N=�(���LG��Д��Ё�fT+ghA���O`�oG��g�|"��|�;���$���215��k4��|�m�{�=�Tc��Q�*9��qmsvuIH�s4��.uP��)��ӽ2�;�;���!�Ћ��(�e?��_��m]N�<'Ym��w�ʍ��k�s��w��3��~�!�1��{dO�z=OP��eX�0�(IE���ɐ�=F0v,S�1�&�ڽ_�{��B��:�r�����A<����Z���u�n���������:��D�NZ���A�;�'OF�!��X��k�15��"��ӧc�mo����jz��+�7���vY�2�}C8�:Y� :Q͜��p��b���\RVE�q�dG<�@�V��E`lܓ}�Q	ע��J'�c�uz��{O�}���@ڂ�"o�뉮{8F��8i;����A�γ��d�-�8��q�M�&�#���YƧ�A��nI5Ys�`��&��<��������{�-�MF��k�ㄇ�����YEϡ2>�O�'��Z����\)>g����?�Az|`ԣ�:3Ғҗ�@�؇�L�c����>�m���������C����0�b������CE�2u�M��`Eұh�n��Ǿ�ɦ1]�FD/b�@$�bstl�wK��Rm���Unz�SE�|�����z�18�����aZ�a7�}72<�܉.��P&����KS���W���;!��/�����99�*��Ȟvg����=��
���k~8>_p�e��>��v������Q��<6 �5�iD$��.F�Un4�N?rA�41���	m����r_x��K��s�1��ߩ�Hw:q�D��'_�П������(�1�3zy�շҟ|�;��Q`1%M��%?7�\Ow6nS�l�=��k]#"'�߻����@�*���W(��E2�\*�D߂p����<9�=�������;2E����O�yL79r����z�c�Pi��q��8����X?7GE�:�~�.e< ȋ�B��AO����e��j6(y�P�����S;rԕs��YH[G���0,������d磏���g���r3>�Z^XqjJ��w�]�r�UI�rb�TFGgϩgN�k��RF�.���:jM"��1}W����4�F���n��j}�pƵv}v��$�lУ�Se�;<��;0��r�[��p��6�;\Qy�X|ǱN7Ea��~�J�����UxX�c���6�����Q��2�\�._��M���K�}�\�U��j8�̛���T�s��^��*C����x�����3*7�/G�!��daf'�k�<�̉�qs�����]XX���0���c	�#��O�Z���`л0��]l�c"td`��z��S�?�)R�X�5f�I���9T�M���a-��N�nE�9JeQP�m8��2;Dh�����=�5pvd,iՈ����Z�����z�����؅����U6|��,���Goǹj)W['+��wB1�"?�sN=��{$�Ă���+w�D��9-s�:��#�9 aeӁO3K�s����U]�����|^�;9��>x� V�e��T�*�0����ʴI����e�ixQ���w�yV�Tٻ����"<�T�A�Wh�ڇ����^���>����Z�I����7ކ47�����}�#v6��r���4�y����W^���PA��O�	 E��5���j��MJ� �շ�`�9l���E��;V���tTp����:�p��T�_��g(�;LT����ۯ��:k�DGP�An|��EW@�VF�ȉNd=}�{����ch�Ҍ�� fņA_� �ʶA���	q܀�JU�sސ=0��p�S�y����S�r��j=U�6�!:���笸3��y�Y��1���mB����3���Ig1b5�μ��b9�ߧ�ߊ	T̌BR<	�!&��0^�}Q����:�����N�� �g��'L�/��N�;��W@1��,�����=�l�G�����`�ee�w�6��3� a�)�B�K�6*�s��7b`�|p�\�ѱ�#8g%]�v�~�4r�D:���c�+kd�VŐ@���Xi"J�>;o���k%�]�*���S��*_x�GF�᧕G�}��W��B��AB�9ɜ�xs|�����s1_�ȡ�8+��vA� zF�*�K7��U�����{�܄������C��y�����Fz؍�#�L�Ƚ�BpI�ǅb��#*��v4"�ګ��,�Ie�����bA��9B5���$6��Lk@�Q��k.������jE	7R�,�݀�9'TO��ig:L�����@z�-�N�f�=��lO�#R)�8��\ܒ�Ā�ܐ���{�9�������&׸h]r�\����]U?e[{f �Y��ʌ�DB�֝�ˮ^Y��>[������85���9d>C)���n\e���7�Ï *�^����O�lS�x.���+� �gYK����(��i�Z��p��\'im|Da�*����fA�~n4(��1���@?�#�����*��೪%��!D�f��W-}�� ��H���3L������R�o����Tjo�%��Q����*��cS�H5i�@k�m���s�' b6Q|"2�:'8>��^wJ� �+��1g���c?i���$�h
aJR�m�o�IÔumg]e�e���R)��?4�Y!w:�uT�e��]�Iվ	�?V�Qn�~}�{͙+݊ ��~�\!�<�z�˙'�Nئ����<�T���^����ٍ9���7ixt;"^�"�̺W�UT-�56y�_*yT�����bLj<���3�7_UE�_9�g����S�q=љ�����`l��Rtb��w��1ཬ9�� s��4��_����Ѿ�N�

�E����r �-�p��,�2Б�"������f�iaD���k���2�A�
LG��"x��sّa�ǀYt^3"�<w��m���ܼ�F�g1H����\�^ӊl�%��^��'E��w`�D�y��D?D�����6�+��<���(6���(E�Xfh̝�4�"Q�e�I��zn�|7� ���š�7W����G�0:��%Nؕ��.C��
jx���Z~�JFff.��j������#����^�$:{R�$�p;-c��$+լ[��+�"_V�0�1ؘΛ��7Pp}||�#���UJ�~�Ыt�v��e��0��&N��]�(��%\��X[[F�[�x/g��OP�.������Y!𐚊D%iŅqa��LO�>�����s9qЌ������Q�(y��~�Ԗ�#/��y�0�E�-��_���.o:*�]deXUu�Mt�˽�EO�:�'�{
�����?�ĉD�����W���w���f��=F{U; jX$�<j	���ko�|��-"�z:��.�=��=�}��W��^c}�ZE�8���h��z�o�!�!&�� d�ē�=���^!�aJ}����%r��0��z�Z�.2�n!�?��O3qk��R����8߽���|�|����a�4@�4���!:ު��Ó�ԇU��L��Z��:��H'���X9�<�NGC���u΃8*vb���"
s��SM?U%�UE�L܇<N�P�mR��C��'_�x:)ν:q�����\���2w�u��W�Z��e��c�����O=`��r�'l���gL�䎇:9��R�A�c�s��Ge�#�w�Ȗ��&a��K�u����z�)�².?a����8��L� ��6�m�{��{���D4���mrYo�/$�Z���MR�C���dnBv���������2��!(�j�N���e���Ι!O�����
I�`���)�84l~P�T��f�	U�,�j0@�1�|�~x}�hܻ{Z4br'|ɇ|�M����u��7/_e|�Q��Kn>IsI��1z�x�uGO������$6�T]p*L��c�.�M�RjU����xWRq06c�қ_�1��9�pO�$&��ػ�m��Oe���>[�0Φ|r��f����K��zoTrT�&~�y;ޯM2r�'�gE���l�_D]�kV�U�@x��<d'ō��������~"�)*
��9��g��]kN�����T�0m���5�}�א{�g��<X���'��C��o��oR~8��i���<s�Ӕ�����iﾙh���_�ٴ��1(f��@|z(���ϒ�勃WW��s��5�����K#=rpo�s�\�����rg��6D5[hv�s�v+�t�γа4�g�<R*��E.���}������@9�c9G�O}�3��'ǁ��0b��̠:0�o��?������1z�?��#UyR���;\Wo�؋�F�L����~��ڃ�DZ�t����[x��Q"�����}Ϝ�xl��P�9����עL�E针��hB>qo�>��������Jp/�1���b}���(h��J?�Qw�屫���uHe:!F�ƛ��N󘈘��N���\f	��1E#��{��S!�e�)c-�2ט���or���0n�Ͼ�zD�y��g�d�v�GE����1�E]�a ��>2r�7��H9�;)�%����v._FF*�M����Rb��i�=��=�#�>�v���V5�IY���W��N���\"��$��9�t�%z}T�x�����M�}��i��+"W�A�m` c3F��t��n
nQD�o=�7X~o��`�	���d=S!�ٽ���2�to��R�5J=oA�=Js�Q��V��w�R�I���!����d+<��L�z �A'���\ۜj��vix�)��n^+o0�R"¦q��Q��n&��m�����=�~�?�<6�C���v�7�=L��##Мc�SU��U�gD���=K/���22��5��5>�V sw�S�;+�e_i!v��ߕv��.���9O�6�hW�b�U�|�{*�:o@�5;��d:�';���4�p���_E,�/vf'2�0��:Vt�2�y"j� z�1E��^��D5�K:�܆�r��vb��;�g4:~yO�x��pxV!�&/nt�3܈�0=�3DgG��ƭk4~���a�v�/�����
t'�	��NPw��ϿH�j:���\(���at8�۾J_�e��u�Ɩ�Q���7�z4r��>��:y�<C~'��Q�H������1��ҥ��������ν�V�'Ϥ=�G]���bf�,���xz��gXd	1rO�\��M�q�f2�~,}�ܫ�3���~�MӐ�"�-���ٗ�L�	��L��A<ξ�A�x}���{�[��׿�o�ЧH��M%�7�u �j�(�[LU˨���Ԙ+ha_ｈ�#�Τ�\�.�$�aV�ѧ��,s�����Q�[�*�ؽ�t9'��X3���Ǟ8��x�D6��äh9�C�҅�OV���"��f4����� ǏReџΞ=O�M�Sj~�j�^��;Nx�q:��p��\ّIpվ���2�ɹ�<��=�EO�)�㾈���\�y˾`m	)w����8c�{pY�8�ΤXY��w�����G�3u�	(�&�<w�6�����i/e�Q�z�Ug���8�a�=�̯��Cu䫏uQy���_�Z��#b{[��z˺!沮O.�Xx��0��>��M7��g���O�+��!��UĔ����v��£���Ҍ�F̬�<V���"q� ��� K'XN�&�ue�\0F�14��25�2��W�8�
���ƊP6BL}�L��S�8CfC?�z���R��F��Ӽ�s���vʛ'� *���Zc�:G�Y��66���q�\�c<sj^�d�^Lw��Oލ�:Ƽ��$d��#�/�떍�4��)=OٵC�5'+��Ӷ�F��(���!���^_��J�J�a�g;E�i�s�������t\3M1��=~�P�E�_�cXI�t���۠��.�@��]"�4`�{(9s�N�����0�ֆ��]�z>���l5m,�M��ۿ�W�2��l����C]�a�F���{��p/�9�#N��S��ؓ}��XB��sr���>_x��������9i殹x���0���|��t������a�k�+i?��Ǟ|T
�HS�����t��Y:�O߄D8	j2̐�	j�u<��>7V���ܽ��9�pEkQﵭEM�X�o�ܞ藞SP�|�<�F�[5�lU�fX�hm�i��a˫4���u�i�KT���h�i�{�aF���Y���pax�(i�ҿ��c2�u;�T�"�#�FbV�
|�\�!$t��ѕ��4��Ng�r̟��'�k�x����-��������Ty�d9o��\G�0��5���ӂ��$�'��@0��}{銈,u�61b6��V�L��ƷM'9;��]��o7���Q����"��R��4"�7��C����\3�BʽXom;?�)�6%���z.�HTܛ�;��<T�B�K�Lv�z&�z Q��^�ϋnMG_����)����T~OF�2A�~��3�� �[b�i�]���q�7�х{�� �n��*%W-���Cd�wz׷j̀{5Sz�n"���hّKғy^K�r����܌ja廜�Ю�
N�Dr����gr��e���4Z��!��&6Xz���������+��+\�L��(8|��l�c�g딬��.e۫FN<�ad��U^mؼ�H\g�#�!d���|�I��"w�W�һ`����1ר9)��~�^��4p��޷o߉}�zn��5�,7����N��L�%*3��ԟ�o�FqF���T�]�M�՛W�+�~�aY��`������n�Ay�մ��,+�q|�ľ��g�A��8���5R�ְ3�3�R8�C���?�v R�c����F׷��qbRTUde���i`t��O�D�^K�����rm���̜t�A��W����?�����E���0��j|���v��W��t�#Np{.=KıB��2��ƨG�vȈ9�l��aZcMi��0���V�^��� ���a^��w�UGe���xUד�x�f.��\���^��N����bY��A�V��%v:z�No#�h�:��$#j�W*�ƿ|]΅ǎnp�1G�9��aSO�@�b� �G����h{;<2��6��=06�D�;�\%ne�F	��H��d$s�;w���1�<cT/]�2�^OҨ��k�+l����Q�X��`������V��A;u�"ts�}C3�I�K����y�Fs�Uk0w��с�B�;@��M�_�Be���M��} .�v��6�ݻ�:����،�>���9���c��*�nm�!)I����ʂ��d��y:9��r:ݔ��oP�Fi�h���_��p�\[�@��^��}d�'�x�5k�u>TU�Ik;��\�:p�|?��)ҡ�!��m��>���C�?:v��3�@Vԕ��%w���aγ�OF?��b:Pp7�p�W0�9_Vh,3^,ܜ�	D�Y�*����VT�BCAt��m,�]lP�U�����2�ݏ�>����q���UN/�E�m��r9��(�.�������o�`^T�~��mY�v�y���-s�*Ԫ����ݎ[ű�$6�p�"�-�f��"��%��g������#�9��:o�v:56=��ݲ�Py��F=�nA�@�lA�o^����׾G�mO4��x�YF�j#.�֏S�"W�L�F����"��)Ubf���d��"����`�����~"��ܩ��[o�{���W������G��Q�1	AU��s5񛪈ҿ��s�YAi���Z�����J����~��`��4|+��o�)��'q���L�1�w��)��u�Ht3�U������1�O�!:����i��;��`y��ōk���Z�=��9�����VV��=�XN��z���(STũ��r��N.!��*gV�1T'��i�Nw4��gGT�-:�5���,5t�i2	M��r&y�-#�����|�e�a�������g��m�o߾��x� x|���x%��x<G��i�$� ���2��*������'�y��tz���A�He@��Y�Zx���2F��wD�Az$�M���B�Rk�0�+�8�D��ip��	s�7q�MMeҠ����u��Ȉ��#Jg����qvGA~N�<IJ��{��Co����bOLl�y�.�hG�,�auD����࿄!6�s�s�N�0|>��R��5�x���1P��`91�j�����Z/Q����B)�>��1�zf�ğL��] Z�Xu ����0ʬ��A}<4����=ֶ,�d+O1"L�ܬ|\���'y��^�s^u<Q�Jt<�Ji�W��>��Ex����A;�r�&ǥ����v�r�F�� 	�!:�5�@#&��aFw�~q���+%kE�<Ɨ�AI�	;������r#�|����!������h��Fj���yɡ�Sn��|�}�g!��2��_�x)ݡ�:9m�k�C��n�i�e�l��^~�&�P��dUO���Ї|�(��.ڵAI�6��'_�z�����)�sD������ݝg��
�|�ȟcحrDaF�J��z���۩���tg~�{���;�+�d5������Ì����#�NyM8V�֨��/���P�\�����t�����@�0��o}�[1(�5o�O}�S�I:�E-2�W�thd�(b���4����=���֭t��Cm{�6���;�������R�iQ���fz��7 %����G�o�
܄W�5��v�����M	�~��)���ʱ����Ga�-�]ű�A�f��鞸�9����p`b��:�EB�Q&���/׍{�cu��e���e� �?oC����[U ��g@9 ����q�y���C����h�kt�T�w�Q˽"J���8u�T����v��`Ȼ�5(Ά�ꢪl�	�#b�,rR��O%�Ÿ�j��%q�������_��ݼy�gv�:�"���>�qtC����-Ċ�X�������@�,�?p(ƞ�q�LL�q����=��R��{8��_#��>����=�!��{4��%���<�.G���r��+~:v9&6O�d�T�5���>�1p��Z��qo��Y�(C���p�n߼�=s�* +�q��Sʺ�A����G4���} �����zsd{�5��޷�|�V�aHd�g8.TQ�����\�QAE�w8��#z�Е
�u@Lya����.`��3ѝq�전>B��\��H61��t~�R��s��;���5�l�ةw�܇!H��(d�f�s�Jиg�2	$"P��弝LV_������%�F8G1Fy���۾��,�~�4�H��6�O,W"���(���Q�K!j^U��ёp�o G���K����(��/s�{����U �{�΍��P�f�,�I=���Ŷ������u��u�r��j�NR(��A����qZ O�&�/~��4��>gڿ��;��D~)�о���G6>2�u�$����r+�[4��mm�
������'N�Z�D�k_��{�6���F^�����*���A����~�k�FIΥ;(y��z�V7�D�<}8������H��_���,�sm]0�q�������O}2}��[����c�ƹ��&�K��3�r�bz��m=��\<s����sl3�r��ͮJ��k����7��#`6�y���T��8P}B�U���a���ltɑ0w�~׶�QD�D��i�+��:�F6�=���N���s|��4��=~�h|pb��2\��;9p���H+ؒx��Gi�j/������e�IwVh,1��W^#�s�>O�� &�  @߿z�%�r�E�<cxWWX���:�4jqo��c��Q<�W4�1�䵍��Q������V _�!_���L�o��0��pY�Ni4�721�1���>;{�lZ�w;}�/��g~�i2�3��@<ۅ῞��!	�[�����:�a�ÜD_W�J�u�Gu��J?�U�&F4�S����Bh��D��^a��>��Y�RNG)�,M]B�����Ξ+�h�O�9U�;�Ý���~P���t�0��z1LyZW^�y��R��Zbmi�ss�
�*��X`�T3��s��s���y[�����To�����a�6� `��h�R͜��ߕqvJ��p_�g���q��Q�^q�$�Ԇ���mw7cH�4c�8��k�P�tB�Bn������b��%�H��R�9J��4�*��(���F�����Wc.Ԯ"�3�N��FG���*�W��U�v3�0m҆U��Qo�?�s!�EJR��]��)5R66�X���ܺP���T��wL�����'�Dc�e��m]� ��l��wD#�Ӈ2�(�-#�1��.�O��L�obh���{<=�{�y�_��o�*���P�Y���0τ��S���Q���K�^cr�ݯd/ۀG�A�f��L�r2R�V����9��ˠ᡼!%:d���b�{h�W��e�*�>������˫�1t�ֽ�t����?�7=��)��D�sN�Wg��O|�}���R&��B�m��a�<k���Z���:<N��9e�?�����/�wY�N�N��d_���[��7r5�y�㸹ǁ�u�c	��6`��TG�q�%܃N^G��#���
���rg�B�|�.�������KW��7�#�� ���k���v����9u���7�*�q������ud����s�3�k8k�������X~������$�p��?�K���͕�쉼u�χ�/���sI���\(�s�8-����8��^p]�~(�]G`��;�1r���Pj���Y!�S�|�Bb����Wz@�~V>Sv�ׅ�="�7Dֽվ��f�����W�B�ބ�rCx`0n=�J��=T���8	�;oE:Y!=���Ơs�v[u!��nN�d{�s���UD�`L�A� h��1�ܼF�z���_8x*��Sv�l��u6]�����X�kHr��:�4���d�p386`�L��	X�����ߟ�B:�Tb�x:�6ŀq����R���t�#sڈ��`��W��f��@�疙9��EW]E�ѣ>�Ϡ(�G�d/��.@�$4{�ˆ^ �Q�h���c�����yB���-���]�m�n�7ڐql�5�FLAH2B�����;i�!�^��D�^�~.a��M��oI���F�J�KKx��a"�IF�.m8"���瘔5Չƛ�+igdb�i|��E����N�,�:�=ޭ���T��}��f����(��R�v��8"k˞j[s����0"�hʽ|��q����v�zI���_}����uF���ޤLO��#����Z�^���ι���}7R��ƶx�A
�,#TW�G��n`�q�~��E΅��{��a6s$�ݢ�o���ƽ��^h"̽���1V=����Mk ��W�/П�繺CC�w����- Q��0$��L����@f��2G��GNEU�0��~�m��o}땪�RU������]H���Q�Đ��K���L�N�n��R�E����;T[�u�%�����Z�b歍�={���7���J�"tZM�,c��B��w� )�)��H佽�؛샚�hN�!u;˶�8��:D��$龱W�U$"��Ȝ�N�!t�"r0��c*B�hG��Bg��3�r-l�ZR+��mЦ�_�~:��I�H{�y��.`'���;���[�hdu��ߟS#��*8���s��\��0��������&;��p ��|�Y��誟*m�P M��|ti�5��Q���z��0H.}�~J�6�����ͭ�16!61{�>bL%"�Xe.*����Z�MP�D�l)�c�C;w�#�[�6�ϡLʙ��t��F+����&����b�Z�eF�1N3�����N���'�/_J��*j#��P�vF�F�Swʦ6'��ly��1Ց�$�P�Q�A���	D'�$a�rI�Fh%21�l�YX�C����U�[o.t��{d�˼�4�1�nr�d!	J���Їu�4c�s,��m)�{��t��T�'�wӣ'�{���/<e7�w6]���g?�I�?�z'����&��� �>r0����+o�M\	��nh-��/�җ���@�z��(�:�b4E�a,<,�1�]�k@h4�7�K��VwHq�KU|*������_���@�1������|��my.�X��'N�"�M�Xk$]8w�c�� ��v��(1�m��SGN2`7Xn�]J��o�Q�j�s����15��8�z2%��,�}���t#Ƞ��>������r�i�k��� H�����_������d��&�[L����!+Z��,p#kj�W��_�W�b��K/dh�{���o���?�/"���Fp_f?�Q�(#l1}�3R���7߁}~!]ۼ{�9�O����K���^���������	62�.Bg�"~ s�k�*�o���y�����1.��"���7�*�f;3�]�̙�w��x}F�����}�����{�W�/Goź�=�@���[}�S�;oaۙ��zq��H)�][���bE����r�}���>�_���;�O�O�g/�eV���mP��`F�L�I���r�W�{':��[Q���C��S����e�<� �Fu��-��:D����>����οh]�K��*����{�4J�U0R0"#��A�F'Ӟ�T􊸄�������t6a�&����F3s/�IwX���4lq��ш��N��J7W�?Ls��\T�N�yf(��+c6�cpUFl&�f#P�������-ꞷP�}���N�G�,��+*RHo� �|d�#��pݢfya�u6�i�U�g�"-qst�g��7�-�w4d�Ǿ%oY���������㘟q��(d/�9?�۷`�Z[-\xY���cR�
�s��(�Y��;�k��F��Q��J���{�3z׸�6��Ds�(�1"뀾Q>W�m�t����%�3ju�f)F���[0��hr�\�w�|�hMp.��ޚ��i�r��ݺql.=v��������=��Y�S%Z���L�j�b��sS�,׌���H(uv��U-:\M����D�C(�}����}�u3�޿L� �e�Gg���~`Rr�������T,Ҥ����sms9zD�`^[V �J���A�K��k��;>�D�4�	'�{0 )O�Ns5��7"�?�ǁ����8�g��뷙5�à�aCU�&�ڒÉ�	�O ���#���w���������N���sW��>s�t�C�C����~�Y7�����}M{2��n3,giy;���p�W)a޿E��.�>��6i��6dɨ��Xc��_A��$E-�k�r8�h	x� 2C�*���"`�k#Ĝ�nw�t�-�M���+Y�nv�<���]�Y{F�~�id��������0�w�6����kئlԡ4�� ��O��i��8�i��7�x�4��4J��C��`�qFYU	�|N�T���42�ѹ*2�x~.;"�b���&4�C���c�Q����N��o�L.�X<>��!��^��cjѲz9n<�Q�Cc��J�t����7�n���$���m������hT��H*o2�d	:�����qF	�1�10/�XX������S;0u�BnӃ
��^�*���DL�I<6��nu��jy67��;d���d�8���sΞ��N{%L�n�sf��,�$b8=r_y�Z�[��A�lAL3����;G���Q�؅c��ߛ�]cn�a>3V���!�k`��ڐQ���(�c��Z�񝷧'�ϫ��v�1$��K^�ƍ����(x�M�%ʙ�B��IG0����K�>�,p�X�G�<�V(͙�&ơ"�H ���"���ppT�ܛ��B^�I�h"��0���^Φ;�<Ɍr�A�qm�R��֮�(>�;�Ǡ���+�џ��1�ͨq��>��t�Ң���:z�<�8�����*�D7(Q#eC��Q�QyW�t|ns�4��q��>x -��$-ɗ$�__�&�2nL��������ԏ37�3H��;LΛk��ܐ���a�9���Dz��' ꑣ�fr�鐺�K�	�a��l����Gy2���O��Y�|��)�D��Zԋ��@F���e�?�L���G���VFM��Ҭܝ�}��q^�Y����O�_]�@�FS�^�1��=�h� e|���XA�5ʜ���}�W��b�򟥙.�y{��D��1?�@�H��%pի^A'>:ʹ���#��c'���#��Y�m����D�~б�wJ�&d}�Ϩ#N�㻧��9Ώ��EΣ���[��\��BW��Bz'P�wp��|�����A��9�� ez^7�Μ!ec�"����"jw���eԐ�4�}% ^�$���Iv���k�N�Є�φ>TḎ�Y�<��-�M,�3���*<��a￞�N�4=�Dd"�+�Wu����N����RK�jiwIQ\�
):Ё�Б�CA��`��[�r8;~�̴7U]�]�<
Hd"3����~�7��F���PY��g~�5�����^'(�%���|\f>r�;��F��ٵ�؃������ƍ啙0(�3��E�tT��|p��܄�j�Z�����欢@k�>��K�dAF7�97�Y�%:�9�s^\ղU��4�~UvIzs#�J�\�Ŝ%ȩ���N.C8��Q^��n�H�!�y�T��T����>�\�ש`2<�O��p�NaF5<gP˜���Bx��YB҆5bfW(Ց|�2������JqԘ�G9(�+X���q�on��v���@8j��h��Y���D9����K�n�5<��� ��=���KQw�~�g�P���>���_�J�w�ys�C���������¾q�9��thң�BZJ�а���Es�3O?=��Ю9�������v���!7X�4��g�@f�q�
Up��۔�T�$�f+~��ÛG��E�ԟ�|rx���az����е�����ps�
uʴ����`�݂��|/�_�[�=�n�9L־�R�y���e{A��4�
��p��eD���@�kX	�\O��6 �u��x�eK��g�}p���I�ީ�S� ]��ͺd�.�v�L$*�|�6 �S����q��~�i/R&�U*\���(�]�ڰ�Q�EzWQ�a��XU斲9x����<f�~�;ޓ��k�4W�;
}��Q�@ćcM�0���q�.0E�d����x�{ɉ��X�W��M'�lT&|����bIS�F�@���B�{��n	�{;����~�j��:��QP(g�ؖ1^�����?I�q���B�������(�Mj�I!<��/R޹�F<�{7��34��FV=zγm{�`_�_��T(�y4�'�)-��Vc`�<��(h��||�<J�v���}ָd�+���V�|��y6M��12���K��t���D�6�Ñ�.�w�&٫B�������2���k�~��7O?s���Ք2vS8��N�Z�g1օQe������ʱ�g<XZ�|�H��o�Za�딭U��.�,,bU��ϋ�b=T��˾-�r�xZ�S�/�e�����9�LP�!�� 5�=z����r7W'���&Q2Z��w%��c0���~@���+�|�w�����؊Q�m�ok��a��5�0LyC�E*C�~ӭ���J
��r�)��2�$�����<<|�k_~����#�h����9:��e3���|>��zj�m�{��E t�w#�9h�u���9B�6���z�ס����h
� n�+�B�۷|���JD�1iZ��q��>�8YB}��z�ں�p>aK�ȏ�ﴷ�k��'>1<��8�d�N��7�
�[30�i��)�bv��	��	����g�6�D�0��+��`6n.�lf��Ƞ��ʶX�6�0/N3�z��N�
a�
�u���m;��h����3Dv lK�4�&�g��^��^�!s�*�� �������_|�TD�!M�#��/рR
~AǫT�z���&߭g�:����Ɉ��`�1�e��	�O�M�zJ����P���g����Шb�뢸�:�]���
�������ծ~�rk9�d4|�J�l��#�n�|�֍�)��"R1E�,PsI:c
j��B���(���T�Q��q4
<�3�w��wϺ�Iń��J�A�_�n_�o�li���x�ﱦMH�� �J��t�̲>w 8���dD�`#4�%���d�_���lG��dUqD���!9�d3�%������-�P]�+�5:u�2?xe��q��b�,�Y2��9��7��;�J�Q�������Y-���������}`�+G�x�܅���&��'T���� a\�Tt�����Xҵ���"X�
Z^�m�,2?k��Ŕ���Rj3&;��n�FS�k���y���B��@s�jcT��[�j�Tv�Λ����b��&
�v�n�y��Y�:	 �p�
^�2���o#x��K(n�d�~ X�鵌�H�1^�D n2.�
��m��qL�&���sl���Lk	b��SbrЗಥ��zVU��w�p4�=�y;^(FBp�põ�'��z�R�f�eeW;��D��gO=5�c`��]�]n��C�J�x��3\���ԗ�:��y�?�2��dZ�1�kF�w�ߨ���Tw��@@^<�@�&Bt�8k`e�@NOe�U�ч���[i~2	�ε9�J�1�)�E���]{����6�}f�XR#�E�hH����$(�mÆ�;�q��Ls�m�6��O�g���V�f��wNCT2_���:�����~�����v�\8��;�8��ȁJ��8)�-���Fֱ-P]ɩ��x��Ž`�9���v�LԮ����?�O������o��E��VX�R��u�^��8	㐙��~m�b;�8ѵ��N�6�^:���?{J%N��8ƇD.*�ԥ�`7�Uk5k�cAl4�����x�+�c*�x̍�)�����"-_���Ո�������c��:
@C[�R�����n���K~�d��D�M�)־O���W�'�s�N ڻ��ä����{]�������?�'����I�i��<z8)�*M� i�^X"Rr�H�%���FC "Ax��·���D���^�k��#���5�S�څdX��*.M׌ �̴�ёwV�po1#J����t��-Ґ����Ż�ш	~��`b8�	��c���ZF`E��}!W����*��y����������O~a��]E��vZn�ƑTy�8��c��c�LO5�.�Zd.L�F��|�,?�>�A��֭G� !ͬ���:������hZ�wPp�Ϋ�����-���9����L\{u���]�y�V�u��%S�� ,���<�==�
����رɌf,���&;u���2=���\��m�нvcs�����;0��6�Q�·��XכһË�[|ۮ�����B�0<�����*8S��<t�=A�����-��tj�7���Q���
����'�R�n�E��_�o��,!4�i��e���8��[�p�O����}��%4�O�g��M	�"��֕rk;e7dp�@�X��V�y3���xف�2C�;�N2�;b',#2���-��
��1^�.����E>I���G�f�3�{`���<�p���R�=i�����&�._�1�2�f�E�!���m�F�8sb�v�h�}�3,<�
����'-� E�$��%���S���H�yZ�J�>]R�w��,�w�<���c�7�G�W4����0~�$�~h�%9"�mi��3�#��g�J]{�f;�	�k4k���C�|���'2�I��ly���\�Q��m �M�1^8�:���@Hyq��To�%����v���2fU�c��_y���F:F��@8#d��w�U�8�DFDƔW�:�ڊQ�)�Liio�4FUƞុ��ٞ��ַ�4L!{dA���:c�\d�8�z�Dl:�N���=ua8��%�^��i�p|�u�wX �֜ ����\���I�C��5���`��a ���}�y�x�&޵W^QNX�Wk�c U�� c<��%}���T�<6��7��'�Rb:%�FX��`E��52'n!�
�x�>�V)t��#��c��g����8O�r���V ���ڮ�B�buǕm�p�Y��a�W�]B�[����r�2 �M��B��@�ZJ��.Ű_NW�8�(�p\]@Y��XRѸ`Y�Z�IQ�5t�Z���I2�y*aTr��1&$�H��ROE��PEzji7��c�	�����LT���*���ɥһ�n(U�{H�β�bh�\$�w�Y%���$��ң��;�����{ �J̑�'<��@덳�6Jx���/>��':���p@��L��c����<�[(�1=w�<�gsk޹á��Z�Ks'�o�O����P&W@�K���$gj�F&؂dM~x�K̽mu9*��fm��Lx�e�nBO�9A(�����Q�;i��O=1>�;�N� @��78\<wq���A��a��.�'�~{���� �x��&���?�������+.��P�� �׮��wT�����`�\�K�w�����.�bVb��]��9/�C?�r�!��Է���~+F^M���Qk��Ͻ/�}�	���n�\�^\&2a��1@��ɯ�5C���X\��W���x��'�O��F�ʯ���5$���2^�aۊU><K��Ǣ�w�1�r���Ly�}�:\Kw4D��h�pLꕪ����k����zԦL)�r����6l����%r�D%���s*<���#�t�����E�d �XP����%�>�����I;����s�u�ԃQ�-��q�F�0��1�R{"M�"x��0?T^,
�����لe��.�k��Zv0앫�e�c�{��ks\L���p~�f�G#?i�ȍ��yQ'٤T�~�B_��JGȵ�D��}���0�/��6�lɫWn([H"��nc�Nccl��[���y�%��Ƕ�3�_y�����~����]����O��-�լv7K靮CK1�:����G�g����%�W=��j)3܈�2g&zSkv	��X�z,*-��<
��+E^f��׫+�5��@	~����0���*-<צ*����}q+��-�w��+7lj�Oᚐ}ج�5��1zPe!+Nʤ�-�9�#,�}�;�U�� ~�0��M�bO�ڋ�* �27����{z߆�7n!�ņ��L�$��'��%�%�(9p{��@hNH�Bn�p��'�[��o�]�����fix����f�5��-��׹��P�T�8&H��&��~d�ZH�� 6��F��ܨ��Ry�kϽV��)���]#=�RƜ�E��8�Ǹ�0�D>�^�&=�ُ=2���X~�:��ɻc\|�+_��<�Z��?}8�i7ф�u��cPt�#��ɑ�|v� Q��\��ћ�����o}�ۑ�W�x�1I.�0j����S���!�'�}��j�I�$6�W_�FO�I�I�dSP�
��D���]��)(t��rҘ ]$� \ �\�r/ZFI���������[O�"s��x�����R0#�(]��6�%�*%���$��0��mp��a~(�Z&���m����L�Գ��c�i����Ch�{�0|�j#�]��Vx��m�)3E�`l��a:�:ߔ�73.�p҅��Iz�d�Mk�Y�}���+_��p�=D.\+J���FGa�)��x��)X����f���f���!�7�r�̕Ke5�{v���Ҵ*�W�qIu�i����!J�(��x�A�`q\�?y���+SLڢq)J�7�`��S�~t��_x�5�;�OS�_��
�{�H�q���A�J��ߢ����<t����_�����N����GLI�D�R+���Va�BC\��Bw�ּ���]	�߁)����V�H�\e(�u�P�z�-�%��6j������k��P��0P��!u^D�h;v����<�ތ��^��b�x�mg��o[ϓ�U�Z �p�\|�i��<�PP�}��A��,��Wv���q%zj�7xm�0,�}�ӟz���ގ���n������ �!�v��e=��-йN"ף�n��Zw�2���(�D��?��'��Ƶ!�BӒ�I��D�O�?I{�9�������c�/�s���f0�(�J�͒� z��5��;w���g?q�����c��L�hT>y5A�y�5��$�C2�|ψ�mČ�	'5A�o����3��N)�Jғ�������a�N�M��p���-�����(i��۷��ӱ'��m�6��l':aG6��pϮ�i.C���Umt���Ȯ~خ����p��ùc�������e�W�����D�KD����Fm���Yd�^��4��Nb�XC���x�x�[�a��m]�L��rr�s��w�v�&��m�u�p��2!b�ph�+�q�d1)Wm�l�a�2���B���N�m;�O<���ڊvZ~<iA���1��
\ov(u�w�X8��	��V��Pm���T*��> ���<W1,�s����hqJ[_ז�O��jW��Z�B�Z�[\���[ ���։bg��pΞL�9��5YND���^dYK�i�濍8����0��geLg�3u�J�ƾ��-��,/�(�
�Rk�jP�b�l����ޠ�dR9�翎����t��0֯��p�����c��.̽{շ��p��f�Qj�f	C۰���[�зl����w��k�w_~���$N��l�U���%˺<�0"��V�	aC����V�YU�1d�<�N�Ŵ�XQ����0��&w�P�D���Y]��,�p$ǳU	��뮞Q0h���X�c�k6���_ee�0W۾�H�(�2�.h�RD�x����u��M���~R���yE��uF6t�a�Q�	!O�2F�(EXM�W�����a�4t�/���V���=����?�j�
�OB|xI�7oC�/S:�)eb�jl�4k�1\�%����G<Be�2�q�W)�Zo�6vٻ�0���gO��0��8�P���?s��u8��:ӿ��"��9b�IGx����:����?L��4���u���9T��f4E��;,O�&�J�>5S�ݔ�P�.�͠�"%��o�'h�Ǟ>����/�J���TG�ݯ}�K���\��7a����Dr�S��.y�s���:�w�(���v;~�V�G��<����꼝�!r�OS����[#:�^�u؄C�_<�q\��=l���wE��!h�2[	��zܖ�i��� ��>i��:D Ԭ�� �ÆV����@�u�dp�`z�l����p׽���?:�ѷ^"C���f��nlD��(=uC�2ѻ7�S�,��,���TK|�}�a��WJ�0����N�MˈD�&UL��P��x��{���"�g�QD/fm��~���S���Q�c�#ytx�����������I����B ʠ�d�>f��+�%.��E�q��2�?�Iq�E�V$�A�L�)��.�D�b�G�3S����?]�k�EG��<��M$A�կ�9&�x�r�����YG���K��4Q�H��%�������=G)��ĝ�O���w�и����EW��w4K�3�R�{���x�{�|���G��� �InZe��ٽ��5Ž�s��y�wֲǨ�U_�U*��
�o�R�ň�*KH
ei
GJ�D���X�k�O���/�����ԮL��S�{��5u��nk3�͚�4��U����_6��\�2o��x��c������q]R�������{e���+�&-��9��q�ׄ��"*k����F�v�4��$�|彄�S�Ns׎�����?��%C~v�j�������h8r�����(�q)<���F��/������<�|�&$SX��U����CI���7��h�-v��>�9��%r�o�x������?{f��W??�s�]����3m�̋��?���{�Mr���m*«E5���F��<i����>�&m�a+�b��ukC�RBB�g��~��/��}����cg��|c����[�;�ޢ�����W py �>�����W_(o^��n1 rw_@�|���"U ۩8x���<j�(&s�7{!mI���xſ%;O�9�!(-+��)n�u��%5q���VR0�8�aX���gO �˽tB۽�s�Ϟ��"E#�����4�y��=l=��%h)��"0�I|��6�a��l�pN/�J �.�3Ģ"&à� s������Sy�t�.�|�*��0ȯ��H׼�(%"oi�J�A���?�2�3@�%�{����Ç 7�X��p���˴Q��P�����B���V��R��
{(���J�X�1����#�-M�W":������҅k2�7j�g��&��Y����;y�"��e�2���Bq���q����uu�5YX��B�wR1�W�YƉ�B���֩4��$ұ�$sc�@இ��ި�u�r�Qƹ��po��3�k�Þ��U�{wm9���?�������;R$�ۍ�̏W~���jG+,�{_�e�zy�	�6����j�r�}Y�1ݬ7Uv�����	(��[H���:)p
<g�iҚ$���Gf57C�k^S�#��0x���!G���1�sݖ	
��M<��w�G�K�Q/z�3�M?��K ��s�3�`a#�3�����R:��!#��g~��_���XƽlD��s��!�;���c�B*��`F�z�ό�}�ci}zLj[!ZٶmԔ/�` P��a~^y����{� ~�S�/r���QH�ڥ�=w�B����e���,�kMX>2\:׳^'c��/~ƶϣ$ls�n8����Os�i�f�9_��?�좘��⪬�{���m�7"���'�D���V6�]��)
~�o�wf8z���*���^#n�&#�҅m^�������/e�����9X�^�zI7���������;qb8��4as�l>v��������K��z��$��e	͆mZ2N��3��,��
}��<9U{ �~�V)�5d��z����CQ=���o��o�?�di�{�^�#"��h��q=Jr��q���p��� �����KKj�~?��ہ�4�,�0��I���oL.�ߊـ���(3��NT(3S+�V�W�֬�:�k�&]���#n�WSf��{�H@�и=����/y��̺`�v����/�w�F(�]#L����w��%�5�c0r��,�*�5J�%E�]k�Y����-T$$����)�O���;�W��5Gc�	o6�jL?)O=?qz����_o
=NA��0���{�y��1Z��]���%�)P��a��ņ���c5O^CZ,�<^��������ڰ�ͮ��1�x�#%:A��߁�2�w�㱇�g�x��g����I9U<���s���p���5�Y�a�Ҋo���D(�n�D��k��c-���dE�w-A��J�N��1�7c���OJ�������]&e9�)˙��[���4�n��zфI�,m���4�1) �qC�l�����[u��C�}<�$Q���<%B��]���ᓟ�ܰ�/�ia�(�ؓ��m��wJ!k谾Ma� x'a�250C�Q�b:��Q���h`9��۷w �߆�� ��V����7�%�l�T���xQ��̅^ ?|  �^ji׏�Y3[���nS+~c;��_L����K�W�f��"͘=���A���Ͻ@TPʒ�%Qė.�^z���9�O~�b�,��$�n����a����Ry�z+ˤ�Zܤl7?Í^�(4��Q��3y�UD��_��%���w �}XU��n�p���p�<쮝	�26���/e
]�"FM����?:a�}��í7iȂR���Y���O���V����.,�N����6��OS븧P؋\�d9r�/��fHl�&��1���o��'��U���W/�?>9��֫ÛP��Zw=`3p$   IDAT ��sg�W@L\���שHI����GR�=�(q�e�`]�f�ӻvS�G�|����%j�W��H� <�&�c3F�QV+{�4\lz�r2�y�.\EIHH���Ű�J/_��h_h��C���-Q�D����s�6
�:|h_�yS����ktE\�f��zɇ�������p�,� ��n�<���N?���kF}�$ʽC�h�"v���E\E����Q(<wu�U���uu�a1�WO��,��~N� �}����!�}#�E��T��	qT���~���!�Ns�]$�˂��֭���~!��됏S�O>{���1���Dy��`Xo�`o��L����رuәO=y���_�z��.�!��M�#��4��^�9*:J��p��5�\u-�����%���Եqr����"����a�u��z+�o;1L��p�g4��k�߷�f���-]��2��ɵ&/�񻐚�C�O�y����� ;��#��	"�)�w�>IXj�*���>�R(���X��'�dNQ����o��ɒ���N���ƾup�I2�	J�P@v���[zQ��L���.f��P$S!�XG�}3 .�Ֆ��x��@D:G3����{(���Ո9�iǦL��s�]��~�>,���_��㝆8��u�'��ƅ�����2���w89P�E�^<:�-� d����C�_���c� d���7�S���E�4x[�z^JŁB5kb�e��hS	�9Q����zs�+�G���-�3�#�-s��= �1<�1�jv�}�5��1@;��N�B�(�����e8z�I��g>�����4�X�i��.�X��g�NtK��.�t�ˆ��v������7|�k_L�ȵ�X�D��(����}ï}�K)ۊp��ˍ�,aI�3�x�u�FB4��W>W���L�<p�R�Y�SD{6�ʄ�%@?��7���^��v�wΞ$�����o�9n�zy�:�r����/
C9Yb%��{F�]��F��Vߔ���м��i���>o��=f��b�S��r^:OKң�R�~6��K��$G|S�ԩ3�(cؐ�غ�ѫk���]�DK� ����LYY����)y�#������@Ύ͕5�S��5P
�=�w pS�~4>�m��y0ߡ��s�Oc�})!��}s�^�ޔ��9�������e"(�]t�څ�2GqF��LR\`�X!�*J<ӚXc�	�vK՛C�!Me�v
�[�/Wqn�
vv�3�s���M�J���u^�;����gXf+�֑��=w���o��KO3�����.�{X�gnҸ+�rU�ٔp�[��n�}}1�3�e��Ϧ�!%[��RSC�y�Y 5�D��S7)*�M�a�B�V`�5���$A1��U��Psj^��z��	��Pg�!a�(�Q	]�Ra�s�E&)��kž�\��a��|�S�L��	���g6�?��%����5�^sjfʜ��b�n�粘Y�q��w3j
~�I��aa-o�x%l�=�^�u�� �}O����E��^�
��;�E �Ea	tQ�o�]��Ӥe���xtR��g���ߖ��Ǐ#�~Iu�e�C=0a���}P�.�+�3������a���a�P�8�&���.��>�3 �g�tv�4���p�R���j���kU�W���/��ʩ7�o��!]C��q� �	� ���D�e4�"BO�G�<$�˩`@^~�C� ˗��Z��zJw2����w(���A"�|�u�*,p׮<�;%Y�� �nP5p�p��y� z�(3���݈�߶g˰��^<�}H�5=4�{��ݤCLsT�9덥��B�S��gݱ\E� �S��;�4v 㬰V}t�f�T�Ft,s����MM��=�=�%�ћuo�r(ίwm�Pǆz�1�܂��_!��@����$�	W�%�(�%���3�g�\�S^�v{=�G6o @�r���m���ڿ��3���0����t���*��|��!�q�L�[6���h��S^KU�p|tye�j�-9��+�ޝ�ȟ�%-�V��U)8���X��w�=����������Ż�h)��$�M���X�R `S���L�'0�&Ѩ�qN���X��A�}׃�Ҏ��bL�MCvc��N���S�S4�_!�b.�ֳ�_�^�^>j*���=OdpE��sy����y�����f��q�,��&����@�+���"$��e���������K�}a~��tr��D���圜�!P�pܧ�\�Mq����QZ�Vv&����Z}��t3զ���B^�ҵ���Q����5�n�W���lFØf[��	[ī͢�+��r(�(v�=>7)�Ǧ4��
�i��(�4��#xƳt)CH�=�k7�bl�M�N����>�ȣåk��}`-�C�[ o�^PP�Bɰ_Rd�^��Ԯ�s[��קj��
l�jyF�-(_o���Fw/{������\��z��Ȍ>�ƶ���ˌ'������ߊ�sp��t���������!�R��?}щ��aɟ�y����>?������3������C����jQ�C�UJ�n�'��8ky����k��x��w��� tS2�]��%�QV�����MWs��i��g����)B�A�kt��o΂!=�e~0RTl
s�3�߲�������w�G�/3^��F]�g!I�a��O�1���&Dy�����w�	���!L��庶�-MX�ߵ-k�P���}ix���׿��a���Q�B�v#,),�~	ı����qu�J����q�4M�,ˤ'+�y#&��W�g�̏�����5��^M��p�ܠ���w��4�n(︩:�M>{։Խ�B�y+9ߔ�aL�/ʧN�IҟbR�s���xQR"��h�}Ɬ�N�$��=��m{��)<ދ쩭܇��}�ꆅ��so�Э��쥌����Pi�5y�z��H9A�+�%@EdD�Q��v��.��&K.���,H�y.I���*4ܛ���'�޿���ZJ%����!�Iw9&�.&� �OR�'���H�T�:�K�j�rxb �4�Jvi�o�Ny��?���1_�B0I��"'�UvIQ=�a9�v.^G��&G⸭��������:y�FiН���:�� ��,�u B7Q���kM0�����dB����+� D����/�f����Ͼ����჻�ڶe���k����|�Y�Y�|1¬��K-��b������ب%Y?���:(��� Q5 �lY��Zzx��&W�V#_%�&+5��ZB������ZZ�*�7L�MKī�׸������*-QAx	>��3C��~�)�0��g�ҙ��~�7~}��'?3�M���?�%߷��������JjcJE�D�δIHVȣj�+�h4�'�rB�MIHf7��G�=\V�r�9�/�vlx�$%*ze�ъ� �=�����*m�w?m Q�����
'u��[�m5w��-��?��?E!��瓠��s�F�ʹ�\�Ar��J��V�[�.G���K��g#@�c����pe�S-�IP�y��Q8(W9�7m߭X�ב��G*@C�x 8m�⨨8�"��fg�ۆ-c`�*�OJy����U��u�~���a֓En���s|v�I#E�k��/�>�w���O=	z{wJ�ާ�t�70�j�v&����t[�V��}d��Pqz��yǍk�*aRk�mt��·���h��}O�a���s�'IL/�4�SY�G�ʬ��84U��X���]�z�f����w^SI�$�o%��G]宁gT�p�5"H�C��Q,s�c���)����¥�wm�wH�=GD�hɲ�!]a�K�G��rͨ�
x�fOڹ�u;Ѕ�^/?.Cɢ.��L<�R�Պ�=�_JFm���w~�H�|���F���N�:����L}P�R*H��%]!�`�E{V�FS�Yl	����j�UT��=�h���Q=�F��%���á8��Ð�<0m���^���%o���I���*�C�)��͒�g����ȣ����~]����ggΜ9���G��w�;��0���[A�'���2�^��K��O�����B��ҁ����7���uǮ}����z��g��^��JE^�Qy�U��|�ۮ��s��*�Z�Q��FmSb�TyQF�Ik��
�z/a�&L�'Ne�{��Q���d�T����"�L�eI��9���T�CKڒk�> ������"��V��!*�x��	��+�_����-�YM^}����?J���h��y/��-��Q�������ס ��]��6�1�d����9���}�<)0�9~��9(IסP���?��0�n�<���	�ʾ�Si�zk�Z&��EU0�P�i�r���pZ?��(z�P����������ީ��׶�'��硿�x��mx��8��MԺZe�o��@޴��-���XBG���ـr���
��J9�ETt��4����+p�V����e6��D��M-���eD),���M������TET�W�[Ě(�ϜuX�4�l\=��:���(QQ�z��p,�����~j��ٿ��9؆kW�%�:0L�x�_�b��q����DE-�E%������L.�֏�[�KC���3q�~bx
�)��\g�T
�5���������fW!������*�5n��?��Ea���q�:��Q�����^��d���*j7�n��+�y��S�� ��`P��|;������4����5�*��!KX�w �`����FH��f
$*�~��5���ipV�ըb��x�h$��M@a�A������8�.]:�:�+���g�Rr
 �c��O�%2v  _��0)�2�zym�%�#s_t��=ȝ�G�4�w��?���vqn�I�H�5m~��M��cvX�YX98��!qg?�H�2��o����O������M�lCf���ʱHxK�P���&�5?~bx�w��w��K����������^=1�B��ށ�a-��)�Z*Z��a�����^eg��?��|���6���\ˢ:�94=|Q%�O+�𼻕��Y����
���h��i���q���"�=�0*h�ɍ��k�(�<��@�u���\�}0�݆bs���[g��t��3i5-p9�}��7�W`esL��'$��1��иz5�p	�4˝y��l�QR�6��1��=�Ǣ^�l�����s_���Ly���)�E��� ol�4�����x&֏?�t��{���zX�.&�.��yʵ.#D�?9��fx�╋x�(h��' SQ ���+�ߢ��p�#�u����y��e:�� hs
��4h�M�\_�Z�.�i�L	Hm���lԧv7+p���x����5I� ���1s�G��*�W"6��XVS�<�&�r��v��t�T�(`1����=8C��0s�u�BL��Hs##��ٍ�l� pr�|pRx����N����u`�v��`=;OZ�����gZZ:&�M[��;aw5Uc%^��DՃ˘�xd�a=�Z7�Ʃ�� #�i��{ډ�d4�j	����S�yH�����ϕ���A������:ɕl�Xe�7b�x�brR�ǜz�@����#�]Z����C��F,����AX�~����X�{Ħ*0ĭ���M{$F�n*:�C�y⢦�ϖ�o���eZ]q�#�zİ��+G��%V��҈Q�z��ƹi}x�H�87����V`��#�脚��]�V�()������O�E>�qSUE���p�)���[�Uhf�t#6���w�t�4�j.a8�h���q�5M#{�Ƹ��F��y���qw��H��$N���˟�Kߓ0e�Ͳa����`���8�m�9�1��իsc����?��//8rd�ʆ7�����%�'j�Fb*�lH^�Xÿ.�"7���
�<(���КMu��X����aǛ��G�'��煐�Nu%>�@4o$�X�IՁ
݋�]��}�@d�ғ)O.����rb��K��i*����9?=<3Ӈ�SL㍢;�%:�i���کKo�{�@���}��a=1���ئ����3W��|����
$#�=fd�KƘc/�/�kq�5�����|��+�P2����I��N��)�Z0��G����pmx���ၻ��m�$jq�w��'��m�zʓ�06�K?���������[�3��w8��α�c��BJ�^}���_���߰$��U?`Z�{�K��?2����õö}���H�_���w2,���7�d׳�Ab�	�rME��g���6{|�0��+��(�|�<k��݆��`�`|�"ѕ�aˆ�Y�z{��	�TҘ|;��;{)���h������g �%-�yB�7�X&0���ݧ��vq}�v�Q������瀢���(^���r7�n��u眧v<�Fj]��.�x��&��S
?u�*Q[`�	(�s)��1����Cc"���@�4)����^�͂�gM�g�R#ʗ��� F������MR����i�k�Gc4��8�6j�ǝK�
�v�(6s�+�Z1�&0� ^Z9Ri�n�t9e>ηQ�	��@	n���y5ũ�X�f����u oL�D���c�TT������\C���M�D�8��K�Vj)<(�q��,F��=����OzcF��w��8K:�{��S�v�؅��X���?�1�	쿆���7�:B�[!��6Ǚ��@�h#r`'�4n�y�ell�BX1��:�ە��#�ޑ
�|��+W�����Fk�u%�7S�g�k�;�e�*���� 	�]�����7�?�%8T�0E��WCI[~��S!ބA̾Ֆ��a��vQ�6��@������+x|7�ӕxb'<ͩc��*j�i��v��c\�7*� ��ZK���r��-����٧ W9S�f�i�T�����)���QɋEl���v���k4do����/,�0�����-���K����^��PSl����K�\AP��K%J����>4R�6Jƭ]C$v��\���K�;��<�0��9�W��?ǂS`���\`.��֓��G#���
�/_��'oE�l ʰ9\C���6�w������@���Ȟ8y�\�g��g��ǟ��ߠ��������<ш�B�d�̟�Ռ.g_��g�3s?�N`<Qs���%m+V�-�6?v7��6R�Gͮw&�����dK�k0�8�m�����9kՈ��@ ��7�P�J����W>�E�4��R�r�{�H>r���[�AD� �8��:x/=�w�N���c�""s�����^j���KxY���R�!	ھ��1<zs�̉{,���3o;�4��GaSa��p�����)e����*|u�"@*{�k<��V� �|WJ�*/<@�9a�I2њ2�Y*oհX-Em�<8� �v�u��=])�� ����o&q{����}�Mj�E)���-\���D�d�xp��H�m��|(��ua�o$"b�}�X��˓��T��.����īL��z��v����k�y-2
�@���w�h]_ZEg�W�?^�W,��{vo�[��ƞ/�k97��7���p1{v#�� �i������x��?ל�er=�Y���\�r��D0����{v�[7|���sL���~���W�&�^� $�ug?�H�~�ԩ#'O�|�H	Z�g�}�k�\�n�s�K�IJȓk�6�6��<����+ִ���ʭ�{�&- Il�EBD�(�śsxy�@\'$R�&
��XS=��[���%c�;�E��$��4p�������Z�s4���5OKp�x)��WAf��\��2��xM��n�̳�F�e�bU'�[�\n��Jql7�����J��S���KM`� �������b�����
Ԧs4�0�+�ױ�4̰�5�цʧ��yB���T��Rꞡs��Z�]���F�	9�Ζ\��*�m;���_^y��S?�MZ6 �[��(3�&ϼg��?98xdx��W��������tl��?�6ㇵ/�6^��
䓟�7T�������_O?�<as��o��0�#�>1<�'i��8y��a;(�6Rw����a�#wSK|	0�ld֒@E�!;q*�Xza���[���0{~�Da3uT���0��4Ѡ�z�T��A��r�m���f=���qHtf@J��:���������$o�>�Y�BD��W_�P;9���Cۜ(��}[��3��/���0|�;�a��°�mx��	��a�!ް�3_��D�l����w�f ���xSU
֍��\E)��P�p�bK��Rajy��i���h�0��|V��2"��*R{�4���u=K�E9�Vl$Ǡ p����{7ǟ4� ���@���gs0�V���-�#�jS�4�߫&+�����C������f�=�j�ltG^�TwW���N��:�:޺���&��#�+�z)�b�@)p�aq"�`�h�YQ^�L�t�\U��C��~§|��$��6�zj�@�D��b���F)�ܽ�����lX�:<��Z�!Z�x-"gM�1:u�-ڙ�;{8<�1rɮxa��K��O}���U��t�A:�8��ݘ�ٹ#��������I+��O�}�cOgE�)�Z��0���J��^�Y�r,���az�aRy��� +ih��VN/�I�h^,����"�3�ۻy�N�3
������R.D�,�V��Z�a��0y����}I�����uLM��ܼ%��dֹ�mEY��1��8�}��{�2���d*��e�I,/���?<>~/����1/�cv��"u'���x}w�;�H��l����*�1��o��2<��e�ȥ����+Ϧn �[�y��+��� ����1x�7 �D����Bk	��m�l�R��r�E޿�k�@�ior}[�������={@�~Э�
vD ڿy���ã�?>9�o�s��e�;�?�$u�0�!�o���۱��Or�7�_v���������!D:#rnu��AY��-AZ�^f��1�)VÖM�v1�i̼9�����q�(�~�K�n����7o�����H��F��9�3' *�t��E�V�` �9Ble{��n7���/��E~�����X�4<���ý�>8��|��&
�j{��U�SC��S^���U�rd?VɢUU3o�Jo�P}�k�ʍf��C,½W������(I!�et�Q)�2���kz�r�e-
�2����x�B�=L���R�֪�M}z����[Qyxe�Z���g��c���g�Lm�5�%H5��>+N�D%�3�-�]�'�v���-���G1W�M��y���0������.J�v#��,�������h֚����U�2�6�W���z�y�Y���*'� �`�H��{�6�� �(s�M3���t�#�~��0	6F#6��ѱ�TZ�N�Bރ���r��q���C��Ko��2|�3������9�L:�$2�f����8�n�o}�[��A�_^��X��(�<�z��E��z�*$�Hy�.P���Sh{�fO�AY� ]���p�����V��`^���������˽B=	�!X�B�)�E�P�T1�L&����k�
d��L�*2�AJ���O��|����P����+�����������p����ٓ�-x]��W����_{��h��H�^��vj���z�8��`	oE=��iȴo �6�N����}�;�^���8V˝�97��R�FTz��8�����\)1���P���z��P�2���%	ḗ6��Y�v�x���C��#��M���`���u�@z��!��/�K�,?F�$?�n��'?����o|*�Y��]��3��=���{`�]8�#Q���?(_���(��n&���YG�b���%X<#��#mL�5E��%������4�'�ӷY��>V���w_}���9|��?�`r�(�R Nӡk����
-�|����oE%h��,|��vh{�8�~#8B�{ȋ�ݵ���ѩ�T=l�0(^�����u1AM�}�e� ��جE���T�,'R����*hhS� Ī�-u{��+��27�?Rѝ~��ձ�J�E	������f3:����X~�?z�^#@iS�x�[���|��gYثƇ׬7��ZU���O'R5�an%�a�u	 �����5��,Է��������:�L��H����R�f$�Vz�f�^]s9�e|�,f�IZ���?P�>͞�c{B=�����i}G��|ט��|-)PC�R�{������O�����wŎi�@-6�5��/��c�� HSeas�%��H����s���N0<S�dY'���8F�E��]���q
���an��.��Օ�����X-ބ�0�W�2�c���7gABzq�&�{�����^�E�j��ўoʂ^^�:���K-��!��Mc���Z�|$H�\��t&,����Vw��b�1S�{���)B��Kt�EX1NE6��K՘(�H:�����A��n�@�w��+�Gu#I����w���g>���y��~���D���&����B�*u=����e�T�8C>d��K�'��	,L��j�R���o�)$���a77�|�O����#�d3�]�}�ʟ�ٟ������2��K���>����j�5潯���M���µkW�9���!�Y��h��2
A:;Pdy� ����Sǆ�}�Gx��0���W.۶n8����ǿ ��hޛ��q�TX.�H��C���D�G��Q�+��9��� ��f�Vk�Qҹ��%�#�b+�I;�ɰ%"�҅�Ʌˌ���ު�����t�z��qx��'� �w�J_n���ٽ{���{�)L��fTqæ��&hUJ��Ш�DK�Y:��Z+�כ��@���_<|�Q:f��JPy"����p�K6�_)��0�5���������%؉<p6o��%����׹���!�p�3KM0�
��k7:���5�P�i�,c��uվ�7)*����J*+8��Kz����M��S���oʥ���rhL�.�
/z�ɨ����tS����Ys��ʊJ��/��U������X���rn�^���Y9���m���6�/�sߛL��4 ����-��m�L�D�؍1���dL�/sź��E�i��%��sϾ0\C�ݼ��)t�f��p��W�N��N�_�6�z�v�ǲ�m�RT%8F��d1
@Z���N@�C��<��
*��+ ��Ʋ+�,s8�Fe��u��֠��{���oi-������ ���cK�e�s0;�U%r��Y~�c���wNʞ�/��]��>�$�,Z)jK7�����!��%d���B���=Zk!2� {��
�K}^��#�w��1�ع��!�	��M0�i[}�����M�]�=�֞3ɷek��\��yqL�k�֏{�1s6�X/��(=)����T�?�;~��� �.�^sk<�����k����o���5����4���8\<w6�Y9����lۼ5���#o����֛o�}�I�~^�Y��s���j���O��?pee��7��~w���ߢ3���e�jo�;O����ې�,P�n¾I�t㪍����B�>s�Fi$9��(@ْ���Y(ry��D) Tѐ��*V	N�>}��ik���9@�=utx���Y3c���q�rܟ��'ׇg�{
��/�u���}e�C��}򙆹w���ߑ������F@u�]GH�Ѓe����
Wp�X�~��D>V�,���V�.�=�V)o#h��ve�Asz�v��;.#���VO^!�R��5�*�ev���s�*�|��#Q���s.��7!	�\B�ݨ(@^u?sYW)��H��}����*��[C�;^�?`(;2�Ej�ZY�)����Zk`3�cٚ _SEa�[uh<�^y��̀Lz�jR_	���l�x����ｵcf+^4�b�T��x��Jw6E�j�)"�!��I���H���%�[M!��A����tu�PQ�p�P��"�_:2���@�ۺ��-�jkc�'�}FD�M4��Ϩ��1��硳�& )8�l�rΆn4�2#�P9�� +����f���N|�A�����Z����5�/����c�G��[�3*�l(�"�<�c�Q��Z��
�y���'y,ȐW@y�����}gq�x�89�5̃Z c��+��j�+�'�h9�E7u���&��J�S��&�R�\�B�?s��qΛ�H�
;a�e�c�Q<����rs�Q�H�����Q&��L��N���K����*��&L��#,j.���n�S;�l޼���թ����+y��dx���1<d�CQH�b�����!1c�I%`�E�X����N��B�C䌽��Z�������{÷��� ��_�,�:����_f>��O������n�Ќ.M��frFx&�	9�,L���I}�JV(����*:�.c`w��>;�I[����E*�;
�G�`6`�,Q
D=8�w��i �����[a�ӈڈ�mH��Gxax�����H�M$������/h�r����ch�K���q��hﺧ�ʹ��;�M���C���<����:aޏ�ջ'T/7�)�
o��,�z��)k��O/��V�r÷���8���{��&/95�A����;��W�t�[�=|K#Ğp,�2�3�E�����lޏ�װ(��I2����$q,�0��≶��;��퐳�Vz6{�sf})�HU�Q��i�����;VT�)���zV�r_�m�5�|�xД{��\�9Y�;�-��5�qͦ����;�&]͘�Ik��X;wFO=��:	5��Ҡ��3���m���b�)\	���II�������|������#�.qx,��{`��B�����KȆ;����:�mP�=�ܬج�Z�k��B(�4���\f���i�g�i1Sn3��>�^�z@tn<��aF�{Nar���u�.��/ٸAʰW+'gs�F��1&��C�TaC�n�p6:��3.���L���~�B�s�Bh�ܪD1��$O�aC�J*f���Sm�״���	N�����`�������-'H�h�H�Q��ڴe;�Q6䖝��\;6�d�����9�$'���(�|����"d��$5�����e<���Y���s�s�����}������ӄ�(���tnnx��W	�����?��&�.ԯ��?~ix�w�	O������ �J�|�`��!�|��������ȼ�2������o/F�Eh���	<ѷQ���|���a?!�'{hx	p޷��x���x}�k_^��������!�g�PP_�i/TJD�lx��Ѵ��A��<(�D�<���f7�Z�y�҄U�;�����`>�z���+�0?����kg0�v ,���޿�����-�?Ex��a=�7o�J�����׿}lx��3����IJ��1���t#��2|��-��CJv� �{�!j��ʺ����l�z/�*0��.�i��h^���+҄�y�g]���\F��>�e*]�����U�w�v���qy��m��=�����_���0��ɽ��!��iŔX��*�g�L�I�|T�:��ngDo��*��,���cO(7LA ����L�-����
�7���2�43Ҡa�do5�X9���*>����.��1�#�w*�����c�Δ�
���(��(y�x�S�����u#/�H���;1u'�U@�6ne,6���}̋��$goy���D�\"�IO{֛�8�K:v1�����l	`�[C�����0;�%%��|N���VB���q
n#�"|�ee��T��s��n�o�4N��}�(,d�BA��B��7�?�gΖ�h���.��$Jgލi�**�S�;fH>��*QQI���JS����W�6�һ�s�� �;6Ӱ�~��� ��t�O�}�� ��S���5"B���{��d�����e1�6�/�{9�
T�?���҇��`Y����G���I8�}(˴���]�	y]�4����6}Y���~��5R��y�gZ�][�O�gi7��I�5��e����zp���'O�<�}��D�~�� ~aN����hs�h|��:��y����W>�	�{�ϟ~*|��P��C�z�_Ʃo~����3�������׿J��j��×�u�t���OS�n��[i�"���+��'ՠ�oC��v#\�n�����*S�V��a)�F%oEr;�i11ů��j���[i�J
��U�C����p��4�/,��8�>>ǜ\w�P<��~�3��=BNCQ��&�o��:q����/_^{��1;���'>9L������<|���&�����;��u\
�E#��ඡ
�B�F}k��؁m	Is/��C�*����[Ei刏B�WT*Qb�%f�h�4��Ϻ���<Vg��A��s>��5�G��{�}��lͻMN8�2؋;��ι~�f� 4��g�P�h��K>W��*(�t���7i�Sv��M��F���N�<Vs��f�M۽.�ȋ�߲���@v]���`��C���QR^�X������|�S䵷��x�Ց��YS���4�@�f�HsD�^y�d�-�����L�����h�w�>�޿�)xD�� Yv�ȡ#�,)7���J�-r0k���N��4沝��TJ�7��!c1ޗX��Ww�_�<�͔*�*K��E�%����OV�ц��#
�l#��� T�#��ɔ�n�H+(���n�e.�+������ G�T
� @1dS)�)������>���r��/ek���@����sj&o���j��-/�+��f(�Rи`��=�^�S�1�W��|��7J�f����8�T�#$~�6���D� ��qi�� �&����l�#�����(#�
^�)MKhl�1��!���o=;\#ל|j�w�xyç8fRֹ��'G�k�]X�[�>�uj6�ܰs���O>1|	������?��!���DAI�aLۗ�/������~��p󔶐���&�ٳ{/����>7�_��=�Cy	P�b�����q��˛f���n<���&�vָ���;����Nb�RY�~�#@��2r��a����G�R��'��/��
Į\h~FzW��G#'Dl4H+�A8rÖ|r�6S9����OcpyXtDS�x5���g]v���9�{�$nM�.��⇯s�*�'�)��uHe�Q�{��k��U1XX��x<ɋ�'#�(J�r��i.�[\��*$^{�{�U;^��]ڌ|:mu�m�T5D�S�֍Võ�=��yG�w��=���=g��yM#eP=T_)����~-Ui*K�vUBW�#?����9�ԭY0 �{����M���B/���D�zrƽ����7*��������7e��bP�0�qf���B�B�!�,-á��4���Lc�-��C�	\
�<4�����}��
��K�c���apY�D�^���w��Y�^m>36�9u�ʹ?~�RFJqSx��o"%6�!2������;����f��~�s7Zk[�j���4�,���8F�7:v'�/Ys��8]@JyS��<�Q�,H�ۿ�\����YңY���&r�	����#
���|�£�}��*��*@DJk!ZRȤd,Q�*�����"�'}�4MHT�+��ޒ�Mo�����: �;Գ��%0Ap����m�o���g|���BWc�R2r��?�5����ʖ�J��F�)ޣ���Ux<�8�G˻��}
�Ǉ�߆}o��"�ۻq���?5��'p��/��^y�h��\Ǥ��`� g-����5������_�M��p��O<����3/����3̓�Dy�dӪ8=���'?	(�������?��H4�x!`$n��/|���D��=��*_�	M��pFs����/�a����K0I���W^O��M;Q�S}���g��k�` vC�b�{�3�=��%��5� 4Ȱ}b|��]���r�c^���KYPи�`�\��B�"@� �m���z��.5c���??{��̰�0u�m��EVKM��FoX� ��
^�x�唧}�49������%l�;%�$��t"p�Kaj����Z�5�Df�hzs�����uݮ庽�^:V��jD�y��1���d�,�����X�ʯW��iT�=z�Q�1�/e_���纛U ]k�2���y}�d��yN��x�8˒�P޾{@�Jq4vY�8fW��j'�˪E��;x]���^?+���U��)�f@���Hd�7�(wٝ��3��������1��ˤ����CN�〔�km��,RW�� ���k 8�,�vd�:��r�W�4�#����W��)�$���� �F�ڏa�)p3�8V�6�x�-	p<��`F6���#ֲ�&��r�0rk¹���|�Q
�M��G?��,V�����V������hÅ���L�^,P�`��[���e�*`��L�Yeq��ꐕ\Yl=�[�7�Z>���d��]�]�v��+��9W����dfj��Ά�����+^�m���zhOm����%�o���{Q�����E�{}��a��yJƮ\�?4�`�l��U W�k*48�V:��M\������������_�2�.e���M	́X�n[�n׻+����<C�nF1S p;������O}�zqx���	�/��~����ç7a�+ઑ��6 d�]�0���!ex� �Js������n���3���dO����I��v��4���/����{��<���O�����!B�[	G?��G�9Q�O���[���7Ŕ/I��Z�f�J@ #Q[��Py�bD��۴�
bY0d��.g]��׻��-�}���[�����rO�5{�G��q�r�p��Aal��M�T�N�e2!�Jr$�IL�z�0�����9TZ�,��d�3��V�(�W!������cG��1c�q��{di�3����{޻ל�ptO�i���,t]9�Z �|נ͌T()��{�}?�Q�v���[}��GB���u��~n��̬ܽ^2�o�T;��%ru�a���e��5I���ܱ�h5*B�f�ٟ��ȇ82��Onwɓ�1e�t�\T�)�j���N(as{k�ȫ�p�}�O��g��_��p>�����0$V����0��j!{�X�l������ѵ4��l�Ȳ4���D���HS~��|��oڴ%�OβOg!O�M��F�w�$ߟ+.���H6���c���W�PɞCc�CcD�����������O6�8���LW�[��^��Rh%>|��|�Mn��6�����,�Iȭ�a�V*2�t��j�$����vd��^�Ql��h���]K'�ڣ�G�l����YU�����{n��[��p:d��*^Zh�����ߞ�����Kn�����S�~�l,�m�9�P6���L�?�ϦәD�o �d*ہ}��Ki�x/dQ(\��>K����DT�D��C�x'�5������}L�j?I����?�]� ��A�g�9��w�����Hd��2�Ԡ���2˲L�m��ݽ�����y>��!����!����r6�������N����	�x�)�H8�p�e괏2{���� h��Ƒ������0 'FJ�4R!�ܭ�w�a|(f�"^$�0K� [)�R���R%�#�L�b�p�"Q�׋���K/?p���y-��R�o+�����m�bZ~ @rT�����@�8;3I���x��`/��s�ɿ�]V�)�*]�4Ft����,&�b/C�{��Z+=��7Z�֑𣯅��s5�|������Y�^��D� �w�=�<�����n���8J��TB�_3Ҙ�nxS@�K�A� U[ Mf�H��	1)�,�P���c��M���W��F�E�P��H�e��oFs�[i�9�U�ՅLˑGV4i��r%���#�6�tM���/�f
f��4ڀ@i���_�Ѽ-�YZ��(�#d{��B`��d7�S��b��j�{��H�á|-�/FZ��rz��=�E�;���ߊ�p�Tur���HlAm).����;�q�y���>��F(�� d�<�nE�NK�Fk
=��'Xko���,e*r�Z�m��"����Je�w�����nm�x��{��L��4�&a��ΑQ�k+�_ @���,���r��3�	>�X��pC�Z�uWX~U���إ���W��A���,��a@��S�w~�\��q+=�������:!Ϋ�$b�Bmۻm�����@���8�>��SO��ng�(y�8\#�o�7g��T���WX��l�}Ζ��_&��kJ�1P�\�����F\��:(d�%�sM����kxBzG��������S����y3s��~���(�z�P3�5��o�Σ�o��������}�5�(p�+c�o bq�<HN��T��z	��e+FK�֣c3߆��θ����'�u�R�f*E�*ذs��fH"T��д�sK���V��9Zs�\]�^IB�K���~���Хh4����6���y-�N��A�G��h�7BT@�y��M�����4���AџV�Tŉж�ӛ�Q�Q��k�k͌���1��Z��w�(���W��AM��y���8V3 z���1G[�f�DqW� �y���M��g��k-������F/4g!�Z�q>}R���k��M��Wࠨ5]�-ͷ��w�D��0���.ӡL�Vg�B���n3���7۾�d�h�G�zW_�]�-i����/� ����\�e�bD& �MY�H٫&�F��^�c4�{�5�J���
H����JX�q�$�XL�F�ăhlIh�ꭽ���h�w�c�|�F����E1�n�W�IVI���r�<�����Չ�kz�g���V7�/
�5�*�qU�>��,!Q�����^���Œ1�����`��Z(�V�1�b/AW®tp=W�������P�7���W��v�,�n`�����u,Z�)�j:Q- �����t*�z�y�no=Y���V��B�668J�J�{�@�������yrŷ�w_��8�y�°o�V:��;��ß�8<���Æ7OR�}a�"%G���)��_*��AUT����#���$
}o�uq��+U`��{�@]7\N�8�1� _$��"����OϿ���6%p�xG���A=w��}-/��a��}���[�>�n�I����c������tx���4*Am��K)����t�7�����P��I�?׭"R΁�`v��׬���鑴2���/��EDs��R�ոEF�.&#9l��\i?��2f��1�k[�>l|�w3�o(�+����uޤ�d�&>��P�e���I��+ݨ�2��~p-��Y�]�n��+�5"�bZS���^6���Bm�*��Z	Z��U%�k�r׵_k�:�=��=�C��T����f;_|��xӉ��q�v���ȃc#;�	�(1XP�6x
q����T����T4��4X3n倗��tq��p٠�0<'0(g)oF���07Q_,�.=�U�s��}�Q
�	��t%�Y�s�*W#FP`䏴ՙS�42=V���-{~ɴ8�k����B�iRVz��z�[Eb�A��A���:���=̽	Pv���#�|��F�4b%��m��Z']�_K\�y�`D{|h�?�(�A�p�¾����J(����U�וe�hZ��nĳrsIo�7ls�ڂo�0�$��)�ڐz�E=�����WBYmA7�]�YRH��R^��C	��
p0�FEF���]`}������k��[j9��W��(󤫛�}��ckxK.z:��:�����@�z�Y�c+����sP���?�~�F��oP�{�wO>CD�<@:��#/��e�Ǵ>{^�u��A�H�R� �����0� o) ���,�FF>��:���0�K���5�}�.���s熟��-j��&m
��G �|����<|�;?޿���H�Ǭ~�����=�������䖆{���w�O;^|��A�+x���kdJ77mH���?=&<�m[��Iى�fl���&c�1��1�N���"�+ox����ɡkTVT`TL9�1�;���?;�ri5�ˋ����ֻ �_���3�o��ǳY�q'� $/ꞱQ�� Qj�uv�F� Mq����*5�5sՌq��c�� ��"���hSކB�Zc\b��y�M�3�Fo�(��騇������
�P]Ft�A��!:�Nb@��0���Q����+�����;�-�v�n��D&�b���c��x�7C|A�8&_�+�w��Cw-��߰�ְ�>�Da�k��_����4P_Uy����پ�+B�oZ�����^���Li��Lo�����,)Q���5b�'"7��E�卶r��br�_^_�����`.�!�S��9"Fc7���q�xЩ[̚:+���~��>��Z�B(��p�{`���b�]�eQ�ps����7�0OSB����S�mPJ�0su�*v-�n~�o�^NS sh"V�����r���{�̬��u��� X��skzkB�E.?`x���t+h�ս�
�l6�OE_���"�"�ۜ& -B�Q�[�Hoī=��Y��}��n�(y��7m�3����xi[���<���e����O�1?�Gw3�����Z�|h����.���Ru��H���X ?���K#�5!9м{{A�O�5�U��_���8����u�S���L8X�vmx���C�������ej�	0�a���?����6P�/Ѧu�?.�6���\�"s�l�P���Њ�6C}���č�6�g	�������3���-��F.HJ�m���0��1�.F�9H6�$�qb�R�i%�rM�#��՚�
&�chi^>��'�o|����֤o�y���i>��/�)8;�ɀ��P*x���۸k�(@r����ֱ�6m�B�:NK�-�=�qK"T
�x�}�y�zkͰ� r�}��>|�{�#K� �H�댏�.�{J�����Z7��
�%OAH��7��4�Ka��]�F��89^�	�3u ��7;��*�����t�6c��~�Ţ��;*_L�I�k?t+;D�+�4		Us���m0�h)m��&�`�J�d>8����������jAJE�`i�(j�O�)�N"�H���QĒ��{�7I�#(8�)�fd�as��%��TZ�����d&z�r�#������NOɵ:w��|2�Ӹ�Us��>�{����WW{��O��L�И�p�g"7ȡ��|Y�|�?�(�����w�^"jջ�/緹��[ُu5����ݤW4�PS�<�G4k:�Cڦ�=�Z�������
ǜ3j����\�.μ��)�%�)��P��(a��H7k�r��ꑚ;�L��c4De�ɱ)��y6E��|�k6�(�M�ӕ�L�	*��5�?��φ�|���w�X�tk�p+�q�\�o�{.�BnY�eYS�WDK�D������M �I�Ys=A�BW_+p� Ebz]9�-�f���Ǜ�J������Gh��5J�"��-j�W(��K�O~��c�.��[�(6����O=>��Ɖ�,�>�����̟��O鋾}x�����)5���Jr�Ǉ�jr� t��Y�7����	P��'{;�B��Ĺ���>�ܳe�����C�+��0�<vt8~��a���^hi�E�zvM��0L�p����*ty-�ZE*�Z����a��-D6q����箜N�x{�|��a0�-���D��wu��ؽ�S�ڷ��),q:Hv`c��Xi܆11{U�^(n��
/ 0=��ᦜ�k�M'O�L8W�R?}�T�M���|����Qڮ�"g�x���?�I¿<� ��s���pp�sϽ�0�QR�wD�믿��nݺ5���h�����p׍�k�-�U^�7kY3�{DN�g����O^���T��Y'��������"�Y�� �hr!	�+7�\���HY�8?��ui,�=����x�T�Ƅ�[E��v[��M
%
���,�&�j�c���\����Z�m��d��;!��u�[sN�������v��s=�o���r9�F����>����Ez�;f��I��m���3��Q
���|�H���,�&��̳��k륈*�X��QE�A���&˛��訁�5�o�x,�ֳǩ�#[Z����@��D��l)甴�+�yچݕw��&�=J�" �P��®m�{�N�مO�x����:
$Ta6�iE<ե���+KL����
�1��S'aJ{B��@����!��ߦVy�ҩ�F���ѐ�������oa��ڼ�w<��m�D��eYz���+�tF�ڔ��x�.02R��x�O�����&�G��Y����EǾx��o���J6��Ǐ'�y;���ԑ�0����dmMM6".�;��WQ
;BV��<>|鳟`�@��]B��޻cx�8�;ߝ���mU7��^�u�R����������D�.s=�9���Y�k����3?�i���=�P�׸S�����u=/��Y�H#fC�����g�n�Y_}��ч�J�s�>.�՞=}�����X�>��0	(K�ۀ CzR	��^	Zy�6�֡����8�d���]�az3�t�Wٛz�-�j��������E'q�w_�;��RN�V�c��2��u�.�s�N��e<�t��[W�
���n��C䣑,�׈R�������th$��)�s��w����5Ǣ����n�d�k�l@�[����u/�YN�c���4~3d�|�HP�5.sa�,ƹ8�>k]<	 ��q)��7O���NP`�]=ٙ��ФB�M;.Q_,1��;�b.|�9?A���E�u׉�ۗ�"or+_-�#"
����7�y���m5�E�y�R�	�s}�ō:Ǣ7���������)�ߌ������b�{u�yO���f[�G�G�"-�̄�*�R�]��?����-�PqLJ�E����b�sk�6�w�m�,��!G��hf@��E�x��He����;�vi�֕z��=G��5�ۯ�[�]��r�CzG���a{ CQ%ږ��Q��Lo�7���K����X�1�l3��%0v	$���[ J9t�p��֣L�ʑ���OT@a��nº��Z�56�w6�f��κ	n�v���@�V��!�P��[rd�:щ2F�'ᮢ������w߻��Z��G��v#H�3����G�G!��Ƌ�H��g��0Ϟ� �qc(�O|�I��_�X>9���?�yܲ}3����ȁ�a��㞓���4�x�����&�������{�� ~/�~�\�|��utػ�� �u\�E:D]&Up2i4���WV���R���\��7�.�����v@ͻ�Qy�'1�0��>gc!C�*o@�!�HJ�K���>�������d
L�������7m��22�,
}�*VE �U��M	(ح��*^��h�}MaV�qC�O<N��S�վ\�ߋ�+u�`|��ƙ���>�����;�9k������a������~�ϩ�ϝ;/^%�7B��o�K�����k�Nq�`bTX#Fzɯ
�&K:um셖W~X+}�y�?¸��`r�(�h=�uܖz�*6Z��rH4,��hY��)��')#[G�xU��O(����4�m�j�lU�d�w@/����xOw��b����u�8e#�F<����\~�Y��^��R�e�{���:_��r\?�f�7���@7�˾�~P���b�5���<��&�1E�%F�-Ѣy҇F��N~~�(t��A�����C�`o�23�_)��������-?�-�t:`�OdϗE6�A�BUڝ9�+��~o7���X�t����[�\�fh��.��j�����G<u�Ӆ[`Q����Y�e�S롗�\��uޢ���cu���R��R3�M��X�����*����ϧ����3�����n�ӛPN*_r�7�H'�/me��3wo�ܚQ���ث"���|<����]E*T�=ק������X�Ȉ�9k�y���G?�E��c�ޖ������5��o|�f-W��	?h���O<pװ�<�>j�=������H�����?HJ`#B�����	Ť�FB̀t4��[]�rz�z��p���BV�-_���	�TLw�&�?	�����j�f1n��矘Vi ��^�0!Wю	<�� �륺E`	��)��P�\���(����]����"`@�W`�KȚs^����>7��?�ï�G�,v�����l
������k�,4�[�(�+b#%l�W��j9ZX!N�x��jM�h��o��/�˽���z<�*����D>����Hw��um�u�}���������<J��~뷆�{��5���=�\�̿�G�1u�Y;eT9^�D7N>�[h�Q�牆Q��׈�l"Jt��=7���`+��HMzz�&%ʙ�����^ެ�짢�6���\��S>_sQ?��R������
sת)'c$"�h�^�~�sJ�Ǹ���_���Q�5e��i9������`oND��k=W��{.>��J���%�<��C:��l�Į���Y��O#���1��"w�BG�����K��e�,�n�L�h�Η����N9�A����hH��7y�7�z<�B����⡶ܕ�7���zۅ�A@?_)��L��(�����{��|�Ub���J�F[s�6�\�޽{�ε��9(�N�2�GE�G�ExՄ�IU�Q����O�a�!�^��׭ �Q"�c4���h�U[�҈}�r��hQ��]�|Kr���n��j��X���P(�Z�ʖ�©zo��?IL�f3���ն��ݸe����?�~��p��{���vv�P��Aj���u�	�k�b��رe��8m��:���Ƭ�׳J>Snup�[�D`vflطs˰o�f������O%�`��+���a��)��
�NB�I�����@t@�#�m�r0�bL_d� B=|�
�4�m\�ᚖ���5ap�5||��}ۇ9ش�	�?��/�0�{�]�wP���p����UfZ�Mo�l��1�!����o�*8�C�Ғ��ٸ=�n���es�0r��b��5o2
Y��t�o��o���
炈�n�t�rޖ͙G7'���`���o��o�*ٵ���?�����?�T�a~=��Q0:0���[��%T�;����[��U �*���v(c:���%�l��:t0-|Oѫ�ƕ����$�U��dHV�.���&{]㹸�E��{"�R�떉h�����1�k��g\h�)�M��7W���9+�E�O��<R�˿Tx�^_�)c�>��wߥ��,�Q��-]�ܑ�^@l�܂����¹T�K�Vi��{�E��ږ��MD�<�x���8r�k�q'>�c:��Bbw��)������n�(,חs3��Qd���@�6!��(�f�^���	�7?� 5��\�:���u�fH�FF7��*�\�n�[��d� l�Xs�������������C�>	���m�;�+�*���Ϝ�w�guғ�vh�T
���~���'A�ޤ�ZZ��Dy߲Fk�l�[xL�+�&���8����ǌ���� ��:V(��,���Av^��f��{�}��-�#J��-��*��E���ί�Xfvf?Cx{nx��w��(�x��C4��v� �
����1_�{�-+�w��&*s�#`��K���]��jt��� �e
C��m�Ƕ��nڻ~�Ệ};T���/P����7��4���)_�F���(X��߂���D1�W���q|�!bDJ�_&��2O�h�Gț������͖?��<�;��&"�v;�A�s�P�����l���l���VCv��102�����4
�̈��s_ۣ�tv6�{�n�s��\� @��5�mKW���p(%��8M�َk�4��w�}�N���[���{�{«�?
�Ν;#+zw8C�K���.�F�Y��?���i,}0��(^ߟ=��>
(�s�1�F�~��50T����A������ʐ���"/·�S��(c���Y��g��M��ɦu�T�>�3�7���,�ri^w*���_��x�m�� *bX��jV5Wt_�۔��ټ�;4����=(��d<�eqe�z]��G�s��_E���˟�RZ�c��M��P��j�@��k���+�j<��C����Z�����(�UWmu�nҮ�no
��z�j�`S�0����o�Q��?������=?߅A���[�Џ;*$Fa?F7t��)4քb	I��
�E��+]"�4���l�?�Nݻc�p�&%�+�l����T��p��p���6Qص}�p� yG6�['N��C#�'�v��ݥid�5�= �>K�Q;��Ү�iK���3�"n�f��m⡇ڻ���Y�	��Q,�9E���H
�����?����fw�!�p}8rx�p�й�����I�[��u<C��i��ѷ	S_B�V7�!���Z�	[5� �	�z߈
��K�9�V�o-O�s`����y�Y�֍�$>S(���w�������h�s�:Áh�ٍJ�gO=;����*�-n���]KNr{~8�o�h�V)����R���hN�q;Ƚ�o��<h#�P^�B5C[�M ����nb45�Ԓ�7H��A�T��9�Q���}�����]�T�ɏ�Z��5:�#���jѺ����U�7h���p��)�	|=��6�ƹ��5Q�ʖ.�R��?y������G��tע�9j�e�uv��0j�����Q��R�DalK@��t������������.>�{�	�d�e��l���c�(?J;K��Yq�s ^���2�Q���V�S��R§-1*ڢ-����P��{��Q���ɾ̚)o=�ʳ22Jn�����7�F>;5yss�`}֑4NZ$4��KK��~�:��FD����M5�e�o��T	P�:��:���Awd��Nnl�P[J�>(����f��bM�M�׶�*���2эW�j�u�}5��2J�t��c�V3 |>z]=?���2����qG��hnԋ��O������W���%D���
�`������,ex��������J���ײ�������˿���w~���� l2=��~{��o=�]���KU8��Q��Vm��Sl"Ѹ�2���u�g��R�+�2�e�!lJ$�$}Y�e�7��&2j]��O�y��̰�u�R�g^<6������ �]'�2���a���U�<l#��H�۳-�����7#`,����\C��S�fl���5���MYP�w�OOu���Mݲ�ĺ�nnӖ���
���;��T��47L��4|����7�7�^�N?:��ҋ��I`��q�,:���j�eв���MflU�����O~�>��)�C�.���#�:Rh�_>���s����Q��_��Gk/vƶ5�u��{4rE��NCjd(մA�����d4�N�@�����U������|���'w�a�
�P{7��LH9*�ei��h��}ͰY��O9��%� jE�a�8���=4$� S��S�yLgC޳\O<O��k}���>c?a�1*T���S�ҫ=��R��3|:֞K�����q�K�b��V$A���K��h��8$�d�ƃ����g���Ջ�,2^��@DO��i
��Ƚ��R��d���ߺ��z��0Y��qݻ/m���w��_���;��W)��_����C���L�R�n�[�]Q�z��F��׭ U���J_�i7\�!�������������z��������]P�U!�l��F=�n��ޛ�x�_�����֊h�f����7���~�f&o�?�c�y-�pѐ-�mt�?�����������~틠�g��{�G�Y��K��rnzۅl����zЅ���0�n�Ox�����"5TQ؊��n	�dZ[}V��۱j�Z���;Ǉ�����S�%�?��q������B/G�F�eI�U��%� ��s~��ru���DX�&�]�(��0Sy�#��m��=ÉS硚}���	�n�p��$��Mx�� eYi]���ؘ����ר�>2|ꓟv��7��޻��edx-���]x�@�Mn�h��ER"0��ّm��i<�bP�%|�s��\�
�����Djv��5|�����/��] �9�� �u�q�GgyT�}�;U�s{29��k�㬳.���`8�!�3\Iʱn5jԍ����L�ݣG�����T�e�B[�6���~�%�Ͼ՛cz�/[�4O�����p��<��0���v�}o�W4|������0o�1�u�U�ݵl��q��y܃g��Z�Y������:|	x��c���V�o��&T��S�T��Ζ�aٮ�ͫ0�t��7��=g՘e~,]c���2p�|��j��viʚ�&8���2��`+�:��o8�(\��/�<ɽQ����i;;��v�Yw��W�{*X�`�}1@[YH�K�z�,�K���[E�D6�aKl/�7�Ք��z�j��D��|���FI�T.#�&'�n2oW�����
<�+}�����66��h����G�ص!��e�<i�[ϑu��n���\{x������u�н�Qo9ۢy>�!����u�r4��?߿�?3������y,�;���>:< %�|��ָ��7!��I��Y��4�_��}cQ+�(�ϧ��A��A������g��9rǗL�aL37E�^gдQ��Jd�t��x[n{�h�Bj��#X�Ӷ��筀!�܎������/\{�rϗ�^@#��]���G}����3x��gO��6d=9��1�vQ��q�x* .]�Fkǭ4����>���G���0 �zr���_��_�{�[���l��ȯ�n}�|������5v���/V.#�P�x��	��^v/�)*�)��~�4��8�,\ ��ֽ���wx�����Fʤ7�x	e!�(z5�Rd"�-{��-����������`�_g�N�-0��ݲ�~LĲ���!�[�W��<�����YC�b2�77��R��&J$X�2���Ͼg�am:]7���={�D�-A'|��6JU�7��{s�/��O~�c<����U����Z�����h�L���{��dS�9��FJ�D�[�nOo�/�6��r*[\g(m���c�ZY���!�j!�!S�1�A �Mz!\��L4a� ����.���>֣t�`���q��8�[�}�S�(�µ�b�����W���0�;%�ڸ�fƎ%о��{>y���{��'�
�b��$B#Xͮj��=�W�N��p2��T�{D'}��g�y^)��}L�J0j�Q�u�C�lE�-n�*��s�Z(�K#V`�b�/I��O�$`\��K81���nxY����e���W�%�u}G(tۦ�����)i(�`X�G�3d���p��mH�q#�k�)��q-��J��(b�U�������!�
�U\�{��~��*Pםm�wME�4�+��Χ�{�l4"0���itO��u�~?�u�
y�g��� �����4j��};�6kmA_o$7ڕg��k1�/�?��	�mg�Y�0�-<�}j|K�Wc�r��k�f-��u衏�ٞ��Q-�^��R.����̡�b�\}B+k�}��gs'���_p�J~Ae�W�P��Ye4~�^J����C�!���}N�7���� l*���ܗ�����-�6�x�
����ϜZ�z�9x�Y��?��? Ran�B�Ρ��x������K/��f	O��h�������3燧�r��q�|v�ҳI�#Nuy��I;�N�7}��(=t�$����~�l����r� �T��������0�M&�z��^"Mq�:w��BC�Ϟk7H����W]ʲB1T���	o��.���7��K/z~~nx���
{۶�	���1�~5��~����)s٘��U�~�*ts�c�4��E�\�.�B_�1�s������J���eª��F�Ч�;ʯ[�GTN����P�>������˯�!��ڸ��&���	/���L�A�u�^5�S�1S"��+G��[�i�Ҕ��<v6I�t��������c�����Ki�깍�X��PІ���(t�m�l�����95�7p�(e��C0C�IbR�s�wf�C����vu�u&#�^�F��Zf�<��g�o९g�\.3f�Sx�IePwʫ��
�
<�����9~���ϟߨ��W)�:�5�����ە�h.�a}�?�P�h���g�
�!��P>k;��Yx�y�	�y"�JД ����Q�|�����Vs~�/��[YJ�H4zz�$��$f1̥�+�3��Ր���n����.��n۾u�qe���Lʦ�)�m�"�6�%��%��"�eU�G��_�R�.4�35�\�p3筷" ���3�
���}��/������o�XZێ}��׋�d�#�!
>���.<�i`�1�۟ky�8�xN�t��7��<��ؐǈx��L�2�L�����U�����+�Ϝ{�p�L�4�
${���\�vO�R�#=����÷����ЃSQd��W�-�ҵE�f��\�K 	�- )>���&A-"#�8��+ MF��\��@�� fn��	x���o�8;��{�~�Y�^ZAK�ת�|�y�-��x�`=e\���Py�Z�G�X"(F��[��]�"���{4*�\��[�p�H�ji�� �����0���zr����o{I"���/�"�z��1 F���{�ˈ9���fa�#���:���>j�/�e^r��ި��� S�f]C��a_u����7��ؓT�\�L�����:�'��� �Z�U΁�[G�r��|U Ďu�TY+�3U��s����cgiժw��hߖS�G҂��F?���-Nf�m`G�Kl���<N�b�A��9��t׺ڻ�tuH�0<�o��P��x6*bT�e��F@����i~��կ�Ɨ�O��S`}ڍ��w�9� Cy4¨H�6.cD�n�4RH4��'Bb�"�X�������kyF]������:g�'���M-� "W��kn�
�S��H��g�w䆫�N)뎦�������9�������tEdv)�B��
ܩE�r)~�gz�����[5� �'B�m��=7���ٗ�W���|��# �����h���$U�;���c��8�Y�Gp�q?�!j�F��"F�X��n����-� ��Ƚ%�g�K��X	���E���6kg����S�4%�ؑG^���N/�OaE�M�VC�K��ϡlqu�Z!��,
\����4�Y���5�w�|���뷇̈́z�Onx ��ÃG?��χ��.��we��{_��'���C����e^�c�Bs��q��<�Y�C��Q%f8���&Ü+�k��p���$��s�
��̪���5�m����Fhĺ����FV��S��UE&�󺥝���Z�Q�%�/Ɣ���\r���4���6"J{U���1b�=��=�M[*Iic�y�2�z�E�\���ź��H?��b>�A��^�ىiV�U�K�m8����#G���q���s�o�k��~�����);���� ���AJwV`�MZ����1p?��G�@gv#@8A_l������@E��-�@�#b�ޔ�:+ݬ�D۲t�����{8���$R���/%��������n8�u:+J�s�Ȝ���r�*��0 p2�eK_�A�ԛ�"��DO\���s���%�$g2u���Έ�ն8�~��ᕗ^.\<Gl��я�����9�{y��+�n!@f>eD,?�#��A��PC����x�:��>�;Fi�y�,��iQx�uZ+)�BGi���&,�x�=��Ӈ�o����[�a����5�[m�(�4�(��[��t/�pV	ʘ~��F" �e�5���g~�_�j��ЮA���m�K�ݕ7%p��z_��X��{/Jo'!M�va�i�B���h��W��f�d���
�*�� �s�P�5끱�R>R@!ˢ�VƉ�R��z���������1>ڕ��X�e�!AS���>�я �"׆!���/j#���u�� ��x���ُ>B,<�y��:Ы[��	ᎍBlbry8t׮᭷^O>w�P�ۇ�ss���9̢h�y���"�˒�,"X��?@�pWB��6�nϽ���U_{�V���r꺩B�u�R��88o奲��b�s�r5*`O���4� ���jc�w�][�s�<���Lx梢XkzA漛Kx^(��2iq*𫕒i����(�n
��"�[��*�[��]!�G��M[�q\]�=�$��6ڞHڠ�ٟ�Ǽ�N �T9�� _Ŝ8$����a��k1*/{$��w��.��[5�c,U4n��&��c���Ű9���b���H�l�Yˆ�3�w��1�sx���a����ṗ_.B�,�KQQ����h�u���������2����pP�e��[���#��]�"E,
r�����3��.^=���f�y�sMkh] �r	�}9�O�:�{�N4`�u`EMR��e���s	�s��ft�"N�k�6���d��w��sx�q����k��Q���X C�n���އy�%�o9�Ir+����" J�s�$���#��#��s6֮��>��? ț ��Qm�+�nߊ����mu�eE�T�������2�f'kg���s�)��ZM�T{�s=�f����f��hRX9���w�C/�G�lZ]l_���`�z��)���]��N�"̇Ww��S�}�P��m8�Ojbϱ)i\!��_i��uz$��m�w�Ǻ�j_� ��|Z���Sc�T��<�֌"�o�aT`¹*C,�临s�2T�;9~�A�y��(���T��76�g�n����<;<	����=4D�~d?�����˶m;#��1_����������7�7���ςt�}��hn��j��n�lټ�\9�0xЏ?~������6�˞@���`��W�ܕ2�J�Nzz']�ҧ�J,�r��kߑq��Z�QGO $�)�Є⽄���4ү<���j�-�g��|`��S�	��.n�ǐmt=KD����mD2����������2�cIQz4�\�%��'/\Q��T?O��O��ؕc�p���MŰm��TYx�}Ҵ�����/�@�6�`�Ɯ�4�*c1'��� �^P�*}���R|�׹�{w����~ޭ��HKk�RX������z�}��5xMFcV?��3�e�]!�}��9s������!R7FgX��bd�}����P����#=�Q�PK�V�T帷���I�"j�G���������0�)��m�bӤ�Rk������笖G�B�e1��+�רܸ|�"J�<ǆ����({@��V�H*�5���U�P,eX j��Y���,��")�i�?�#�����"7xq+�RX6:�����Snq?D��%��kb�Zl��N�uG(�3g�<�BO���+�����z�iS��6⡛�r+&�Y��*�X��+���9�icu!��fߕ�6��c���s���Lj#զ�{���;�4��{�B�!�<��z��Mx�?J3���B���`���Xʆ�@�^Z��� ��g7lb���>	��1Pۻ��n�]-����t�76�̆1:�m�x�}V�8%<����j��eNeP��7� ��5�F7�F��品)��Q݋��Nݓ�ס@�GP?���^Ν;3�w�����'N�&���]Ò�I�Ɵ}����[��O�n���$�~�zB����p��"����'��>|/��pE�;}�8��ΟG��$��j��'������������"�ERQZ��Ly��1�w*ʤ'cX���
zh�y^��}��s2��642.
�r������n��H�R�Q�#�L  ׬�_On}3�Ķm;�Ӕ�A�*P�9ī#^ߖWh���:sN���(`�����|��.i��uDy!�ס�r�
��`���a��O�� ���} �>ɹn���3�=֌Q�������W^ɱ��և�MYT�2��L�YI���=��B�Y��+�h�NX-Ӎ��ze���.v�,��9���,l-w������NA&$���mɟ�h*��>����6��������SI�ŕ�
['"�ܽS2$��Wբ2Ճ�ܠ7�R��:a�ײ4s~�,�n��>�T��l��c��2�������w�?���`"(�q��u��
Q�MD��Ll�>���?}���J"u��@���J�	4���A�,�X��LDjy��Z|�9� ;��&;R7��R�"���
�f,��_�˻��|U��M�W��G|���"��;Z�Z�Z��_�Th���Clk��&t�'\@���� "@ݿ�6��iJJ�VK�l9MYp�������[��ZN��H�.��������^}�J	��sӊp�w��Ʊ�o_%4��{�j|���sj8v�,�׭��]0�ɾ�&�j-��]z`�|�:���p��C!����r���gtUEZ!��t@�E!��ߚ�^5�F���Uom��ֆ��`UI2V�Q΄w��a�޻�m�ۆ?����e��D��$>t� ���{|����\,��#�5���mG�T�voR�2S9**s�zW��%���T�m���9"�����3���֕F��X��EB��[��x�έ�h/�r.}�υ�Ӛer�1gT���w�x�25N��c���i�#+[^���3ˏT 7m8�o�q�hog=�{�ܮ�q7�*���LM�[e�rDs�^\v���Q���C��*�E��8[ޫƶ�c�N�I��(�E�]o[e�O��=�r(t{֠;F}�o9�=��g?[�|�zT�6e�����!�M��j��e^�zu��!2���Ip�U��~�a���I�b��2I�<��"(|���x�W�ȉ�B����4�=},J�,�5���ƧX�V���$� ��S�Q�� �Z��i��0R!�q����
���-��#wz*����T���62�<�D5cD�1;IYޖ����w�� w�p���ͷ���b����ڹ;�����4.+��!geEpB�Ş���T2��NX�Ls�� �R����H9.r���k���<P�S�3ރ Ks��J@�EZ�s�W���\�!�p�v�U�����T��S��p�:�E)X��	���������?�R�ցy�]q��v/~.LX-�չ��ZW1'�Y�OO�ŞZ���.G=��Ʃ�o�p�I-ߚGIlH�j�Q�P�r�����OH��
���m�=KxT�Q$2�ݦ��p���]�B��j�8B�{HZ��RA/}\����\�%4���!�Ǫ��{+߷�ښѓ�ݷ�9Of�a��C�G��|�r������e��SAn_��֕݋x	�	��MO�p߹D'�˷��4O�>B������w�'�Ͻ'���V���5t�|T
ȉ25�D)oU��"ԩ5|e�c�f�_�����.�w�����w�Ee 9jR�_�.zzZ�=�6󻛶�2�۶��Hv�|�k7�����w���
k#T�՛ẁ�Q1w�������?�P���u �RV�[���M�Q�_�җ��=?����~Ơ�4�/�9����>|�p�ǽ����tf;x�`�D�خ�͛[�.�1<�q�FdMS��=�X**rRh}��B�:�A�Q�������	�)�8K>)�Ҡ�-�-�#�|�=*Q�'Ξ��Q� Ϊ¡yԆ֙v#oF�R�b/��G�?E��<)�E��b�~���ĳ s�DU�H�sF2�m�3��2zȻ��dcM{)���~���(w90h^�yv���C�'N�����~�I6��(H�(�m�Ml�_
�N����)���%ݓh�t�|���d6��	@��k�~Y�Ub�s���{�֠�����]X����M��4d��js����J���>���-g���u^�|���Ek{�cv
��q6���Z���%\`Z˱��܅�����GN�*�	���b���Q�w�y+��'��cTN�SNzIn��`�?/�{7��� �*�����ق�ۏ�|=J`7V��,K����+g�#�n��y��"��*��P�lS�b��5���ꡊM���/��z8׹�z�l�h�.+x��H�iSr�0=z���g?�	�k�W��5�x��g�W�=?� t�G��ko�z��p���{�`k����t�b����x�g�_z�<��tM�Rr4C�6y�n�jX�s���6�R��������E}Ҕz�K�oW��QЈM;��s�Ʃ�1k�v�X��2���:��N�J	�]�S.��u>���}���Í �(9�[O�\�PS �����Q�=e��K��<���<W�T���1 O�	B�c�NA �kV��P��+�����%j���y�Uu�4?A��iM��H�ֽ˦<��?��ᩧ��5\�ç>���պA�z!���hL�^^�u�΅����a����^KeI�,�3�l�����N���9�V��S��%4Gj̞ ���l.�����������s��"SOz���sou�խ�4~���';����3,ş�531��͉�S!�l{?�:�G����4JR'Kz�Bn%�������)Р���|2\�0g��L�X�
嬍Y:�>���wh��j�@�9
ގ�\�ԯ�������3_���Q���L�y�kJv��tp�K���7��%]����Q����2����1�k�rh=̷F@SԅO�jJ��(j�`?�r��s�uW�w��\q]W�C���̾���&�^��l��ּ�|�+Jx��a�u*�q�P��7<{�w��ل��|d����?�DاކDe^�V��%������/㼜<���l��cg����.�R�J�"�f����@�������.��rk��5���RM(s#@:��gl&�2?�2�ַ~2��HD��������>w�(E�ɻ����S�����a�7�z�?x�p`��E9\%���5�	#����s����mÏir�}a~p(tǡ�=z��p�<@'�����H�2�����DzJ�V����?uo}���+�[�~M��sX��G)FaS6��1�Z2�Ud#�'���[�����Uۇ	������a<���!��#��5��ZR��/���`ޗ�(u����hz���l�F�D��D9��Vqv,L�Q��7����}��P��ӷ��}�N�{=�֍��Y��Z7J���~4�ѽ��.���2�O/k���p���|yf3�݁~�z[N�oi��@b(��jD�d2dD2�m���G0'gUWA���V��-E�<Y���JmY9!�����U�1J1�E�}e�16*���f �����LJ���X�_|��U�֣�+��\UfDC�� M]W��?�U2�j�Ү��q�05YkVT�ڒ��r�D)��"2�1q̲8�kʥ�C
����%���1" �_~u�:s�{k���4���Rv���x{�΍����B1��{μ�����Bq5�ߔa?��@��m�c���7a�l�2`�r�.�)��'�7?eN� ��eyf�g����-Q[���e\ʡ{�i��Z�Bp�!@��\si���;Gy�g���������3}���w�����?����g�C�JJr3�M�lm�I)'�����o��mO�|�������αТ����FěWQGn� ^ۘ%l�l¯{D}�z�aU�	����|;f̬��lt��E>���ڸ�p��~�0A[��k7�M��ax 2Y|��q�����;H�ov�����(��D*���P�|�^��%�!������a�{�O�3��#��y�ҕ��#`�� ������M���C��t*]�z�5�N)�R�k���|�s�:C�d�B�ѕj���gZ�b�lhpp�S �'	�&="�&�=�z�!;�ځO��2(rrג
͐�zz����i5)3��l���Rr�%��='ajäajc�̑�z�5C��My�֋w������W� ��a��n��+��݇rè]�&-`w<��xe����R-"�>K�u}�G����&L�x~��Mi�B	I����Y�&�{ɩpP�7q.I9��Xq2����3i����8��FA��|��� ʕ����6\�Y�ab�=�r�4�̌M�4o���Zn�Βk����S��=���P��X���
4Jf ����Mos�+�{����>M����|hЅ�^
�nql��`��0�}�m�tם�l�,��$ę���'�vX]���o�B��c`�MZ��������/S�<�R����J�B�6r卺�ݰNg��G��g���͔������&A7á�[9�`�����л���aʛ�`p3&Z���T_{��J�Ɖ�w�6M/�®�:W'�螺���Z
���w�4c��P����_�����������=>|�?�\dr؎�����j	��畅��̮�����aw�:�����Q
��Q�S�Ү=����5OsT��6��hj�CeT�y��U,�\=�Z+FSd�ByM"<�Pq��e�wx��O�tt�D�r�z�1�x��i��w���"B�'?{a�v�2�y�>x�o���#�w����e��+����|�QhUOsN���<��ZO��}D�����T_Ö%�Ǩ�^स-YJ՛y�<b�A__�%��fx緓"���K-��#���	�p��В���Si�{^��4+��y�*k�G��ʡ���1��쑶=���(��U�A�Ⱦ���s��#�9Rk��!�,���wc�˓��F���B�G�=�vT��T������'(���xW��37�!;�C���b�B��?�1�/~k��_���p�VV�+��m�R��:�*W/��]阤ɍ��5�������FZ#@2�+�A�e8�H78��
Y��5ra���o���Qn��D�lq�8����F�d���H������4�����9m�i�|r�e~OM�&�1�4��9ڬ�f^���0�:=9}}���DP~exܝ���
e>��:!�C�yB�YL�lkU#�_�X.��̟�O��B�k�. ���7��A[�ϒ~=t7z�\����~U}v1m����ũ�f��"J=�t��P�
��W��r�����x/��&XFQ�U�ܬ!~Yb�P[��區��|s��?q�������+Ã�߃��cSA*�y���G��Ͼ���ir�z2vW��(�'�9�#_�|����kx�����}�P�lKK��tn��ix�]�����G�B�Ѧ�� ��Yb�MJ�e�s�?Ԗ͛�d�w�����A�� H��x�s���_��_����Q��>�7Ets�"���ӝ��Y�ǆ��憓��"�0v8�5���Lo;b��A���|fEՍ����u��o4\���w[Qh#z�q�أj}mEV��0#5n~�~�)+���D��>�:_?W�f�W1���s�����Q��ڃ�Ǩ��s5e\�R�JԆ{L�Q~w�܍�j������xu�=A��``��J>���*`���.8�{2J�Bc�K4�Y�N_��
�<�x��u��*����Q����\���$��k*��eO,�[��0��<�g)��~��P=	L��d��r���.�yE�:t'�����a��&92���&�����+
ԁ���/1?�5��SsD���O���C��Y��>�(�]>�k ����=`�1X0S$".��O�y��*+34x
�D����إ�2cB-�T֍��+�:5��6���y,*:�Oڕ��W�K�B/^�*�"Y����	��ԡ6y����jFC����\3&�<���,%t��6r���Wy�������ǝ�SǪ�e�{�J)���+d֭i�k���6�߽:/,��D5�p,�1�h�в�G} ����
ݟ �	�:t��a��Y��o�V��h4�%o���������α������^ĳ�D��B�(:�����w���|h�tZ�>�m����{,��ͨ��4�J���LِR0�~�k�~;y�4΀|�N��������ʅ��RΡ��"�,��kO�v�5�H�iD;l�=��sk��m�<u�*y�R������6K���z���Rxױ��ڐD�`1�T�� U�5�1��)���T�.LyFx��(�}��#����"�%V�@��:��.�hĪ<슆%E�wM��>�����hV)�5,@E�T�������wϹ{�l&���D���kc�#{�{�m
3�>�a5kꑀ(�6c)!m�be�+��5KT뽢�'���-O�I�����>�;~���ʔ�a]z{��M)\�5��	'��x�z���`��yd����j2F٤�d*3s\Q��COz=�����b��{����s5��<s}������*״]�i��9�U�)sl�<�/]Μ� ���p�'Z2V:�#+E6��+e'@�h���z��8��}��Np4�Q�Sj{���9��^��˝���x�n��iEq�t�*I���Vo�O˥��9e@n|>iɚ���R������*���??�������y'e)�.��F$k)�ch�f	��{k�i	l_QTA '�)y����%)�>���zt�����P
b��
\����b�,ky����Ob�9��ޠ��n�P�`�+;}�t��NQʶ�4�y��%�X3��07"�� �>j8F�>D��=F*`�UJ��=�]Uޣ�է�r轼�MY��T<	W�sm��n I��6֓yS�Ҩ�UFEnb���ю�.ӣٶ�-L��z:��h^B����*%��=�F���t�����Ի��^m�_OuYԾߌ��F#k�"Z.�>>�H`�%Kr�w�Do�K�(��<���h���HS��Q�az|�h��K0�k�w�olM��e�c�T���b�O��t�X�{�Ae��Ux�GBۮ$�K�޶�✶�(�`�ۢ����ާ��{����!�ƷzZ�_�&!�Am�"����?��9����
�������Mb�t����hY����5���3g����F5�VQ)SqQmkժ	�JG��3:�	��Gj)_ݏ䶎�bo�1R����V]E�z0m�۞���H�^k4K�p�f���@�V�kx�ļ��M�7=&��Zr�L�\�``߀��=\�z����.ڤH����Fjh�T�����o�B�r��y�ڟ��i��.&�֖z�i|���bv;s��Y�-$������.8������~yM�Dh�Φh�7�p��>���)!ַI���ؾ[a�zV��UY��e����QF�E�W�~�1�u�q��b���1��w?����~E.��5���m�ַ�v.K�9�?NC��I�S@U[6A�I.+�AE�f#�E�P��@@��(3 z���5��:>#-��������f<y�2�����;k{oFa5χk�h����H0�P��@��WB�z�M�I��egT�el\�u��=�Tv�J�ܐ{u�?&��T 7��+���y[3��B�z�.�&l�zZ�Vk�4��¡|�cN
cQM^<τh`��1��5���m*m�6�I;;c~ݨԜ��6;��S
��H3>�;����^݃	�Σ{��*m+��P1���]%\��|u��XZ��?�Ԅ��	����)�B����	�O�������
�I�*���zծ�%<r��_#�B����^7��:��m<*���)'t�Z�Жr}�9��w��-��.��B�1� ��K��\L�u�q",R-��^q�'�@e�"_*_���a�X��,�+�a����^���WC�d�bn�P;�1oB�{��9N�H)��a�^��%d
�G�;M=9Y]v�>*�	]Y?�IOl05��b�!(}o��톗���Nw�A)�p!��۸@���L�R���
�Eu���ѣ�=��#�v�%�-K���^8�'�Sea*����j�Py5��l�2˴=��%dz(�^[n��[vUx&�[���E4���j0DpU�U���m(Y��R��$���u�Ⱥ�ٮJ�U=p]S�ڇÐu�Eh☨���_^���\d����,M*u�^�C�bG%�)��^}���|�M&$@�R`��{;J����	��̦�k��Μ;�/�yj�}P�NTh�<��S.����",9�"�Uw]���ސȩ6h^o�n���d�&8Q:�!�Lad����g���K8��)�*"o��pl��W�Q�"z5����A�./�6�h�7�h�ʻ���O�Ys?m�eR�km��(�����ϭ�mK[\��Y?͐qB^��ܯ�$*L<t�Ή�78�!�Y<F8��K��/�YI@��f��$��2�{>����;��<���nh���K����{��v?f���ki�"s_��<�2��x���9�EO������ն1����iH���R�#�5n? ��k���C�޽��s*��+Dk�����'��K0⥏���m]ז4���� (lFf��Pk�)*CNe�m�v*O ����3�z�<�7���j^Rk,K�-��e{���4P&�Ȼzm�tq�J���o/B�;sȆ9�k�g���9p���x�<QRx�a��]#���q��Q����iC|.�c�ųW���&�u5y��̉{LB"C�v���!��3�\�ק!��s���D)�hJ�����I�%,:J�I~���j����. ���޾}�y�Q^���WA^�-�x�ݹzoL�
OB�X�.Feg�^)6y�K��քf)��~rj��Z�Uy���V.�_��J���%�ʫi���T(
��!���C�B��6[)�R>�g7_��X��������F�<��M*��?;�ִd�)��˦��'�@�{MH��3�۶��{�ߤ>���,��T�7K_�^��u��
P6��@�Z�@v�R�ʏR��Gگݼ#�Z�PRy���ѨK�Om�* �c���lZ����W�s��{��a³�'#�6��&�<����Jr��~T����/��.���`��gT�/���}h�;�QcR�q��￴n��w�W��<f�Wj��J�����<�0ev��u����̺?4�g��)ˮ4�Q27�qZf��M�]e�����s2��v)L@�k���5����X��8 A���2�;kZ�r�
����F���c.o<���_5�뚺������fhTX�;}���r�+}��w}/�9~Vw[��zP��A!7��N�UqKh!k��׾�ȷ��&MaҔ�2FE�܆���Ŷ85�-�z�=����� �LЪ![����p���-�YO��fY�LJa���(ps�!���K7�ٴL;9�?q@�>�E���W��G��dm�����)�6���H[����d+��睂��7U�e��xV ����FoH���ۉ~�=���j!�]�:�؛/���E�_?v�'�U{����UٔZ6�ĄMF0�vSx��v��\t���_^y���th���U�>
P��l�'U&����y(Z�10*�ݏ��S�j�\��%j��m�z��Qǭ�o��n����cc4gY�uab	� ��A�ڰb�^Hb؀�傈.�c�M���CW������ȩ�7�S����=6?��z2���F;x��
��Bz��+]�ڍ���{ }"�Z�l�B);���S�4�����c͛�^A��B�"{�oC2��0��ǉg�G��q���4��R��L'V9�7\���*V �o�{R��/�~5=���z�i�#���[e�Ե��e��(���
r-z�2m�U�YEq�P�T�i�'W�{-|ֺk��5�Z�)c����r޺�j_<���j�3�BʵY#{;��Ws�μ\@n���`��x�Kq�5��汃$;m�,c=Џ�g�r��d���-K,�n����Q�F��+�ןj���^>L�;��W�n��[6��KM���	ʫnB�R���%�������҂��#���&3e��m�yx�Y*�m��s6b4y�%�4�z�\zO��et�,��7�~���;ÿ��?����ȅ����x"5��?��&A�Oo�gh�D��,q�݊r��30�M@_;�ޛ�^~�,kCp�DL��m�k��	��d����q�J�D��g�Ƙo�R�5Cwc�4��_nz	��"�^1߹�My�M�_em�J���>��+t/���CG?����>��G�6%X�E�4kcv[݄V����&�`r�Γ�
AB}#V��݁
�*p�KU��4)�ڿ�߫�s�.�VC�K�ӂ�X9b��{[S�=4�OX�#&ESh֌w�VB��R�ȚR�p*!���ߍQ��w���}���n�������y8|�a8��9�;A;���*���i6�`8��oË�lF�t�Nf ���)��<*��Q�y�yTR\��cZ7����v������3N�kc/��-��!��X'�ە��Ä$׳��P��'J�NP�FAX�[��Խ�&p[�fdI���S��mf�a���J�u���rƨw��F�:F��wM�B�R��R�ˆ��AY�/�/ ����V�š�5��~����s��(�j#�c���ɨ�l7�_�^�ųF��a�ʜ�~�O��z��$��:�F���q��t��^K��t55V��bX*��+�>U��y|O�6bX��wc��^�㔜{���cu�ܿ�e�����e�6D���X�\�+�*gL�AnkX= &!��>�1�-T�CC��`��K�?;���2�ub��*�uQ��x%�aD�h�/j����N��6�n?{k���M��Y�SP������o��_C�&O/=�S��<���;  � vk�7�%͞��nn�A�r�4w�n�ȟF�4��8��<�8������X�ʍU����w"�M��U#ZC�K�#{�{ǨY!2�����Fd��7��=��n�S_�#���;����?��z��=y��}e�ڮ0k���pvE��	@��(��5r6��<�EQH�� =B	=����Z݊��̇@6v��k�W����B���c�s���n���	�g����,WJ2��#^���4ή��M�F�.7�@aQo����5���ۄ��<m���_�:]������#�
|賳�C�)��B��nH<�T��f'����Z�BF/21����.�T��K�l^�jv���~j�k�x�M��C��i�;��7�:>���2��+�ʣ��Oמf(��Nb����$��Dq�[gw*�+�޽��t���HJ��+�c=��$��,�I�
j�����%�]�\��E2{�QT
"8�'[�YE��z��.e��d^�:�*�*���bj�� 3Ӎ���b�FU�v���2/]%Iŋ� ����K�����\�,��U�dH��hZS�}-�*G�"
��\�H׀��^�TT0����m�w�0G��j��?4fF�p{Wv݃U���y��2��L�w�^��52�'��S���q�0�:X�1�Z!�c�_�QEW��3(���W�:I�@�E�1Y='H�Fi3���ӛK�E��r�9z��4<�{��ڍV��5���!u������[!�Qyʵ��z�z�vPGi
,��S3#(��.~%|E?�ʆ�|Fj��ŨK�
q����ˮI
�4�RX]{Ԭ���>�#�;&,߹�Ǯ�$z��8ձn������C��#�c{�С��|��?Y��e�p݁�e�/����!�B2�w2^��C}sv�9f��@W����
��|��n�_���B�a~k�ƨU_.�W�TB1��w{��V���}ЈX��KH��I<<�t6t/-��xS�3' ��*X/|��D���t��Job�-�w�᎕l9���ۆ{��3�w쨭��?K���;�Ev%!_�=��B��ă��J��W�:FJ	S�Gypx��#�������O~���"%s�-Mn�y�y_�M����e��	�"$��5VB�<5�����T�^�uK�� ���j-���-3����۵�r�Q��b�1�mA���o6��'�y�(�DE�U8z�*2<�fl�Ll��"_O6�B��ʹX��C�UZYG�U�M���:j�����8�����.��¶v��._c�R"�xg�u�鞴M�s��(Z�Ѭ˵����m����{�0��g������7�A+��XU�^\ka�sKeh��51x�qk����:#���i��Wb�pv:<G$=����(�/i�J��hv�)0[��Wg��W�k�|1D|��ܐ7@5�0��t���t�#��
�����Kjʰu�ߍ���;�W�]�b).�P%,�®����V��d��Z�σN�awK�TO:)�H��}g�ȈT9W����PTk d��+�g��9���9<�dSR��35���^ܼi����ް��Ũ�y�����4��,���?��]������] k��Rmֲ"�wt��EZJ@uϢ��`x�6k�F���9z^~-?/Ɇ�
���̡G�����zL�_u�����댣�Y���{�ĭ�B�>�Q��=Gk���l^�<U�P��k�`ޣ%����������vV�1�Zл�>D9��a���({�l
P�l�KW/�l� �6C���'e.\�ݐJ������|u�N��饾m��i��D?{;%A�;#��&:rYs���В���Oȶ����]%΋ ���'|��޲hh)��j�:k�c��f��<Z�)�!��8�8���m�r��u�%�o!�4�����%�j�����4ae.Ѷ��6[I�av�UpH��F2��F+^�%��j���Y���TI�_�*�)��������fR�C�e��HE����"�5���zԥ)��e����#���IW���ݦ%�M�W��IG�U	36��>���Q����y�NI[{G��:)�yt�|������*�A��=`��P܆g���r�]�b���DO�*:׸��b�2ec�=ZC-�8�3w_�̽R�G�ɫ�W�[`Π� r�ȅt�t��G��[���J�VK�O�uj�+m�cV�X^s��
`Oe�.�A���k/@Jed�8�!��ލ�T��J�D&�y[���]�r�����U��u�[9��l�M3p���yҶ�R,q��;�C�bi�����~�.^��Qf���P�׼������]�zJ�X���t5TX����c|0�6�ɏ��G�A��"A��^������V=� .��߫�B����2WY�
��l岎�CI�b��x��ݴ
�>1��-�������{���.j��?{:�}{�K��
g��=á��Jٚ�]��#n���e8�4y�rB����	��^�
�=V�%�2�
*(~����7��|���a~� ��=�W�Ͽ���/}���{����E"Ԕㅌ�Ӗ���8��lл0-�� '7�"ׄ
�Tȱ�v�p��U��2���Ƶ���`����q�2�eIR��4�D'���
 #��z�7�'Ә�oh���oܓ�Y+Y]�	���nƳ3R�s<����[_��D�f@*#��j���dnу���L@i:��x�Q�^97F���������(k��1P����K>�E�������jF���\��Wv�}׼lE�*ZT{�Ǩ1�)�W#Zm�z�<�� �|W�V���u���YJ�Sk���5$ś�W�?�,W�=��<�1�9n�x�*� �r/u��u����]q�j|��Oh�y5�2%��Ek�����Iv|�$��ک4���u���b�����@ȑ�Izs̧�ep���-31#��! �͏���R��V�uQH~�Qr��ַ�H��-�)��{K.��@��Z�R���㱂Ar�肱�M���������m��y����Q
�����y�Ϗ�w��/����K���Z�K�W$eTi[��.����~/�h4�֟w�V�>B Ѽ�x�V�SI�.jw:Ey�׌c@?nZ6Gg٪�e�0Z3.�N�W�ݐ=��kҋn�<=��x�
�ΘWQ���a{J7d?��к�w�=>�������'A�1K��$��=�n�V��u�Nj��ފ��8,=w�MenQ�ý�����HR]��WYm -23La\L��,��%��MH$��3�����O|lx�{�	B0�m�����P�ax�/�� !�t@l3F)ڵ�j�x;z��n�2$��x\�^�� ���߳"!���(�b�Wͻ�y�m+�}g�����US��\@���:���J�֋^�V��@	xv��2�*)�Ne�3�l>����
N!hl���7^YS~/ec�q�P0�èxg��MMiQ Q���Nn&҂����^�K�YuM�窀����[�)+���j�J�;k��o�.���+S��ז{r����=�l����VYiy�Ω�[ՔݸU�������Elb��66��B�IM1����E)��a���SbxM�fK���A[""S1^�Hw�a���7��0��(�Ҁ�h[�iL���#v���W��rx*'�@X\{תUMO�g�ZQ��X5�W��
JZ�ܴ��ٷnc�D�N@ش� 7M��ē��֔EmϘr}jb���)��=Z�g��ޫ���j���Kn�@����r�	����p�X���8�k�ڿˡ����ۯ{��G~��o���'��ϔU�� G7q�Ȳ�w�':����S��,����Pt��.��<��9�JW��ʼJ}v�Z��ݒ�����楤�(���m�\rX�>��CV���<q���(��u�Lϧ�6*1IHS�\�~�1YO�x�^�����7}��|Fp�ŋ�$U�	~9�+�Q���:&��B2U/x#a�l@@
)_� ��鱨#VKj�j��-�tFJ	8o���M��]���E������	�y�y��O~�Ӕ�m^}�ᩧ�f0��&0�rO��q��-���T膱+�Hge��7���q*T�9�x�h4���_R0�KB������s��R�׬�@�[�,�v9�z�Ƭ�o��wc�tLq�e�nb4�jVeC֓�!<v�7�w֫�+���c��ެ��I�t\n�n֓��+��<���n|�=�=��yo��e77i�+�3^S�����GԸ:FO
]B����W�\�cm/f���n��%#
��A����B��Q4|R V�s��)���U�P�0��
bI��j�M�����0Ÿ��@�9
�F?R[�����9*2_�������%Rs2�z�o�O�u2
<`���Z�;E�8�m�\��kF�
8+��ll�o�p����G�40*�P��Nm�y:kc�h��e�)�kQ���k��9�~t$A�Ǽ�fER�g./��������ܦf�u���n�%~�?�(��Ɠ���o��O~����εw�
�mM��O�K!���n���&\v����=,>������r���ѫyLSAjn�z7�S�h� y��D�aK0G�E���jy�,��N��j�7=��5�^w��%�J!�ICZ��$�p���s͎9}�\@*ָ��>O�tۢj�Oר��f<�^�8U��e�w�<��)�cJ����ޞ�VaƉ����Q��W�x��p��iBㄉ)?9:i8��+
�+��u0�{�9�Co��Y 
�e�����KW��g�l��:k�>Fu`���=�ha�H���$ż�B�:�fg�����&-��Y0b��3>�ɉ�]θ�<�z�`��I�2��LI$j�D0����;�@�}>��5g��)8}����S�8������K ���L�b�U� �8�\]Wr�^7�3*�������`��)k]�6��O�p�S�Ѱ��2�F#i�8v�b�����V�W�T��徎����;�jc��*��h�����^���ⶣ�y�l�^��,O��*%F�>3��ܯ�o�3ctdl�0�deT�'��r�P��!�=�$+C�s���|?i(17��ƍi���:p"L	K�U]m��Ϥ[7�X�ф�yp �)j[>n���^l�`�#�m���^�p���]7&�]�ʯ@K���*�3�\��9͚�TH����&�Z��I�*��xk���7���ٗe�u�wj�5O=w��#A� 	��Hɑ,ڎ�ر�(�Z�W����%oN^����!��Ȗ5��(J�8�	�����y�y���|>{�SU���$f�]`��{������w��8�~�?S�a��7Pָ�MGLL�v�'{�;8Ws���_8�.��.=v��O<��^�I�r�iC+Nc������gs��{UH]�In�X>��Ra�`���eБq�ߏ*���ռ���11�AxP��ī��JoR��5D�H���n��Nh	���	�<�!�:UH��t��aN5	AG�t?1N,��_uPlf����֙�����|t= ��M{��(��o}zz�����(t����x�ާ9�������`�" ���qOӄ�O��b��&d5r���	�,	oI�e�5��͓�C!7������dx�E�t��s�}9:�eD��
��e-]�2��z-r���t �a�<K�B=���~T&��ғ��zD�v�pI��=nz9b ���ǈ'�/#&�Z�'l�����
�\y��K!��3R���Cm�;�>��6I�Mf�x��Di�h��8K������ @�%!�#�.�>P�]N��^��=�w�2���	�vjl׹��$����iNg|w���~"SIATi���9�N����?YϞ�^�=�)o��3M����|�^ON���&n������om�9�y�J\E)��h�x9������{��l�׾�$�ͣI�/���
��Ԅ���=�1B��h�#fp�!�f<��D���(��c�mD<2�������*�#	{D����� EZ��=D'H�"*�L)h\YZ��Kܞcq�b�rL�mD����8ׂ	YȵiL����ަ5����w�R9�FI� hRcZʎN{ �ďr�I!�ւ���=w|��B*t�������w��ݿK�����z��<�N�hݛ�R�_g�wT�S]G�7�^���oGO�E:^���*��b��ӷ̹��[�Cc:A�G���BID�7`��M��m����� -�0P2^vH�SQ��^��K-��c�x^
B�#߾�n�GMٽ�����[�6[�k��ff�bn����m�0�ܻ)n}�fl�a�B����/ޖ�o~�s.��i��4߼�$�5<�ȹ������g�����m����7���w�ſi�,Fx�����[X^��:}�/##�51�NR�*���R&?�gM��5������_��*�4>�/��W1,|�Q��Q+N|m<��*<��Fl���]�G�ߵ8��C/x~&L�قYld�#�����̅�"Sچ�����4��^��|vP%�k4K��z�B���I�"��������w��tC�f��b�>�X�_�܈�5�=��)��}��#L����k�e��+a�1��s�~�s�]ĵEt ���;�	����{��Q�g�|6Q���y��O@�%,���\v����D���W|�Y\�on��sf��YE�A�摪�#��ܼw�=�1Ҵ%�-k#E�ͣ�H��d���M����!���:rī%`��`��p���O|�FK��
=B	���@�}@ӢlqluG�~z��s��*W�Ja�V �o��i�\�F,�tn���F�%r����ҍ���m�p����p��zpW�D�
��4k�p��l�\;���R����_�̧?��_|���k͘j
F�q+�:�"�ruq�� �E��S~?���Xy�.����R��Qk�;g'�қ,)��@P�����p����E�r��k9����w�d���8Ɣ�P�{X��O|2����nld%sv��h0i#	B� ?���;�34�ѪwF�!x�D�s�3��ͽU����ݏb��m!�ז�>=�wwP�F�<c4Pio#�`�����������e��fh�SF^�F��������y�=J�h�y���S�>�<���{��a�S6G=��[K�����f��x�/�I�Hң34m+�"������3:�Jo��P8P1:҆QYg��e|�Y�����mg;�"I���m�S�a0{kgiZ����2�c=�.�N}�R�ʳr̤�0E��������A3�ۆ�U��"�h��$�\��k�	��Ur��Y�$4������iC���Q{�3&�ah�y0,�*m�w��\�^z-�P�i�vFa�{��J���!�H[D�?�;���z?�9k�� ��<K��|�:c����6��:�9�Uʫ<��ʇ��MQ����Ƕ��Pj�?��盿���As���w~�f���!��|�f���g�ɕ���7����4	.D����U�q�{�E�u���>װ�g��OC����͘q*��j�l,�I�ݧG{C鵻�$�EU{~8�����q�<�����"�(�Ѿ�9.�=ƿ������T�t��r�������C����6�Cw�9ʚ0�GF���L�c����Q�������޹�Η)�z6-eQZ� �X(��ܝ�3��b�M�  :O�g����zj���G�~4��{�ߏ��'?6*�I��3o������Z/�56�^[��Q!9X#�z���� �������z�,r4j �������ߧ޲�<��#��_jVP��^~�ы���w�!Źs����6|�@��K|�M�'���b�k}����-��Q��?�'�L�4���Av������wx�4A*��ƕ���7�n�^�_��fk��/|�����o7�;�,o��L���~���?�v<[7�ʧ�e��yq�z*�܍��}��ƂҊjy��9�p���X��7��w)nOj\i�v�IU;�$���G�l�
+j�go���ni��K�>�]�a�D>X>�$�/\OˈI*9�~��n�$3�u�S��D5�H<�	�����>
ì�Y~��i׻ޤü�óm��#�z���o1��Wǌ�k�N���E�'1-�B�p�Qw$Y�%��}ֱY���f3݊W^G����|w�+hSU�W�!��f�6��ڴ�!�k	c��"#}���C9��V�ȝ�Q�L��n�|oǶ�e�V�s��G�n�.R-2��GJ*�0i܊Ib��8��탧�@�L��*cֹg�!¬�Ñx�c��b�H�tI�4ܝ��\1��p14㕩^��Zq�� �M�E:#y)��E7�s�^�����ǲ����]�/GbfDF*��d$G������B��|�"�N��k������7�L�\~�М�����<��u�5Q
�`�����j��͛W�����������,��\��W���*�����b�g_K�4�8��1:��z�H1.�nPDw�N�t�Bl��u�������M�ކ/����γ���S��Q"��Vtk�dC�ױ}Ӓ>,�jC�Zˎ���6�G}N����n)���ԙ�a+�G.>�<F}�Y���k�gt��SgC@=X�n��v��H֭��lDH/�1!�z�a��/\8�����͝[6��4�y��aA>>JN������w�S_v5���B��޿����1emO7���'�'��c�P�2B�
+��a�C�J�P0o#W� ����9�
�}��-��!L���x.
#�:�|�B3��:'~e�6Nw�0�{�s�#qy��x�o�8�����1#<1U��P���u����q��p^c�-���vJ�I�==,יU �B�㤰F>S~0jԡ����#��W$!��Tg�Do����фH�ۥϞ���7�RD��i<��u!`�U�������du[B7�z���;�u{;r��B�������E��Ѽy�=L�������q�vv˞���x���"?g�(�ߧ�g"��xQ�WK���g۬�m,��ք^���n�V]Z_l���+�{�7�i�Y���"�z����Vי�
rr�`�
�XnYFe4"$���yn$ͽ��*�`���q���xSWØ{�^	m	�4�����n��`��H%���(�רlG�O&"��Qޚ�6��=}Z���%Ⱥ�H/D�Q���#a$�����5<Ԝ\ȱ�+�c�H��I'�8����с^o���J�\�����ԩ[���g��G����>�~��]غ�LB@�J��=�\}��&鄥Ū,�)�±��b�U�'�CO��ֈ���?�u���+G��]K����#%�?#X(�<#�IC}w�kO�5�2�^KE豣�*����襴�?�GX�=��[���%�p>sU*�ȡ�8y�Ts�q�
�S�<�,�>ǆ�5F����杫7���o�e��ɨg6��W7ќ<s�cΠ�7�w߹�b_aR�B�����:�uȆG��$��������.9�7�4��/7����?�̟:ռ}��8���y֎��
;1�, �h\k�M��4� �О�����'k��4��)L��,+�^�k(t��my;J=��(��V�����l*�\j��x��3���ꈃ�u�����K/k���!	I-�:(��7���i����0�l�bL�G#��X��kǝ�P�~�5l2,�sJ#4�D&�(��ni
.K�_7l:��}�����l\��慳�B�b�HI�V�����_�ͱ��[�/�.�q7׼��G��`m�oɆC^��k�kP˥M�gɱ3�`�adb�Z&{�J�������o�ܻC_vHj�]��
ē7JC�gs�~c����z3C�e�����(�h�yWW�ھyg����f����� L(�rd�^��lf���}��"<����>�� =�>	��6%�q%C>d�F�'øK�Q�j�x���0�N�e������B�{�T����Jz��T���%�HDo�g��C�9N	��T��|�4��[4�Ʊ��Z������x�S���G�x
B9�G
�&G�y�Ԃ��w�1��/؟�	��ӵ�׺�kחZq�%z���ɯ���Ʌ�}����s���x~�ŭ7� �����*i��¢C�
E�Ǉ��\b~���BG�4B���������V�l�}XcnyH�F;�P!�h����rRkz�ȟ�?�k��g�u�_�淛7��l��2���̏����^�����Rs�)n��a��_~�����C(���:P���ϝk��o�6-gO7������?�I��dS{� ��{-<�1�(�Uo�� X�#4y�� B-V�THj2��>��%�>�T�)��d<�x̆+�#ސJc�TũS'�ڲ�W;����r���9C�wQO�^|�;C�[?�)�%_j�@�lݿ�A�x9��}u7"��]�B�1v�#��g�G�x�<G�s ���  v��s'¨[�q#�6�"�>��J4R	��P�vޱ���;6�!���-�3�����9�8�֜��~��Ј�[hD9b�m��kg�DH��Bm��S.]W�a~\�=�����`�5I�������ޛ?{����:d�:�ha� T:�z@Z�އ 	F!�LS��co8�O`��i�Djc7Z�F8-�/U`|.T#���s�w�hʴ��ua�Cb���о�=�H��k�p&�so�h�`��V�����b�raa��S��{�0z�ʹ��0N:^�21�g�fHB�xA)sM��]��ht��6�Q�^�������}�1�K�:�B��1(�u�J�a"�`���pB��.^y�����"�{��_�6�?��k�~�������]�l���>3��!�T��3�jC��wܒ�R<�B<��2����w��5<z+����l޽����vm.P��EڒI����G/<��>ͰZ�b�}v{c ��� �dhSoh��h����~��<8�Q��>�C�PzI��l�"'ڇ��&�8���8��Ge��<x@o������揿�fMB�^o`��)���j�Y�q/f�!�c��U������	šQ�-���O����5�2B�Cd&��d���5jӱ�	��mHv#��� w�ݯ�"7ji�ރ�D�f�;s���KHC)]�C��]O(T�Y�U�&�T��4���83�5(Reg����&N�a)U��a�!r\Sg��|W+�r�&q(�P��j�[$�E
�(�� �m�%�S>�K�K��YcLPo������f�u'�}vx>�[�N��ʅ}�-<�;����5
x�sv|�h\����B�����(0���@C KO��:�{Z���B��O�e�G�]���:��U���t$Q*J4S*?�Cq�U�;��hg�$��OC�&���Wa�߈5�VF�Qe���u��#�;�Ht��}Q���a�o�N��:��G�&Fnlȣ1���my���*� ^{�`��j�^��9�{G%�1u���s�F�H�3�uGe��&�7׉�i � 7��	+����^:�O�� ��'�ӈA8)V"P���:���S��P�g)������qF�P1z8�B��gѓ�)�B:#X���q��,t��/���	�_��^�r�%��]���2��x�D.=@Wwn�g�nT��RmI'0:X0��U�#.�x-?ߪ����ɼ���uJ�!uX���IH䷺\q�)z�FO��5_����^�\�jdW+-��|���l��?j�ܹ�ܼAv����L���<����m`1����M��k��\�4dv�]r�!��O�FA��n�o����|������uE%��A4 sz����;�|x�\�n3G�vgt���;ͭ{�x�vY�>ˣ�޻�^m���ퟆ���(�K�����;��_��P���9�����g���g����}ʯ�7�^G��	G�����2[+�՛��k/2���^�b�(�g���@�4�O���)��}��(� ��屍 d�?O�^G�)rMź���tJ,�8nx��HA��L��F2U�"	U>���m�=�����u����l�t@�7�t�{�����G�g?�k��T���aj�gK���	q��:���ll�JD+r��_�(���d7���gG�Ď�����dx��|��c�I~��6��� ���f�y��m�7�0IY|>���L��U�*i���H;6}'[܃]��h���p�I9aX����2*��D/u�ϝ�5�o���9���1��������s	4�~���W�������Ҡ�%63��|Ny�F*L1J2�y�vfA�T�4�k��2)�2��4]w��Ix2�E0��
V���K��*���&�D��{��{<�0���uי���b���N��i[5L�f�>�T�L`0j ������¹��'�z�&R�1�2�p�=;�L_��c%ω�C���Ɍ�#���,��m���˱P�M=x��7��k��������y
@i4ei�󈨻�)�?�uif�]*��Rb�l����pQx@��b�J+[+��t�o:噬���$�a�'f��^&(����{��6?iX]�#kWCXi���l ����L`�z*_ϣr��娤�̑�ם����A��y����8�ę(g��
Jr��,k�C�������^�.������懯�I�o�}� s�J��L��g�p͌��XgN7���f�HǹՕ��������!B��v��=[kd��\�cey�y��+�_���n�CڻuoeI�����C��B|�f��1��1�>��Q�-�7��<�(����͋W����9r�Y~�W���s�$��m*+{�'	�7e�ut�J�,�:H�2�e�s-�S��NC�F$z?]4I��)T�ڏ�e����1:֫1��"τG�jTH�:s��fm����KЮ��LH��e���V�?���^��#z�����5w�>��k���������0i��w~��f��^ZZ�}e�ڻ�ܠaJ��w���j�S?��#AB��ԑ%f�*M�s�qϸ�:R��]��5��g��?{��5����f���WY���	l~�8��'��x�\L{��p�z�5B�o�%N��_�00�������D�a���p�^�לY1�֘JْJ;����gg�rQ�΄)�|p���������Kqh�z_��4�n��e�ӧ�6��?����=������i8�ϟ�K���v�OK���x�x�^Í�Q�K\[�jr��I�����M��ɺ_�T��{8)D
&g��i�T3C���g�O�;s�Tsc�k�����	h�2��n��2��([;v_�B��T._���/��7>����<xx6C�.��=�p�1�<��Oi�f�N.�͎�SX��:e�לy��m�;B�~�ͭu��2��q��F�cR��P��zZ�Z�6����^�~�T�%S\�z:vO2g�ʜ��dBieu-z�v��h�pax
US)��?w�酱�5��y��K<ћҫX��jum��x�=���Rs�@(����F��!��qz��d��$��� [83�d3M�{����I�+�<N�׏��>z3ؿ�Ԑڅ.zr���̟C��Pbޥǟhnߺ�ܿw�&�o��+��Լ��_n����Z�n���%/��ֱ���E�Y�te|�ĮP��1��i=̃��2�>�f댍�I]�#�RqxHԷ/���A@����ٍR�w�y��6Q��a���(]#��w�}�XV�|�\����d�HG*�n�)���i	��>3��9P��	p(����jDo��9��<�B��
��e�U��Jɘl�0�r����r���Ϝ{Kv4�3��<q�D*#PAZ��W�i	��R�<�%�,E�{�V���~q��ѣnB��;���;�M�"okԣ�/ǈ0|��7ud����Wx�m�,��R)g(7Yb��ez�ɺv���+��c�l��KD�%ԙ>ED&�[C�w��r:��yD:�VUY!G8a�a��Q�x���ᣑ:��VXx��v�k<Rg�y�1.���d���>�>���+ݐ�U"\�H��&Mj\�aH�~���z���ݨ�Q�q�;��p��L�<��M̳/�U ����BD�B�[��
��������K#�M� �/s��9"Xܛ2��F�~�Ȯ�P.R\���S����C�7����� ��[�Bu=��\�����<���Sa�u��a�4mشP;�̕���m^8_3\G�Q0F��uu:F�cG�;�}j 
l�˭G����~�f�����)�]�6���V��I��b�Jx�9ElOp�\�3O?��C����u��z����*ђ��@�4'��W�D-�<�;`P�*����+���[�����?|=�h��]{�5S!$�Cs=lę�y�n'���#�t��50�18��ﾌR��&]������`���A����Y�;��
V��o��5�׿�����|���@����y���w߿׼sa2D�{��5����(�9���fԟlk6�<+�(r�>���!O���G��4�j���k1��0r|j���Ț^hz�9���O�A���b����8^�]��٪�<���p�^�2]�T
��7z�%"��hg4 	R�%� 	-��Q��Z�t�g�Q0���}�{��#ͅ˟h�=�l���?͜���'Ϲ�46�5Ԇ�e�o�[�pm���� �E�kX�~��ݸ�u��p7�\Lb�84���C^3Jś_Y������@�ͧ�����z ��2Jѱ�;%Fl4pɰ��%���a`���G�Bt-����:�Z���.�֥	BF$cr]>փ�����fWF�,i�Gh\��>��@�U�ǕJ*�x�i�E�O���;ʓ�Bf�|��}�s}v�z��4Gߦ��|�aı��дL��9����tc�� 7�v�<,�nu��<FZGtd,������h`-p�K��V	��qQ�%)�S]���e��F��0����ĵ�^��V�3$�R:E��)I�C��SA<��d���~C6�>L�}�e�ܧ|l<to��ŋ��~��~��_�Z<�8�lx6�;��Ps�-��"��B$�L��.��,H���>��[!����IO�:!�5$r�V
.[wZ�)�� ��W~�|�s��1=^3Y�d����M�Q�x����{X����_~�2F����;������fS�v�^�ܴ��fJˉT*���*pC��~��#��ؼ�d�oSC��z�ܬN\�%to���ר5�<nn�c�Ż��^Bl4'榸�G��r���*�lj� K�����=��3͕w�mΝ=�s�^����{�o��5�8H�e.?J�ރ�F�ʞC��%����+b����WX�5����_d^�B�7y�C	�$��ģO0��"���Tx�
l�y���De���yd���l�3����g���n���L�c
�%BZ��7u�A%q�4Ó�2��������mv���-y*�+:�+:�2\�M��z�������Dֿ��Ƹ&0P�R�{�TP�<����xt�
�4@�gT!��S�������R��׽�Cś*��a�λ�4���ꗰ|p��s�M�!��?e��+ �x,���WǛ	���Vct�t�h�t��e����}�?Ԗ���i~���"��r.2]l�ċ�l�2�3ܧ�Cy�z(�}�ʠ�@n#��������2U�Ai@���5B	e����G7�Svz�"i9;E��v`�X>i�M#F��&?}�1�V��ȁ��.\� �'$@��oY�*�SPF-��*�`�aǽ<|�u�����PNd����Y��싈���x�� ۩nxx࿟�{��t�:�m��q�'����WSo��7=�����d\�*�С��J6��V���v�ux	*��g��usG����J�dj����z1Q��.�6�/�oWu�BE���[��zv8�#BV��	)�}S(�	6�ֿ�H�q� a��^��g�m~�!�0�/.�n�U��LY"�72���dS�QdG0-e�7���3��M���V��«�ԃKg�s�ᙛ�X���U(]-x=G����Z��f��Vs���4׮��\��Ǧ"�֯�V<Ke6׷��$��=�pq%�1�}�3��O?Ƈe-'����[5���]�C����pvi�s5�N|,�'�m��6L9�2�����N�����X<i��?	>=��L���qbclj�9wz~��X��g=V���;B�5�^�8u��J�{�;����''�)��D=p�lF�3֖�\r��M8��7n���й旞{��9��߰r�.`D3Z/�[k��[���u�K�X���K��εJ4��?�l?�.%�Z72�Fv{�v������a^����&�f�8��!�{��y�q��zޡ{!�vI����;e�ʾ��7�Pm�U^~�[7��=sv[Ø�F<1�s�˸\�q��MິL�j�K��(Jk ��1�$�QV9e��DK0z���{�ܠ���<I7�F�v��Up:��c��9��JA�t��_{���0m��tEK��g�g�<��3���&����SZ�a�M�0"�٣unF`���1~�������Cw޹F����}Hwɓ�bX���  �I�1 v�$�=�G�!J}-��8ǡ5�>����X)tD��/����޹����=>;�q,�֒K?pi�����R�.sS�rm=����Q���!�k919���:F�	��Ó�i��9rz�i)j��nQ! �[
��)7!���G7��v��<TԽ���;F/�GR�,�M�a?�$��J���tu{��w����:����}ɦ"��� ��\���"tsS�}��5��&�-1eM�������r�+^�fQF���ԓ�4/>����1�2���W_��N^>�O�[O��l�;�V����|��Q�x��K�����ʗ_ʦ74�09��z���W�`hc�)]>2��6B/�A��yB pQ��B��SA�:D?�2�%� ���)��I����`=L�6�?~�R��(��òw`�^^�
��O�z��G��g�'5���x7mM���T�l�ȋ��_��F�����x��k�B������O=E��ts��"��&7	%�`RC{�-��]��0V��(u�9���1��v��*�Nٶ��S�b۫��?��[�|8�ۧ���(��?gX��y�qE*��g�7��"�B�]��gv��$��?4<~��ɳ��bDmӼrx*��T��5��=n��T2�Y�7pa�u`~~��Xo*F+7\�A���ޛ�$���`�1�'�6kr)B~�b�=)���12�b������H�$J��1>9D��0������$G���z\���i�|�:\�&[=�,䤄R۷���u�~�a�G(��u#��ǝ����`��q㔌ҋ�	k6��=��Ĝc�u�:^��իW��~���X�_�9�y܆)%Z��	fy*��n[/$���e쯻��⏥�v��nY!"�Y�VTt:>Cr*�l�ϼp�k���gb�e�z�a�g�~��C�|��]�ܧK�|,�Y�鲟͓����UX����-���S |�l��~ȆԚ=�dB��6�2��R׋��V(�$
z͹�N��{W k��;W��5���G����wjDq-*!�q�(|�<���&����Õfx�Q�\�]��3ǟ���bJ�|yy����#?��o�Ҽ~��T�j��_iN/�i�]��b��UrJ�lQú�@5W�Ad6ro<?���l���<d�g�>�H\3
�V@)��w:%r�H�P�fs��у�p�')���eY]�յ�ם^ZF�|�3fb"�zy=��������R������!��^����w����/�����K`u�����J_>��
��O]���//�u��ur��r��YD�O��`���&�>��,�>�A��x�u�@(i��ID=���Ͽyd�S��;�����ȏ>���M(Ep���"�5w���5��!.�h��k�����ll�ޱ��s�-��Jn��GK���ƥX�pA�8at�e�.�=r�`;Ȅ���r9�{��T��d(���!�q�^v�-��<q�L3-�ޒ� ����!Ah;��C�є��K��e�|�K�n���u���r��ȑ�,/Dއ�U��<�I���{"���0�|��gX�}~_#�O�܍��"�v��^%�؃O�\��#5�5;���8�7u���W��/�����g6��';�\&q�&n���G!OR��`�=�r�a�Oi�ƶK���T��26Y����w��<�DZ�q���fX��
�ŮG�z&q]�����s�����i�q�����瞍\���uk��{�)N��ajx��o[�v���t	��>����GH7�Ru�VO6s���P ĿTT�d%�HV��`����L�a�u�@�����/��4�hhX�Iәw�C��z��m����(���?l6Q��u�p��vg��à%g��t�ù�����fh�^�D��;w���u�I28�Լ��¹-��")�1lM�����|L�B��Y2h�,C�v����;����ľ�A$rB�`>!N��<������4�7�8Ƣ���ǰ�9n�F���$I�kc�)��Mmvv��=u�9�~�d�"�L�����2Z��>C�^*B�>��\ �#���|�`D�Z'��_a��T�"�z���kD:iU:3����OC B�]��#��`�yu��܅�;�h�������M~��G�]���l��������z�t�uQ8��ѿu��)�X&�%��իH��,��n� �����|(Cd�GJ�Tp �_tW�?��w�fɛQ�7����������$��p�����8��zO ���'��GY�VHl�������4���}+64��c"���Q(�_͡��]p	>͚S�dv A9?�|{�K@�;5r*�Y�����G�6鸧w�	���.5��§��g.`���,S\c���&��0�#�M�1ׁ�J��1#'m���?�������[o���7���������G_�vwz�~��vdX�Ji7R�M�OJ���(�|w*��ׅ���R�'9UEg������nkSUzZ��o���N��>m�Q7��,����G?mN�3�܋�b����h��v��Azb�tĩ ����c7�?A�°w��1Bɩ��v�2���|t���q���k�L�<u:Y�[���#�^��<��q�Q=K7�����|^k���^�*��k[�ܳ!���y6�F�����벱���G8|}e�z7l�E~��[;\����c��$�-�J^�Q�`G���x�He�]�8�)��#�w����\���JE�W7����!�%�s��Ǔ��j�4���d��g������o�x���O~�q�@�EHv��=��pNC�>'��(,���n��m����\�Ao���7���g�ˏ_�S���o."�ei���9~r�m�!�G~��m�v|�*�a�ƙۻL����M0M���Ge]�r�Ր�Ǿn�����so�������+���h�'��{0�v��%F�/��G�w��Q������G޽�{=<�xV��������N4��$�m�0�YEA��0�c�˨Lx��%.<y�Z���4J1A�������tOtf�c�8~o�tK]�T�7Fk�W��M�������.uhl���`s��4jb*�r�ՙ�8OCsxġ497b��Z1�4�nkVz7�u�c��vpxtbj�ejl�-�d��ټN���g�w6����4����^��j������0��b�l��Ϭ�_�_����Cy����k��O�x�3����c�A��r�k(�옵C�h�j:7Y(:7d�@���h��ôb�l�����6�B��:1&�K��[�Ӑ��KS���(��gRK]'{]�<��6�֛��A7�w�4�.]���s�Vay��nR?��՛��Ս����ۥZ  HUIDAT�]KچCs E��ƹm$C���6�a�g��i�)���'QGJ�v���åuڪ���;����v�G�a�b0�������^]�)�3j�ǨR%X2���[G:Ӝ=�u�����8�@#�.u}��J�c8�k�)o�(s�Y�gas�*	���n
�s���G��e�*N�N�Q����K�)�i*��	@��eʆ�	�0~����`��S��������,�O��g���\|�R�s�!sb�1^a����
&��5�W\��g8��zΊ�x=S��kع�F�N�7kͳ7=��f�Ju�F2��=h���5�L�"���Ŭ�e�w�4s��{܊���`��rnR�/j�s�v2��*ǣB3��ҋ�m(,l*��R���7�$�U�g���{}��������	G�L�w{��Н�{��U����z�aZFz'Y�9�������vWf*/'��?FYbx�F�|W�F�"�qzvz�Ү{��d����F��N�M��E�����he�;91��n�H�͕OQ�Q��k� ����=��<�ϣg���5�ǭ��'k̓+D�Q���������%/��t�SO?�l�
��I���^�~��$�v�}�`r���w��${f��2gf���~����B�+��o���W~�W��������(�q��a\E
D?&��G������q#�s��ݒubr��0d�anM��XLU�Z_��[OU��e%t
9��ءl���"��µ�a�|���Wv����{��w�����c4�җ�D���[��х.�Ʈ;��H��IbO�X�2Iݘ�a8�G�R��Y���2�C�/>�x��~�y���j��g��^�&�,�y���u���lR'J� %�XC��1��k�������v�2�l��2�9��BIwc�Y��w��H�FmXh���c�q6a��:vi�3���/��1I���Q���|tTNvW�Y:ųرL(�xX�U>�K�)Y��+N��v��`R�����8?�vn�k�k�u�`��>����Qϫ�Z���{���U�P�a9�Ŧ�Vb�_Fc�ퟎ1��������Jz�b��t��:�W��lךs�(7%2��8,a����T�rLI���ڟ5�}S6��s����-¤��#Y�1"n�1b	v��4��mj���q|��c����o�1�����|6y��{Z�m�����������ͣ�L�V�`aF����n�%�BN��B�9��� ��8=���ud��q6�r��>.q��=��x�s��S��)��ӡ{��2��J�,Isg���)����V~��"�#;�g�-y:���%7'K	^7��mSNe�ۻ���Pf��ȥ+��,-^M��5�,=�ه��P����q��%���dD�8n�N�7o�n>�y����2�떽i�sO\���n��I��5�FPE	ɱ�:�
�'u�ɧ�����o�ӥ����/���כ����6t!��UٹI�D���Ʌ��f��Hc��ް��4&!p�N���.��b��<q��Y���e��d����܃R.�PZ�jT���%C�2�������9m����4�Ce�h?�*����ߣ����L���"��%l�0J��B ���G�"7o�Bq,E�n{�u��)��d��4��ܿ���� �G�J2��KO�Y>�\�v�9�7��M�g�w��3of_k矽�w���X!Ң��� ��p��L#xْf��ϜXEvor���k�lO쟊����)>$����>�`�}l����¢]G���Q�J_3�s ���!?ϧ(1Ϟchu�ڔ���Tv�`�~�l�=�V#�����U� c�ǀ�qs������~2	�zi��-+��w��j��=*$"�ӯ�����Mw ���K�A\D8��C�� �~��t��ˡ��k�\�:]��Xt#���ꆸ���t#�_��:ls;F1) x�ܷ}�!�]�+>�9�_�|8:�U��NH5�s��r�=����:��l�%�ށsX(y�~.���EW%�$hp�H㮍C��{pww����� �!H���ڸ$�;�7�������թ�=���s�V�����Y����E]׎�@b�׊�]���xog5J���ߔ.��!��x��������<=�&�Ȕ���˅�u�MҘt�I���Į��_���n���n�\��)~�p�~:��2o_��w��s�<��"a�iv<E��kO*:^NoE�w��⾸g�F�`ҭ�
����U�a;I9aճ�G Kl�}M�S�5��ou�g�= �I4b�e�Mv��%���#�<�ȭ�
Q㺞}hQ�ԩT�0��f�Zn�x=��5�T��� v}ZǍ=~a'�<;�F �ɂ��7���� �*�`���Roj�NJW�Iz�W�x+�V:t�S��Nlj����⪝ ͚�m���ڙ��B�hL�.�儊PK܋���G�9{v~4�&{�3�ݸ4�:W��*�+�o��8ӋR����q6{�L��J���)Ͷ1B6��!���I��e[u�g�v�p	�J0�`��0E�JF�B梠��n�O�ȷ�o��"q����*�H����m�/*]֔����8$�u�j�=-��Ƈ��w��`���ˏ��q]b��I}yΩK�pJ[���<�/�$��_��E$;�aKN�-aKN��&��Drrrh�=�P���Nĺ�U$O�G+��Poq(PCŭ����Ϥ\6)#>n�K�0��1b%e/BW��U�4B�#��k"��e���+�.^�E���T����ާة?�6MZ�������㢶�I��3�m��'�;=N_���8?+����%���t�jcK���A�-��
IDC�]K��(7b�?�����~-��M�r8Hز�E�?�^O�ǹ�H��:w���y��S�Kн�5w_��W��H<E�g�=�x|����S����t�v[��şQ*/_K��D��(�~~�u0�����u�
�LFȰ"i��l��p����k�p��<�Eq"��;4�
nI�=,�(�qm��|$�L��!㽒� ��E���=��~t 9C*F�{�nOcCs%��L��\��|��h��2�(��J��g�J��mE��ց��h@g��;b�Jy <����-W���6�y5��A_殾�/�'-/n��������/��?-�a>,��H��X�����Z�5�	��c�w�fhkw�R_O��2�6�$���mʲ)�]�>���6�����]'���\����/�D=����Q�LD�&�����8��mG9މ{ަ�/��B~���|�f�
���uSc��w�k�@�q�N���&����e����Э��(�����71C<�� ������o����Asu����s�ߐ�-C�[�c�LG3R޶(��y�����H�~C=E|�}.q�w'v���6�n�-5a�QS�m�����������ƀ�K�GLB�<�˔��"�zף���w�����E��w��c�D/�Aa
����~9��6��?9K�G&�$�H��2I,��4��ծ%�c��{�R"�g�� �5�lfy�V)��59�Y9�w��A��1��1s���Y4Bu����F�\�-��FBt@��bz�֦�p����aZqy� �?�\�R�ꯌvwٶr*Lv�s��Ǌ(�ħ�4=W�8�j���K�$B�flٖ)t����0�*���L!5��W�w.� �i���V�X΀�{�\&%!�},�K�}���MX�B�駅R������>��.��K�Uw/�x���f������7�d���ͤ���l���ø�p��:ŔX��@���/�d��������;<�i�}���:m,��~a�.�H�����ox�������woA�����<�1ғ��Vγ=���>�L\�x!^�Ͷ�<�4�e-�2(│�����?v�a;+����Xt����Jç	]�H�l�&��q�͛����@Z����[;X��KS���������Y��@�D�'���!v�M������#7H�������<��\�����{�J|�������6L͡�������-���E�KjC�g�A��V0E�oc�ݍS��>�Dx��{� =*l���kd1���A����D�>�u�+>�͗�ud?��=�[$��d`�4�U��Cy|�%���$?��Rr�8uXDޣ����k�"O�a�"��`d{|UX��4�����T)��vCO��{�Qf�Z\t�WJ���q�*I|�򟍸h	���_�~�����%\����})�Ϟ(�bqsB^���	����J��s�R����M3����ޕ�׋r�����V�L��zʄ��Ϧ�ĸ_��"a��<��o@�v��ߵgu;�L2k�c��n^>�(����S���N�"�}6�?�������f�ݚ�?��H�PSf՗�k���Z�W_(���W���>�i$�M/dA=�����	;���O784�H0��t���8�"q���#�Z�ʐ�1�F�E�^�R��)�����:�Nh1����ۚ��}&�֚
��0��ڋ��R\E��ܞ�h��y;/yZ��X�N��L蜤=����.�8�FJe��d~�}��&H����7ZGϏ��/��uX������v�&f���Qwn)�^0��w������	5�5�4ٱ������vV����^M��1rظ!gQ2ć�A��h�d��'��d��r@��W�����V7�i��c�(�,������橷��j�x�<�a��_t�E	���>�&�82���ܚ��R.+̳��8Vɾ��?IH�^_X���Ą��]��;��V�%4�4'��٥�S����d���
��I	Y���(2t�� �Y���A:sp8[��?N�zs2��/�E?l�Q��srS���?@JϢH���S���pC�U�36�e�����I��%��+j�XJ>�)C�5!Y����}SQ��nA��s��T��L=��`�3����1^��A��)���-}��"Y
����b����Z�nz�+k�DB:#v	ݓ����r)��P�����0��.Hc�Yu���S>4�W��5�$$�;i�J�Y���ß�&1'��B�Z6M��T��?Q�Z	��yE��0Mk��4l��=�V�ߎZ�з�cu�-�3�HbC3����ihB���d&���	�(��w�g����,�?�O> �v�E1(�#q������R��J�?!-X�Ǻ�o �l7߶U��=�H��]�ϛީ���2yP3@p����:z���Yч"�@̬Pz����|I9P��bvFԢL���c�H]�)M�Uq���_��y`��.�i�#]^X�[�*��V��eh�BEn��[!���SY5~�j\	�v���.l�,Mk��>_F�ګ��8�<���8� R<e���bC5@�t��ň����|xa�CdS'��-��5���q�Z�x�=��u�w�#F#�w�fp��ߢ0��i�z���f��]Z~�s{p�e��pou����F"8��CT[�5�����'=��WJ�9�*��h�l�~��BD��G/����-ŝ��D��=jX_iD)��;SW�bt%��2�l�.�_�"S���c4�uJ������إ��v�Ć2�lW���1.L>L�:�l̪P�%����@�/�US/A�1�%0D���	Ks�^����AI/#��U.r��v�=�N�����>�Q	��k��4L��-�w9q���9QfŇcg[no�Έ������U&�rm�lə���9y ؇j4��(�oY���Q�y��kŌp�+���B{�����C��q �� .�K�"����6*I�Z����[�ka�W�^��W��7E_��r����?�m���|y���8�>����no��O�%?#�l�u����6!?�k���!��[�e���438��Y(+]Q�9ñ~C=�௜�#.��p�o�/Y`�3��4z����,�o��nBT���4֙���?��B�Oa	�2T�pL���Q�F��~x���凜�+���&�'@��-�I�D®I�B�I�D���Iq���X��@zy6�G�W2L�~x�V$8'�v�?�쐪XB�#|��︧��KB�OI5�0(96P�ϼ0�c�3{��rj��<Ve���!S�RW���;|�&{�, ������@Sr�)��[(2o��&��w��_BdzH���k�j*2^	
n����?�A���	�������7{_�O(����k��J�@]g�����I|�� 4�u6����'�D��G~u�.�L`���3=�>>����r[pH���5�&�X3�ծ�=��A=p?yza����g��ח\��b�kw�}"ל�<ɞ��aMK���o0N��ϣ�.M��������#�.D�i��r��	���{�\�������゘ݯlx&��	���D����Ͳ�s3��T���EF��	W<�e���#5����c��[|��+߹[���#%Rm'y� ��I�ci�s����b|ܽո�5N1�*v��i��p4�������ƌp`�wyʹ+��ʒ���'4��۩���m*�+S�C�$��b�B�k�}��3Ơ���S��ϙ����N\)Jq���.�^�`$��Lwx^�_tŪ,����TJ�&˖�G��G��C������v����#����դ�-��kQ�ךy�A�$��N���N>�\���gwQ�&��k�8@W+�ػl�'�X��	��Kb;^oL��͹8eo�ocg:��c�ϑI��
d>�8hRDH;���$��{�o��9�<��Ta��p�)����������1�k�k��U�	!0�H�3 �3L�&��#�F�3o|���'���W����,.0bK���ҡ�OO\}#��F޷���,҇���F�Q���j����9�����eM���=�{;w�+b�;F�ht��&��
D�<�'N�e��j^Vk��ؿ�lw���q[*���.L8�[��]/t�-}��Sl`C�U�Sz̡7���<�;��O>nJmc��	���
ϳ	�&�T��2f�JH^=��w��:bj��V�����[ɌC�����Lk ��~�.1.�r�h�G#�Cg�	12|/�@�� )ة�]U��'s���>���y%V0mrm`އ��	�	��M7�6��u ��R�r������}�⯍�1�<�	 b�f��Ŕ�����P�Q�-vr��iذ
�d5�nɏvb��^2���Q���''Zہ;-���OO7t����@=�q��t(W�;�j�����	�� a�phDHEjl��"��_�G���;�!�ҊnzAh���@
�<iH"����Mn���s綌�B�?�R�э�$��=)�r�/�㙮��;¸x�e�[]c�D"��4����Pթ�}J�'�qYN,���$fߣJмD$�r�%JӶi���zH%�ē�$�e�к(JW�ݩ��(?�Z[�P��R���y�$�f��3��a[�?��_ŵ�)[����ET�����_���\�C���
H_Ie��ֿa�Ji�����D6��I�mQ�m���rgM�=�)���	/6?ӄS8$ES��U�V�D�Ub���V&n�p1.�wxaP�+��,s�$��o^k��hBf/��"����M���!�5��O�l��	�j-���C�bҾȪ�s#���S�~��j��I��_8��uXPζpDYG��!�RFvKO���B�S��P�)�=Ձ��(Jиm'���iC9z��W�!V�vR^h91�zC�A��Vvj�V��/�7�!5������?��Y`Ʊ�3�\@�u霠(n��	�%�05?mǒm�w���|HF凭��i�m��Hu����2���{m�i!m�R����Ũ/ %a/@�G����A�T@��c����/��:��5ޗ��v�5���䝯�\^k��CWG\-�u6����7Q:B$E�x��,s�6��Gו�J�9zwX$$�A�ɥ��>��W]p��)��Q�)i%Qض��GG@paA��u�q�P�'��%`�9ٯTń���%�P��!�ݠ�(�~h7�
��SY8�,��}.��Y�e\-��{���M!8yb.��uƈ�p�z=@�Y��f,�R�&d@�A�E������v ~������)�u��+t���R��.9���+�$�M|j���-���`��a������k%t��;��Z*�8��5B)|Uh��ӕ�xM��?�(��aM$u6�����*�C��6�'�V�E�a�<�`�R�E�X�D���?!����R�[��b㎤ܔ�I��]3<�y������8�(�����大��c߂��il'M>��S�����5H�t�%��Cg���P��#����e.�\mJƏe��]&�gF�$4��Q���O�(�`����*h5ص �gt�Yr��X��XvnEk�rz�yW�\�P�/�G^��#���1�Y����N��;�OG2hUǬ��i�Ձ+��E�۟��]�`�R}��9�sgL�//�>.'��*ċG�1S�T�<5���F-�C^'��oF֧u�1ǥ��"L,���u�|H5sNI��� ]���P�<8=��<��ŗV�,3>���~�_
���{�!�g�)�ݬ�БIRLI��U�pĆ���@�鵯���Za��X'NǥUJ����O�]�r��Ai�2>��s�WJ*O��=v��0�oF����\�F!~�E�-�5I��*��ֿ�nK;vn�{�G�����[����*c�̢��|�ΰ�)R�[9 ��)z��|�k�a�Uy��.g{�;l�`>�T��vM����4z߿�g�/���7&%���r�_��U����M��c_p�E�Ǵ�I&���G�Im�WmϹ�b*&�	�P��Wʤ�'8u��
2@K?���]׃Uޢ�2+��q���2�k�!=a,��F���ut��OIvH>(����}�Nd���~&���I�Ęs�e��4�u��m�Y
mZ�}(n���)ީ�	�A���0ԯ�H0ZNUj��P[�V��ǣmd�:&ݡgC@�l��(�?�UT��[/���2GH��3/6���&�����;O�p��
�y���/2�싚CZ3s�u�M�?�d%�t�8��O��Mw�m�%��t|�,R?��FIA�8��_9�����dJ���a�v[#x��Ώ�u�*���U�9���I	x!	�f�ʩ�z�h�'��.���Hwr��� iD�<=����?��J9�i�����t]U��S�� UK�K��T件R8TE2O~�'�3
r��I���>$�V'��^;1!C�EY�Ƶj��c�ڽo��%��S�RhF�*e��t�Ŋ�����A�W��`�A���!���5���:+��h�~�!����ۛ~�Q���� �c)�`���3Č�S���_Ҍ�
���µҖE��e3(����^�6A��s��7�-�~z�B�W8^MLѻ�R*5y�07'#���s�*�9d��Aa���E�����U�xs��&�3�`�WE�����B<����]� �=��SE*.��K%��?��0GV���XmS�♪��%���
w瞉�AT������� �<�V�}VN��bDm��l�F۬8�����S5֛��7��T*qC����+��n�5
_X�^��f�&"=ҩ!P���gG����jl����M��c��a^�j���}s�sf-���l��̽��w� I�7rM���^m�/���x��#!�t���:�ˌ�Zǚw�xy�7��K�UnI����~��� 0�0�|/N��\e�vE�θ�-�:�)L�K���z4�=�5J�d��n�FxN��T�x!E��H��7ܟk��	���K�߰G�d�D
�;҇���⟥�aV�!��>�PJ@�����]=_Fy�vC�eD�.�5�,��DKq��GG�m��aQ�MR;#bfY��s"̳��=�b||�<�{'A�g�;*Kr+;ZR&>9lZ�
�Z�b�%:d�-=������c`"�,�{@9�:���1{��_�{P\{D2��2����ۂh+6PvI
�$YB�8��:��T�/�p�/�l2��A#��������.���-��c��^�E�}{���m]'k45�!fS2�О(���9���t��M�	&�ӊ� X:��%��<w�Z��*�JYJIL��rg ���Coŋ鲔��o
f����Dkld���Ҫyo�~JW��1[Y�[x?MêOl�oG���T�%��f�JUTP;��L >`�~����&R:�X ��~p����ǕeT&B��g�ѯ�ҫ	Ĳ�B��bB�b�xlNE9��pEͽ���eW��B�$�a\&X��휂��t~�^��uGBأ���'�M����_·�;���D�G�g�\i�\,��,h���*�1۵\LqW�ٷbn�z��3ԋ1�t�o��Jg�Pn���pŀ�A_J��1�.�q�}�$z�]k����ɧ�Z��!�`�$�1&͚�O�Q@���ƫ��I�+7��cvߤ�g��S�
�/�ye=�$��7wa�$!�UU)�?��[��j�_z��b=��\2�<�����MϺ�ӥM,�dO�x���x~�ʞa�N���=���L�ƝY��TU�#>Z��ä�\���;l����3������_�U������uZ���Zy@��w˅ǿ=�M+!\��O}FV?���[��k<����Ja:�p�����0�� ~Wt�{v#������l��&X���,�x�<�7��B89�Dm_�Y�$���k��'Ĳ��<�'6H������Ǡ���{��z;s�´�ρ~*΄]���O�isc��?�׺��A��A���	�e���ۓ-Ҷ�}}�Ž_��=��j(�AK-ܹO��?�=Yٿj!'��n7�>'E��6�e�!B%�V�B>[�:���������J���20cX+�>���hpXE��k('��!f���a6�m?��U�U�M�ww��W����C�G@�k�Rhɘ��T��-�ac-`e�-f$���-�4��)���FM�/V�!�g��"M���1��K���6f��L��ƾ���BWڛuA0��5��mqjy�;у�>��7�������TWryգؗ�|oA'�d�9�["ԟڱ�sс���)���1�B:�%D0	�㠈���� �tL�̒n�P>7'@O�<s|����чo��~t0P���-`
#�'ۭ乲)8?��^�<����������_�y��o.3u7=%��7��أ:`��X������L�d��lS�;j,K�ʴ+bZI$��>�3�p������]�����9;۫�ù$�`z�k���O?<[c͐S�1���<MQ�}gH�Np��m�/��CV-�ח��?U6��,����Zx�縿��F�uk1� �\>�u$l*e���pC�=�=�2|tv�e��7zn�;�L:�g�2��S޻�``��V�WNY��$ޘ���V����j��(���6d%�ك��:I`kx�EL�ڸ/ȈF�������X�gF�KU�1��SE�t��z��b�bg39T^9����&&����G"� =�xc-d�2qrz�ӳ�[GG�}~��ȭPU��7�T�䅒q����bJ��8�?�in�C�W�p����u�,�/"���g0D�
�2�9�D�b�~R6�#L- |7�����c�Ym�l8h���x�tm�*QL_�M�u�M�)["����VIwğ����N슓�b����&��'�)p�ld���Nd�J�^������#�Y��<��7���
6�+G_0g��t�I4	g�홁F�'#�2�2T:Л�k���G��v#!Zd�+Χ�_Ґ �oc[�GМ'��g��_���z$��E��L�F��`��i�.�!�c��%����g�O0���k��f<�b�\��X�ڗϸ�)�I��BE���Ō�(%��й���7-�Qv�]��M7;��Bަ���{�"�$-��&�}���˫+y����$<�:%_��
�zξt�:��<��,5~Y�����+3>��1�J$T�6 ���m¨�>�J&x��y@Ȥq�haQڎR}��я�;��{�g�������"�i7B����`O���z��mp��TKl#��vO9)�ʿQ�w2�#ya"wC����D�
TI
pQ>x���-XV�=��!��x��R��j/�H,�U=�2B�e��v]n���K9�yrLƠ0�9�E`q�Pǿ����AZn&KX;��?��˦3�?��\�5R[�OeMe���øH4��/�=@1ܚ X�,�y�]�~�5�T����2!qG�xx	v$���ڒ_z2���^ϰ�=���v�Xۓ�����R�Z�e#�*͊���*�����w�>��(DpBB@y���g�3�Y��^�t�X0���)7W��v;�%���e��h�BIr=�����KH�$��_�݉.��ˈ�������O-{R~��y��5Et�푗lG�K���o?��-ɀDd�Łl�]� ��	�l���X7��5����jZ*�N�GϤ�9�/O7ς��P\ݿ: .[�����Bq	D�d�`x����u�������p	v��"�?g[�͇�3YHh&���ښ��P�:,8����*��$���OD�g�Y�|������r�NBU���޿����(�rC��{���S)�ܝ��l�����C��Ś��i��zk*�<C/�&��$�z�r�Th��E��W>��V^�r�;z+�޷h��`� �%L�ZL���|�ߡI�B++�Y���Վ�,BwJ���x`���XI��c��0a6};#�Ժ�)��Xt��'��9��c =S�{1׷8��m�@)����X�i��c� /���)*�n��ZM{�Wd�iI{\6¡�n�����@�=3G2S�A��_O?�ș�O�s�f��".�K�]�Kٴ�R����)<�~�VK��.�U�h?ݾ��j"��%���â��YV.��j �%��d�����Z2��'f-�7�� ;�/��RRd۽�+`_�d�"��O_��A۵�]��|��e:̂�f�sᴚ�
���&8LϠu��+��ו�����[��`"�����U�p��-v����Т]����۫�0��ţ�K��\$��L8x�o?xeY靟I���H�-y��1�7���ˏy0����X�,�[cC#��O������*Y�^�V�L��I[�J�d���i�vEl	�)k>3���f]K_7���Ȳ&d�1��� ����=��\؋\���|���$�y���K����4Ǣ�x�B�:�G�z�A��A���H�������>�Wf���*d&����}�z�杯���q|2���d�-IWQ�vU������W�b��J�,`S�*Yf�d��M7�h#�y�6�/��J[e։i�9</�1*9��*)ED��H(���P�UBa��VTUT��{��n8���ԘIQk��&���VC�O��;���߲� ���RNFI��FLm���0����jw�{����*���5X������(��^�i6�d-v)	���Ӧ���e���2�r��$)|�����5�_�q �4�hZJ��u��.f�&}��"O��m�
�� k�`u���T����F�"YcJ;�&_v�I/u?CTs�Y2Ӹ�㾬�q/˅p�`��Z@eD���Z��.���/a
w�*�n"�d�}���"Ms�9�kk��L��2'r�M殕���#�ᇶ�t�?F�g���)eU���*!��3,��cL����X	KY��!Іs�*������C����֔��Ѽ¶��5�s�%��T�"ՙdZ�oq(C�c�y��X,�壙7h��<x�WJx��R��MyY�+^��Y,��H!�����S1u\(�4*o�t�f�Z�	K�[ˌn����L�Y���Ng?����"����5"M�x��%9�8�N�����I���gZj�f6R�tE��f΅~e�y���	L!qЕA�r,��㫘�2�Ҷ(H!G�y�����E�VzlQL�i��?=�g�66���HJ9X-��d�+���Q&,����|��&H�����(&3�5��df�ݷI�%Ϭ��bA{�ï�^�)\�S�=��3����ѪI�hH�e����凿�*`Y#��'�:�\�R�u��N%=Ѿ.��W�0�L	T���D��P%m(��N�C�(0����s)=b�7$*)��g�c+�^�v
��Bh6�����$�?����X�s�p��ꪓ�r�cś�k�tշ�������gi�A��/ro&6Ȣ�����j��;�[�����`mx��1[�b��D�B�����-��&V�S�G�{��
9$�#J���?.5��w\8֮H�^.��m�%�)�,+c>���W�kf�f�m�3��4�R9y=(�y1%����m�y��k:-R���2�]Q���l[�*�*�r�T�Ϻ(�����ܠ>GP�K`���O�|
w9��E�ў��*�E�M�����US��fT���o�0�rm	l��jzR^F3���c�����_I��B�]���5G�4�Rpq��|�.y-�#�h!��ṳ7���Lf�k�p�ρ;�+b�������������8D���ڕ2{��e��ۓ�x���:�mֿ�"!�� ��1����mc�,��;|�Rd}N�)+��C	>$	3�t�|��MD�̶�]��Ă��"�`;Sf;R�u��%��<��cm|a����x�	aݮ'a���9&�SJyf�ڪ��ʯ��q ��4�k��}ה��x5;���r�U�}��1�h�Lx|���H+Jt���h��w6��AH������s�|4}w`�h����|v�q,��hY�q�P{2�HYe&w��~9U�0�L64 �Y��/@�؄���S�"���H��j����"ԉ?��vIw�Oj�!��9��,�M֣�\�\ץ3�m�kb���)R4��Nd�z�Y�Wju����5)��C��m�8{Cw�5�xSl�r
_3�KP��D���qH���XƆًu�q�¥fQǕ$�����������t���g,���^���/O��}�`u=$nb?&�V��<���WnG*�vW�mMCav^6H�*�ƒ��%��C��k���=�\�@��Bs�eQ����V��9x�#Yٟ��m��9�DHPv_m��߱N��51�'�,��CP���$�>��C����Ur���ݎ]���Ӷ��K��[�:q�:}UA!�Θ��h,����'7��4se�I/d��x.!��[��#�SR���l�rGR6�:���_��⼒nt�3-�-��z�'(2���5�O�獏��h_]�^!��*�1�������:�����;�sn#��/$v7���2�Q��h͛��}�du�����WY��w�p���	j�nB����-�ȵ���?謨��G��bn��i�-U��o���إ�iK�Gj�{	�4TD�1X�w6`2T��1'tO��Vx�ȘZ����1ĺ�L?�1,���
��鳷WN?��t������R�+,IYZ6�� %ˡ�ǾPj�v�:�Ǚ.sd���~W��pޤ��g��I��g���J�u,�!a�qB��I����l%�8G��{�����.��k*��$n4�7'�V\�M��B�P���2P�
�=�S��֧@*띘�޻���-��$��.O��ץ<�;��VUS�	����3��"�Pg������5�^r`���F��y�����>牣��4:��]�Y�Y���S�\롪��I��"U��F!攴6�9,��T�����0�����{J}NO!�'c7O��f�Ի\Q^��Ԉ%K���{��6�?�~f�wR8U��xv��1�s1��H*�[6T�H��B�Ew�A��㐳�������i`�>��3f��%�ȁ�;L�wM>����������l�k�����2��"�Z�𿑑TW��PK   �u�X	�\  \  /   images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.png�W�W��%����K`鮥;%����n��I�EV� !݋�t�>��;�̝{��qft�U𰩱  ���"��:��&�ߔ���'X^���  ���q1��w��S2���t���y�s�p��z����T�|M ��)���YfO�����~qv��ّ��v�C�m��� 91��3�,.���3��2м�P%sVOV����$�\09�U,��Ka�����fv�6{{l����c}uu�ڻ����\"�4����h�v�Y�!^����!7�)�Nʑ��[��������y�B�{rrr/[��q�$�|g�Q\P\�_��m����?���Z�|�}�X__�-��pM���������O{uNF����0M8�W-�Դ��۱�茀��4�7�/c���'ˎ�{ƀ������ka��r-�v����}|/}||4�y}>~�w�R1)d�-�uYvW��������kkkW�O��V.nn�� ��|'��I����K$A~���:���0/�j�ڍ>�^�,��ۛ���x��krΖ[�2��������I����}b�t�#���3jL�Tp�f���%�M��&g>���h����Ŝ#)}V�c}pr`�A�W�rm('���� � ���0���7, ZB��{����p_�u~�>55��ŗ�L7u��aMH����euU�򢻋�@q19n�ViFq�{$'��Q2��SGv�< ���Z3?d(9_�S���'���Jߧ�kc���h���dNF��1�;U{�K�����B�~�o��JL��S�d���b��*��+f`uy��[!s^���w����%]�sCã�~�����������x� �r�fr+�T�^����>uMֵ�컁1t���!��Y*��%p�fWD�����Auu�]��E�R999�e���R���M뭡��'�i�=N�#U�LԾ��<�ۯ���g~��d,x�>�-�&Inv]_���]����*V �|�������B��.{��,s5��D���#��Y�]��f�h,�2�@������?@=Y-���犸��{ǦvFϵ{�����eI��<�T�ۮ�?�=����#D@c]�!��Wg�>6���g�T��Tnƻ;� x��ú�(���F�����.Y����֞N�;=��U�v#�Q�EA��� ���o����T�����<�]Ц���P�U�X殎1��ٽ���ş��z��ɿ�eN�]�jGs���\{{�0W�5(���f��,4��S*��A� sIh��Nw2�J�l�ਜ਼��X�2h��3x��%Ǩ�j�L����	!Y�@�G�s��*�l���#�ie�	IM�f�� �����W��D�����<;a�+~"�
z��;B�t�U�ť�&֗ff�1ɭ�}q��2JZ����vj�6q�^ c�Ì�M���(�0E�⇥�<���-��~ �*�塈(-�?���Ć��$??���q�yr!Y��:�	�7�M��m��;e |F]Z0�u��Ӿj\pW()I�+)�F�8epr/a'?�޳����]_А��Y�5�����ff��Eig������G��i�	��7?���y���yVq�]�x����
��1�fs�(�/�s��l�R:-���^(��6?�s���N?���eu�-�&�i�czkH��Q]��"uj�Fz�0��a��5�f�H�EK���c/I{k`��pG��ߥ=n��[����ڥ.w�p�a�a*h4�Vb%F�J�觍��vgc����<n�����a��eG����U���A�5��֊	w)��~��+����i�f��uaΚ�¯��k����[ ��陙�.`ra�AlqC�h����6�S��'i���nSo�'�$���ٹ����WKF~�!��%�0d\��Em�O]䃍��+��qLi�\���k>
;|P��&�Q6P40L:G����J7>0�e+��f�Ԡ���,��{*�$��Q��$h��#��~�i��*	:�R=�0O�!�������d�!8�۠( 4����U��-�l*�L�� ����\���ch�*���bh�J؆*�m K�1��JM;���s��¢k=�{�5���l^6�&cW4|Y}}wl��j�i{�y������Q�S
�	�Jk����rl(@�%ݴ'm�ڕm~�����=�tLV��%0#)��{C��@Z3��h`��[�0$/x�t ��g�?�H�!�B�tV�+61��BG�nna�R���o�^2�J����+�Oic6|������$��,�8`��~K��	K������儃��{(������v�>�)�����'�ςE�\���udJ�HG����5�ؑ\J�M���M����D[���#y���� طt.����Z������C�+[�H�����nK!IG~\���@�#.f[��=�-�#�=	�k�T����B-�m�7��p�������'��9BL�[Xvل��Ԥ0��L�;,K��Rd�n��5���,�J2^�A�+*RR�����g���U�)��ݗU4�����s�c������Fۦ`e�m6vX�t����V��X7��������F�M���1��7?tK�z+~>�\�鑵z���.���il0Ͷ��z�����o�j���W�)���d6p�n��X�����5D���'�((���W�_��r�wu�5��b��ߏ�7{4����۔iA2�x	O��o�ͩr�Alȅ��o��)�?�P���/J��(��)>�-��qQ֒7�������q��a$��7�N#&msܪ��/pѱ3���H굪F�H%n�58��G̮��*�'B�87�����%n�p!=ExC���'�'�F�+�,�2���(w�Q���Y�� Y�XO�Y;�2�����dI/#|�%��z�0%%��=J������8��]�@y�? gnd�ns��O���kI�dv�E���E�/%����@���q�L}@N?:D���,lJ�#˩��fh7zC���[��K�1Æ�5��Y��5�UEd��{V �8�f͙��:P�h9_���%\�}����7�E�P�E���E��1D;I�8}��rO�C��\�&�Z������8{3ͭ�M&ވ
 p�����4�BtuP'^
��/�Q���[�$���%��U7��Ĕ����v�����Z���*�\�W�U���gj���=}���D�hR#��E0��fi�ۑ��>5eY���3viܵ�e�����hA�v\z��7���r؇�ҭM�iPP6ֳ}��=����u����!x/�E�`�%��c�<���,G��
7Ŵl3���}S�A�:1��	�p�����_�ð5=߉|Xj�W-G4�Ҧ4�����[�8���UP@����m}M*�Q�CQ�{�nK+hb�M��զ�Z{m���JM�W���1���7����h��PO��)�y�~�6�{�$U��F 3��U_���h �=�������l_G�R*�MF)'<���H�~V��BI��vp�66.�+up�nf�p�y��ˬ�������%��#Ҿ��� *b?0r�p )�ʮ_FCg�^�u�NkRa�lI5�x@�	Ub?)�Y�����𷌌z�|�<04�'�m�r%h?�c�;�_O��Q��I�F��bW��9`&aL�8�S�I)�P��M�~3���Kx����ދ���2���qc��)v���4Z�p�o��I��	�jk���4��V����V6��2@:\WD�5F%�D��o��پM��g�\�!��@�����[�Qxa��F]����/���mA�zl tG[r,?ɳ��h|f�C�f�xgW���tg���	Q�!� ����<�2���
��S�����uʫ�H�1c ��$7ے�]9iJ%��K��x|H��?�u�R��䥏�~�ꄍ������p..�Y�ܬ�ܨpS{�!N����� ^g5K��;U�|0�.~\�p��Y-8/�ة�{^|�1��жٟ�Z:k�2rc���yrS���\�M�A�ǭu��w{ۗ�)���濆���w��Xw�/��}��6�'�Z
��b�!�|��լ8#��;�o7���i��I[�P}����Ę�-���;ɵ��,�E.r���aUț��j���}9$���LZ��N�����Sw�웩N^7+Q�ZrDoo�n&���.G1`��8C�
�v�Rl~Yk���J?:>F JM=߹5���%��'ב�pB�U����V��Q���&3��]M}��L�؁����Ц@q%���v���ߵ�y$Ϥ w� ��?��unin��}�[C�y���a	t³�{�}�^���T�U74L-��9�U#��!`ƕ4:� fPpF����v�N��z$9�;q9���cO����{�m?Z۬.j���Fw�*�6��k ��A�R  ��N�2Ͱmz�����B�?7&&��g�Q7��p�%Q�p��*��۹M�[.ԉ�xKK�s�4����e��".�1* �0A�Yc2�PH(i6D�w�`bQ eZ�:�tb�y9%<�	, �b�����C��+�a���&ղ����;[K�������`����E	�sy֝�w��E��W���������̃VެGG�S��tך��X�����،�����)�U�<��x���~�ݹ�l��{Sj�w�)�ƺ�a���k������y`eQ΁r^��;J��r�2m�慗B�OQ9%$�&Yj���C��̪0�[�E�^l�k��Y���/'�O@mILdw��h�7�܉2���c��_q�������1c����~��#nY�JB��g&jfE�rP+�" bzC�Øp��x]�U��� �I�����gN�@X�5`/9�䊌,�&��>�<p��s�ǆ���zu�k@���9N�v�o��=�	��y�Z�k�.�>Q���+	�R��igF�̚��T�Ǟ	����<D��7w���vUk��ٔ����*�'��'L�.��-�� q[PV���eOǻ�W�q˒0P������sۢ�V�SY�n"�T�N4@�y�M�ܟi��{f�=E�}|��_��#��2����W/4oT���=B�`H�֙�ɚ��JS:Ed�!e�%`��n���q�v\.��p�p��]�l�(��"�J\𘵾V�v�m��g�B5>�w�'�%� ^p
q�nބx��+��>�f������k�Wj��|��j���o��_�ʈ{K`"��vZ�,�[����=*w��Y�R������i���
��[˵��ж����,�"8�s/�(a���M��;�?Zr7(l��U� � 5<��N5�?�Zxn���~Rx�$}I,�OYQ(���8�-�z^��-$�W������0cg���Z�	ȋ�)��R�dA=͸���z������Y�\�+zl���y��8Ϻ�q�=�����6:8m�R��N���`-�J|�����,��!V#>N��Oq�g_�"t�uU���hX7o�m�i�Rr,L��z�->�#8ÀU�#�	6�s���Q69��&��w~�4�~���VC���� "�����y\U��j(�S�����Σ�Z�X�k�O	�!�$�~Q��X5�fѐ���,�4�#u]�1N�.8F=�Пux���|���(��:'�/C��[<�AVĐ!�j����˧��1���:�
�]�}1��L9�?eۼ2K����l�vr:��{��_�3I�p��P���fۼ	O����(a����w��r������̒I|=�����|K���'wJ1OU�#�AT?�^
q.b���\�kr���͸洘�%�Ct3˨��A�|ؕ��`�� �~�Τ$�-�'[
iXS���J;c�wso�H�=�
�w�HKP�~�^:=�!���B��3'�z��G����Oʑ=<!?]`;
�6�������H�&��5U��,/���P�}��մڢ
3V���\[@�e	O��i̝�KBm]�V9�}22�)�u1z��I���B66)X&�ր��1n ���Ph�ĉ��ۘ���BG�AAa��S}}ɯ�*��I��z���C�;i�F�DV�O�	�GV6F�2<��v�����'�/qK�E(�Wኬ��b>��Jbd<���T<�VJJJis]]p�R���SM����3�rW�����BF���7��!�����x����!w@=l̺�㮌c��*3��ڂ�L�/��"U`�*_�!��?��^�S?�z���I�^E��[�ןb��R�G#��ݎ�]���z@�������]ϣ[Cگ,��j=���j����4ݗ=��ڱ��Tu�:$sy�ab���0d��1�L ����G����5�>9�iزiK�VFQ�f���u��?FSS���X^s��Ja:���?QY�����]ǁ�%��[����n�t���>cd�n���5��e�#n�{~co׼�X�LJ���%��2���W�`�ee*���K0Ȭ��RX}	y�q��/����(���L.,~�{�r�*�Ţh�H@n=w�-�˄M�8�sũ
�Z�1����sqw��5?�mVYuz>��7P\�?5�*l���R���"�<=�j�"���3��ՙ����-$ ����I�7n���b���1g$���i�����9���L/��q�#������&�FFJz3�U(SR�S��y�.��@*�'Q1���X]�./��f*�����'��$::��Q}kY�u!>K��~�K��z6x��0晀k�˻:ݴ�+#x+A�`w7�s�dm��q/ɵ����\�ig �ִZ�$���H)���Hd�g��u��#�.����[S"��u:�
8��k5Б�~�(4�}��iM#�����32y5r�`K���\c���׍���g,�d���qJ(�HDKR�Wuk�WY�
�ym�fg�ؒǽ2SI)W����qȮԒ����+�ϡ�36ZB�!B��V�	�(�dϓ�S�,�g�����g�Ih�Hx��Ȟ��|�b��.8x������+\b��O�	������_�K9f�Ð��n��T-�w�s�Ǻ�奯O�F�e3^�����"X���/)7�z
l�50v^���f� �T��剡��O�Z�'�jJڊM�6Q�PK   �cW�����8 �I /   images/996ffe1e-7752-4112-9b94-ba61923e6aca.png���7����D�D��D��	�k�{�u�!D�-z�h���3��� �`�2�6��w���'\�~�΃s�s�{���k�=U�GL����(�Ք������H����/���!qQR�SWR����rtqw��*������#|MDN���N�X�M���#*�(j���d��z-r�
�Տ#�,��!@P)�zO���\N������-rI���"����{�ȥw���
���j�St����?����-��KV�� �O�w?�Prd��:��z;y?�f/}�!�4&"�%%i,�%'_5cdx��9`H'(x�&(�.�J���h���c�����Y9>'�d{kꮞ���d$,�x H!';	�ї�}Գ"�`�Q��l�h�h�hF��yyU�=<|<<ueE� �#�S��I�z���uut����C��<����ԋ'�{�@#b��Z�p��Qq����B�s���\�UhW����+1���s�����G\�DE`/k''sB'�Bέp-F;���������?������?�?�DW�{�H����?q�Q���E�������@z�"��iuu~�Ԕqf��!�G�C�f�¨��"G�*ٍ�@  d&
��� ��:V^^���5�c���$d)��4���Ǯ���(�Kuh�ּ��s�1�l����}���l�^GM��X�媄v��� w�u����A��c�W6IB�`l�
����됭����@��!D���C��_�� ʹ w����heeX�16.Kd�`���ް���p�����Y����/\�l���D���oR-�v�����n�UO���*��X�#vܭ�(� \ɥ�b��X_�/�ǃ��ސ����wm�'��
%�� Pc�kD��K�Z8�L�{�xK���TA�Yhy8Eq}qSr�vX�Ⱥ&}y���M<���o�����=����$�V����@08���Jw�a�-g)D�Ep� �J$e{|������к�yբ� /;�M'�@�ATx�$��J�Ww�(���:X��T����+ޑr��xa-R��4t^#s������F�ӆ���>%}�mMkP�p�|w}�ݟ�ӯ�|H���U"�
��iQPa(����sQlvaW�u�� #���U��11�iDêۊy����L�]����ς�w�j���U;���:{�U�nA. ED�@7�쓌���?�NR#]�=�_����-bKB��WD�2���2�-�Sx��ۻ�*Ȯ {�1�k�nHׇ��W�v9
o�f61�聙K��e �bn�nvxX=�æ|Uy\���_�MҭH@ DD�3byx�O�hBT���C#{U�S|����̋����f��ZL������{ҋ�s�DE���������:U�"X����04��M`.i�Z��|�_Sb{A/��i\{8s��QM��:åCJ��T��I���x~�2(��l�E��'E��������ದ:�4U�y���ޱ#����BK���1��1�,{%�?H�k�#;�b���p�	g��x~A�T񢡓Z����ݹȻI� m^�lsa\[�-ιN@ԩx�{Qƀ.>X5��_2sⓟ���MU�6޼���c ���e?�	��z��O�g$����f^�s�C��R~��28E����B�����=��;Lt�G�>��M�l��;�uI`0B�����/�W�~S���$�)���5X>�����!J�%d��]��K��!��ՈV82=`�ז� �\�^UѪl���ۻfw��wtd'�2&�R㐽�1Z��3v��U���
@�n���]p���>�������j�&���F����Ǧ���O�>�������TJD˯�[�6*)�O���'QV֍�27�д�)QR(������݀-��8�s�1s؉Xq�9	�j9 ���#�ww�b�8�	�_l"؞�4.�~��d���Zt�X�����:�&�����Q?�>b�u�bV#`8kl��KR�q���Z|�֒~���f��=������!�3�'-�ӡC)��D<jo�����ǵ�0�������[Ug��7�;|��w��L����c�a�dd�܏E܇{9�9�Y��}B��7fF�z�YY�O�y��Ԟл���U)d`��O=L�:��Y��b���G�L��xN�K�������)������ӹ5�n��V����30�i�����2����J�%�J�Y$�rjq����z����ɳm����9ttt�}��x�i/x��KE֣{aR����3���r���h�*Xު�M��&uE@�V�iD\�HѾ.�܁Qfc}��.��O`)k����n�I-t��p@�pE�xW��)�Y|[X����ѭ,�ꔨk0߷�>$$t8���	�����m:����Ί��IA��?�"��3��h��ٶ�&�^-��k�����AS^�s{�������]�9H{����s��gӅ~�����W��[
�[Z��[I��;�h����#�]�m�Ϗ�Ԙ$v���Cs�T�^��gh��-��͟�R%�$��&	���i3�9�d��_l�:GH��6���Ȁw7���ݯ3���˷ĝ�����+p³�⫿&���S@Ѝ�H����M��$yЏ���v�1�����wM 0X��j��ʁk2�y�t�����D���	����h[�b?W�n�QNPZ�2�c���L�L]�R[8ͦW��Fd�4���6��^t"�xt��[ݘ���~��1�*���7C4�N�e����Vx�n��4{�ܩ���*�Q�(#�Θ� �t�߯k�z7��c:p�v|���u�e�ӛ3����˲^���
Q��AW�e�@~
"��	��Q�Y^����m�ER�Q�S�(������.������[�ыO=���7]H��吊�I�n��y��a6+��J�lٺ;�eZpCfS���X\NR2dg������P�B�Lh��㪫֚���R>}68�����#��~�t�U飘���.��0,VV�%�o��5�X��6ʂ�t���yd:w��s`����v�^r\�`��VQ�ƴJP��;�_`s�X���fyF����ׂ��6���C�Km��:�����۷���}�#����ǒ��G�YM����r^�<�I<&�oþn���4Y▏��r�|�����l~�\��"[Ĥ���.>0F��I�έ��p[�j=|Jl�l���g^��j�"�-+�Tm�Ŷ
�� ������TQr�e�����kH�+�-�[�����=A������H���g%s\q����8���[����\�v����Wx_��C0F���(���_U~QKQz�|S$&f���N����ܥY�5�ǻ����Ԍm���f#7���t�����K�����~�&�
^�]���ZY� /ɀ����
V�h��B:bguj��L�A�>���Ƀ&���_�ߍ�)U=�11���Z��%���)K`����I'g۹�w�]/���V2� ��
,�v3L|�d�G{U�S�p��8�����U9ܹ�9�Q)㌪��D�R�L��@b90�"ڹ�(�GV�y�_x�l�۹k�#(���8�㵃3��W�l�P���MS�^��7�<D����ijsz^o�L,��!����>�L�kh��S�x�0�2ROE���V��l���@�%�%��G~s%q�D����p���1�قD�t�V��(3�ɛ��_�<e����!7e�I�Sq�=�c��K����`)����d�g����҉��g8f+��Y�LqLK��%�))���U��� �"���[=?m���q������e��a씏ceמ��8V���T7�Y����#��?�3>NX�>��l���D�$qg�S���Ͱ�R`xܣ	�Ds����A���-�E�7j=�h,�����U׉*ї�C�]k�	���U88�gtz%ojZ��GY�U>\:2H,2�0�y:�+���H�`�������)Y����Ta��3af��	��%��������kau�<u7��K��R�`�,��94�8��xD�p�\6�-�۠��2�l����f��p���n�B��šE����e��Ĳ���&D�p��w�Ȫ&#A���t�p���p( :t�x�M���������¨�t�g1!H��f ��v4&�0��:pE����:Gi��[i��2��Kխ+T%o�6��ʒwm��t�~m~;*�ټy3�QY;���O��Ή%ڤDl-S�|BT#��c�SV=�&Ͻ��H D��������Q	�B{�+k�Kă����M�G��SP4�Y��+�U���Y�dj���hRR��� ����՝0}�����P�
m�����eP���DC~k�WPv�|��Hϓ��]G�/�@�%�ȯj��q��?�EO�,nv�j��K���㮈��#w-r�o����q=,�P����������Tf��eI�-
����;R��6�F�ƙ�޶�,�����\`�����	�s#��%F>��j���
�ඞdٻ�e�w�m������5q�{T!�" �X�����s�v�*tc��6b�m<{0���/����1X�y�_f|�7�Z���:�&S���*g$���_<rCe���n]PQV���VfT����'7ݫO�{mݭ^�g˪�y� CEіӣ�-�J�WU�)��� �ŎQ�Vw���c�q��c��F���#,̝Gs���F��#���tQ�P��GW1��"�`��9(�3Yq���2n���u	���]�� .zto8JΝ������O������=J������^ƒ�ÏW�7l�F�٫jT�H1U�[������Zu建��~T���V �݋H	�WbX�B�شa=^R�˙{βj�y�KE�]�pi�����{XC�S�V_T1n.���#~o�$հ؅D"��q��u�$)I�).NVM��fV�Ds���r%6��q�✧i|��Dkgn�Ov�%�r����zx������$�O�<<2��q7��`1������:剹C��J�LC�b�b2��]���:�1	��"���7���u����ɐ��Z�9���
=W➖dvK����0��x�Xrr�p�c����Sǲ�qYYH�7��p�
����5�n��3:m�Uh"�S�T��h��C�M3I7�9r��,�`�Z�UNEҹH�1�]��������K�_UPB5՚w��n||�Vڷ���e�?u�hXᆮE������P:�Ϗ�%���d۾%��
��,u4��$_W)0�O`�u}�G��p}��$��s��Q��T���x�X8�/Ç囖&��?�����׭�N�4Yb4�K�q	�N�"M(=&�����E���ݶ������WT�����E���؊��A�I����L	nB-�)�~����Fx���Z)0m���R�؊i��K�zc-�6�>�~f@�5zHՅ���Te��0�ٸr<���^��^Qq>
�N=��h�զ�ǉ�p)!��z�(@NI~��Q���Ru��t�Z۬l��}&:�P�a�7<d+�t� �Q�E��Z�A��SX�un[j��6B?�"�'"��s��:sw�������0�w��I)����������,�	�wD7U�||!\��I�'}%���g{0���}-(��MDH������������t��I�$�e�á A `_׭�,��=������UT䠑��͙m��+6r� #��*�0�t(�=|�.`���$�:< �>n�3*r]�.�?
˓���u=�@<�1�bd�ʿ���D�L:��6�́�*��d;�<h{�=��]~w?���]��l�w��34���X2���(���f��W{�@&CY-p���b�`A���*��_񚬟�_�>��g�VG�	ӓk-�i��c���eG�ꠙ�9�!��2���N�
yR�z����?'��>�̹_��po���נ��]]�㼭Ǎ��8�
�H�9��� �8 ?�uL��`�>�,��,VQyMt�a�����kx�i��ql������*����@��̄���a�x����݈����C �M����.$4��K#[,���|������U�(���2�}��r`�F��(Μ�n�3��y�\7Wo��5��mv-w�)!�Qk�R�5�G�ݚ�����@59�+�r�������=��C�LN߇C%xjʅ�8�)�?�M�Gǲ�G$���Q���:��,�*+�q�I��iC��[;?�z.�K�?\"������d��n{�o���m��q��8ŠW�0$��P�����Z�*|M-SW�����9�?D�/$��V>g�G��9���J��0/}���,�9��ϠS����b��Z�mH��}2��Cz�Y��?�G��U^p���e��3�[���=36<7��?���K���c0/�F�5-�V�$��ԙ�r�(7��;"��;�G��N�s�`�2<v�A�o�޶fWm����Ѿ>�#��qsj]�������ě��׏��[SL͹2)~�nEGg�7��s��
\��0)z�S�R;j!��A<Y��!��4�X���B";�n���](x�m<9�/<J�>J]�����.,"���&�Zm��/�%2���EG�K�W�$���9!�"4ز��
vѷ�Ȥ��|%$�����n��)藧�vM��<�#t�Q[.��V�]M��˳J��>5��O[0�~_�*��o���M�=�m���/��n���h���\�J:��~P��PԟtS��B=](�$.��+<~.�>>0��Ì���r
ڃg[�L��34�:��У��e����4|�]�!���~��Nxd�%���L�G-O�O
x�=Wgɥ�M��s���a?+ʈ���ĺv�&�!{A�=�,-�+煮B���	���Ŷݯ�_wc'+�o��R�~�fݒA�$���� �����/z���d�[ЃXh��0BL	m��H�hk��|��w�];23Cn�@�P��o"�:)�:!��,��`���V8<��P�'?;�y��<88�d_
�%��W�o��[M!.�qS�Ǣ0J�����to��4�	�2I8��<)kY���+B
�%6�3fk�w�WO.�_��p��߯�;c�_Xל�r����ʪ3������Z�çw�`超>";��6j�ʵ34�F�si"0��nAA�+���v���ʜh���\��>����Ϥ4����^�\�~K��y��``��p�������PƋ���btt����l�E��r�,嗝 ��i{/���R�ԃ��O
Mp�I��5�y޳'�#T)�"g�n�uv�5�)��a��C�?7�Ƌm�y̄�'�T`E ��H���w GlX��슩f[}�桦�4�dڷ"����&ߙ�E�C���DB�ښ�+A�_��V��AD�VR�� x���Q�Fs?����$��*:�
��z��s�Z{�E��Xu4���� <u�&W5�!�g�GӴdd~�nۇTlK����}ź�,�.gҙloyV�lr:��Y�Q�h�ά�ö�x�G7x{ ^V���9�����#'(�ތ����J*a��\��C�>)"����X}��h�b~:��������*�Ֆ�	pfh}�`��Ώ�ˠ�1X��v�A�n��*���N�a����>����[%睽��4�*Q�;��y����=�1��yDس
�$0񩛠��VEIzI$,���$���C�MIVv���G��Sw����&/���Fܕ��/��'��3�͗$k�Qȱ7���aO����s´��P��t_��K��fu���E5k��-�sKu��dX��t���)���f|_��V��$��ۣ˱�og�uՊÌ��V�{�k7G�va��E�w����篘!ѐo%�)��0�8������x���m\�%�)�b2]�{�%t���������{�������l��ߍ��6N������Ko���������\����v0���K�;��2�<���ߜf@-�2����u)�XT��{�*�}��k1���b���#��73<l��i�t�{B�Ɗ��B_�HJɀ����NE:vs�Cr>S��bYS�_1��2����Rƛ$w�2VL�2��G����>�к��.:�s1�����x9k���%�#�S�Y�� ���GG�s�dQ��ȣPT�:%�LYL{oɎI��U��1�yTZ�@�Atc3�G�-��9E�Zw����Kd�wkJ���UY��4F�O]sK�ר�ef���ο�-���-�%p�RY�얮��Mu��\�\lJ��p����P�bhFh����cK-d׌�6������+=�e*ߑ꿣��֚_�����v 4&�����|�5�{��'P�7���E�@@k��d����߳F�	/aӋ�Z�%�a�,�<��_rF���;��������
v:��.��f<l!#T�N�(�M�T�Z��f�q 
���e쳠�c��h8q��p;����"�����s��`�*R�'_�s���?JP�x���d������[\
@�$�����4E=�M- ��9������kU�]�M�V��
��v�@��Gu#^�b����]���|
��>}��af?���
��g��"^=֨:|4�kY[@]@ǭ����<ld��HPz�ό��zh�b����+�[;�?� M��gm�`񇸸)�S���DL]z��f�����x��x��U#��R����R�j?�2�3�8����h��4��Hn���<����^��Ͳ�P�p3�.�޴�X���3kA&��FdD����2�P3_T���R�E�<����/q��<��O�n|�%cwc�DQ)4�`�O��i'Q�ҦTX6���^\�3�;
&�B��47Gy�n��^3A�	��*��)��ݦ�o�x���&g���.��3���y��}^��R�33�0���aŔ��7�ݶ������r8�R5�jױD�6��X���je�W�y+�2��b(+l,��~/�!��!�&�)����oB`��[�g��Ȁv�M"U |�%����șX�$���~�}������6��lB�b{��Ŗ��Z~�0���}��ު��U��	Ct�w�z$ c��e'���*��B�n{R�z�R�]���I]-�"�j�7�S�#�BNt��H_`>�A6�8yR���8���t��;9X9h��+�|�q�/�4u�M��~��mf�ȣtF���k>�>�,�LeM���_���灶%/�� �����(O�
�tqS��5�R��$�>��n�c4<��N�����O���G�Ց��e�-�Ԣ7���E��������F��7hvu�o*L���(9ϖ�\F����{�e[Ϝ
�N�C�{{j�T���-)1_)�ٲ�j���n�߽[��G�@h���(���,�t�Z��������������ce��q��8�	�S�z�**k� @��Eg�"��-��/澝nRw:�-$zr$s3��ӓ���ύ�.Pz��Z��爫�R��o��l;�R@ݿ��:[
�d=�z *��`Rm02m��	Z%w�����T�paw��m�h}Gر>7����ۋ8�h�/N���J��"�g?ُW�x�_oQ�ݨ���@�o=����~V��l���6��QB�nZZ�ku���ab Z�^{�t_@�*��Cy�>ޏ�k��Y:�+g����M��f��,ox�h��c�?��	�O�����|B����II��q������OH�ꑲ�_����ǹY)�F��CD����aGt闅� ��*3c�������o�-�DA�>���.c-�$VD��Ry���
��[ټY.��Z�^�Ye������{�b��B*V6�*K-?:���C�먟sq�>���̺v�l�ev5��M��g��裃wT;�GH�(�5/���TV߀2~�A��J%/��Um�(!h����XY^
�n'ܦ8V�D�t�N��4V���e����O���_RF���G�_aj%g�	#�fs�V�pψ���_MV}�F�3��?Z.��g�4�?|5j�,Ș�Q���'�;*Ry�[1v������v;�}L�f�[3�B�K%�GSt�~X�K+1��6N��:#J�KT�������(sUF�3���F��� ��y�qO<}D#-bF�Υg$/�³K��9�v�#;Y�����?èF3�u�~'�r;ו;}N9��� P ����T9��{�*�yF�[�2�9��+Hw��k�V8�p��QXd�m�^sIv
�4�����_�|f橅!W�-�;1�@�X4����Ʒ�"���"��<�]"T��/�ßM�T�}�"*���:Tώ���.S#m� �zt��e,S���*��vX>wL��{�iכ�f"Gh��V�PCEGl����3#�Q��[��^��~T��c�6�x��i�֩z����PYy��D��3���A%�(J���?�V�˖% �a�}S롁;jX�M��;e0N#�L��`gKQ�@�����!#�W�:�і�Nl�[~�8�M��x���ϝ4	8�{�:]��rsڿW�v�R�.�,s- ��5�%�&
�ssZW�u�
w�_-f�� _J����'-̠��T���A�o@��'O���kS6E�%�ȗ�2�=6Ui�kW$:��% ����L�o
,A|^]��,������C2-�<�T�k��dV{Yd��Ɣ��u�go�&Ӓׇ�_���4��`��.�LJ���i~�*n�[�����t� @�Re���?��wݸ*��i�T-��ws"9�9]h?Y�L��-��C7�	/:��[�����sw:WO��u�vt����p��T�ѻ`��g0y�����b�Ƚ���ȩ�dU(�{vX��h�#���(z$��0ןe�9�Ӵ^�t�D�����}}�<�֚=(��/���I�����Ȇ*��	�&ٻ�F�:O�o��\��Yq��Mܨ��>0-��:�N�a�9t���%{9�U�0�W��O�bsV?YU��Y�j��HA�"��}檂�^��4�
q��QBF�m��&	�͕,�Q�.�#`�����J���2�O�̧~�-��ȁ��T=��5���W$�D�ب��A�`~7�8���5�\gd�X��%�����<(��=*a��y�P�
+�)c19�c��J�WN'	1	A�fj��[E���u�Qn�>w�;fS��n�$��Q�坧�'=��z��ք/`������%[~��}�:q)�r�D��Z��6�N�XR��tPw�G���3:�m��d.h.��g��
���2��!OR(cf�uw�*��\���c��1��d:)�Z�a� ���W<1_��9f�*(��q�J�<���/�/�W��$�$��yZ���ο1e'���Z��6;%�2#q:���:�n�ɂ\�`p	Cn7������,����ãl�JO�2��=���łF�m�{D�T?^Q=�*�Z���!Y����rD�w;0J�<��<G��pYaR#�{qq7�G�7��~�o�w6p��5mËb�q�1�0��a+�zI�Yv������LGE���P�{ySԳ~����j��Y���j�K�f���-��=��U�(Dt(�^ߞb������i0���uk���ڴƩC�v���H�Mᅗ'4}?�x�u9V�;W.ʟ���`��Ӈ����"�a���K���8��X��v!���Z�eۿ]b��^?�"�	 ��B�^�̅�Ҧ�ž뚈3uq�}Yj ��J �!�Ȏ�Eg f�.�w���<H߰2��	���P�h����YJ=qx]ӂ��m�ڂv�4��+ڪTIU	6`����&[�T���u�ؕt1n�ě{f����5�No����Fc������A�i�ݧ �'��j��^�9���9I�+ƝR}v�4Bb/%@�^�!���f�KK� ����Ft�c��"y������D�>}���Z"�����Fv�V���JO��F��������44����W�F=���	��-�X g�e�<�$E�o�7��y�m�<Ga5��!�vz���wL C1XM����n�Fc�o�KZxѣ[�y6k�-P31g��r�}d�ek��r�#�5X�i$)���EuTW��nMZ���$�}�L�{��W��DD~�PP���r�!7���/*����L���0�!���M7�%ѥ���O�.콢��a,��ѬǛ���b��%����N�kx�5y����1n2��Z�w�>��İ?�b�C�8���i��,Xٖ�=������O	�H�*q5U�z�萌�-!��\��or2d���t+5��s��\H�.&R���ӆ����,&���M����l���NK������t;G�w���V�C������Wv�"#{_C��ֆ�f�G��n��X�陔�l8�����]��8�0�axE�,/ǁ�V��X��n�6�Zʨ��8F��\ �nW��������Wę�Bn�2$�r^$�e����j,ؒP\q%u[�#�q���*<&-������W��VVf�Ul�#.�m���"k���yR�Ѓ�݁@P��Z����#�}J7%�a"'�O-���[�X�a"5����}�F֑��c����1g�o� Β���N�Kըl�]]%�'�"���A�H��sr\!�f4Q�u �	���;�K�18�ݖs�����V7qΧ>�K#�r� � ���0���ag��y�cʖ��[��Ul��\Q�iP{��L�#x�xMv�= �e�F̘�R���O������ve#��mJ�.p3GMR�q�<4d�(��C�͂�<�Z������ t��<z�����������~��O�r����?����i�C�m'���j0}��A0��d�Ǚ8>��A$�Zͱ�@屰��4��n-F>�ޖ��%�(��2K �O����8�w\�MZ{��T�8��D�(�1�������6}$ ���=S�������Ji�+���8Լ)"LWv��U��l�"%��Sf,e�{me>�3�h�����M9Q�X�ȭ4�G�?�5l{���������S��_c��ԇ��H��|
zBl�Rc�x�q�Y���P��mE���1՜��*�4>;���4���iM|�MCIlz��D!Rz4��Fh/�/�����f�mʭ�/x�!�ȏ�w��zCt������E��]�̫��˞7��n?�A������V`Q����9Y���0�T���6H�}��K�=��8�6�����J��L�m��|z9�9Cj���{V�͓W��������\�z�X�tt�.�z_����
�R���k^̰�X��3$K^6�X�C���*ο�t��ʿ�*�:3��35_=p�Q�L H�ŗ�X�ҷE�ח����7&g�A"��A�-IΪ3�eB(��'�-����+�\0����� s��"���Z�ͣ�N7���s�Ǌ5]��(<�{��_���{欁��P0�O������J��^G6Ǚ?�ƥ��T���K����o�������I���W.�"!��P	b�2��zr�-I�f���8_�s�d��K���a�"�`�G�vM��͔�J� ��r:6M��*����̪�S9zuf�7;0�W�B�񹏭�žvD�ؒԄ�%ߛh��A(�R��=�-t�3[¥[1ڸ�����vb;ʌ|]:9-��K�n���"�1��[��� ?ѺDQ��h���\7%�����DČ*{��>�x6�3;��*�!6Bu�[ufZ�d�w��߮��7�m5��T��m����T������pܨ�5O��?K!�B�y�b 葽����x���4��@�V(����.LoK8Yl�p�Ö>	ƿ^/d�n�e�z�lD��b��=9��"���u ��74�Oa(F~}�66����nL��9D�� Y�4��g�}h$�����@��-+�e�x�P.���!��^��^�x��������=�A�U��{yX��ja5Y�w"�f+[�E�bu�}:�b��V��/%VY��\����^΂�;giq���ҕ\hΑͦPv����g������GG��?3čH��r�*��MS�٫����@�5��_n)RF?5H�t���t@$��5l��v���o�`'���]�yJ�C�19[�/-�;^�M�x`�C�l2Lwf�R+��eA$�͛�`Z�g��/|@}�����C���a���f�"�y3
�Tna�g�y�����؊���'��:6vվth�y����wH��ۗp�����dj^�m�XJ��BB�rF�:m�S���#�F{0}���q���<�a �/Gϐ�&��dA<�xA�����&�8�D�t�+���5�����ՙ�B�ON��'@s���v�O~��g�xEx�����]��w_�P{Gϑ9#W�i��w��؏�I}ø�I�%q&9��FL��𰝲��E�n�/�g�аPU\>n���6����[���W9��&��#6�����7����r�;�����e۬�}�@���\H��+�k�puW��4�!����i��ߗ���R+)Qf\<����,��Pa|�����@{՟c��k�t�oۈ��v���4b���G�ɣ�:S�L����V�����
���+���r^m*��&7r�zCc�	s?C[[0�a9��$��P��vE�l�6��]���k܄M�j7Ý���e��iKͺ�?R�B��̒�����j^�`�a�Q!���t`�����e��[����l�9�|�����KO����D|�r�><Oe*�j�4ry��B�h���������wm������m�Gͼ1a-���E-ñ0�������]ˎȴ�(�>Z��Z�5��]m�u���}��]��qh��|�k�?&]��g����(��孓��p�C�Mn�.�?���TYWq��&�r��g�
I[�r]~�G���ɽǷ��=u
�!F�0k5äL��#��<��*.Gq�"�2�1l��V�O �<sZs�*a��0����'�(+��Z��/�#6����7~Te��Y�#�N��S%�^ra���Q�N�i�nBL; �j��U~�)��ث�n2Ҵ�e�]����I�=��$2�|M�W�90n��xD�p�C�J4�L����"%h/���"�?p�u1�{����J�;��(���<e��ϒ�b�m(���S�7�XЪm�^��ur`<(���(T~T�֘vDp�I7��.A�hx�˖�p��X��ۢ�,�T3�Կ�������3����v�9��8��^�y��t��%r��/!���t�{]<;h�]j�Q�jo ��t�R�z�4��xlh�1_��36����ԗ�>���8��ATv=c�
呿P?ۊ�&���Z|M�S�9:KcY�o��|�!�ĿRņz��+s���d����Z���g�?M��7�@���b9���]��$�䑌�)���x�{��%>�$j[�f�Ϝt�7���X+W�O�m3�x"Q���9u�p�|�$<�������-a�'���D��~r��on�4.tʫi���JOBZ����-]�N�� �&D��^�9`)[�� HB�~����%7��n��V!*U@�������l�"yz�~?��*���}mE�
�̺a��8��f[ha�q�6�$Oi�d��A&��`�w,�v����.^�d���w�Л�o��"�n�dҼ�nf6�K�#R�pS�����r����S*�"�@�Հ�4�3���� `�7��$$���)@�|hl��J�:��uGa;����-���z6�n���{���;��	�g�*�'�c�b���	T��Z�S&�:�?d%Tlj�'�'�?�	���.n?��e7��H��HWLĳ%��6#��#�-i��#dʆ��|����Ky3���q�(!�,wb���["ۋn��ٗN=f8A�G��Ǉ����<��յ��?��;mf/�,ī��f�yD;J.NV�3P�Up���)�Z+	h��kE�x�K%-DЗ��.��ڥ|b�����Bc�4�Ҏ��:uiY=����n�\��tZ$�ʽ�4s<��k"8;r�&ة�k1��gX�KD�{�d�#�@b�hG싴�GiE3�C��b<�e��{��vbŃ3 ����6v�eU!�w��T��,�Q�J��_Dɋg�QJ�A�i%��n��Y����C�G�Ԏ 'Zb�7��_���Zl׍
�Gɦ`��oa("������v9�6?˔!���é�$#w�39!�#kǾݪ:a�)�B���{����(,�u�L�[aQ2�����+�҉=��|,�K�-r��@�򡼢�T�J��Ik��z�����խ�O�K���L���	��#F[J�yP!_u)�s���t��d북X����B�n_��%�����QG_㾺s�d�����x��^46�k�+o=��N������>^�,�5��.�s�wk�>��;Ъm����ܮo�w����a�m���܆���t��S�Կ�l4j��D�� �3��Z\Bw�q/� �q�j|
�J"KV��_�$��H)ND�sXkrc�r},��e$#�I���d�|����t��_�H���6F�~�ʆG���:��Ag̯J4��w{�갂R@X;��x�3k��Do�0�a�$rrwf���TG�$���pU�F:H�#.9�P�!c�o��C55�ź�A�=
yj�2R���	�á�lȒ�,
	��
���.�=N��&�a<r8�ƾ�-�D.E{�S��#���"gL����3{%���7���sYY~���U�ׁ�1q�!����־�H� �*�8��׼�3�@��f������1��N�Ző��a�J�s&����Aj?��nr��v;���dpV�������������?�2�i=d�/W�M��H����04ѓu�B։#_��9m��;Hl�6��=��;WΥ�6����CQ��Ork��ŵ�8>hk]\��t�� �"|�3������k��HL=��`,߫����@�=�&�!�*�������ԤA:s��@?<p�ZZ��b���V�Ps���8��k0�WY4���DqXca�Z)#�8e/}��~X�P,.�%ޤ5�:�Zdy?���iY Q<�#i��� �Hb��5_(�F.��Y��pJL�Q蕴�F%׋��۝��r){�NK[Y]B�g>���n[�:#���#���i��U�bOP?����6�0�ylQ:'��_���u��<�پ�IP������D� j��y#����A2#�!/+k+���v�}�^������F�H�ݥ���Y�Y����`q� ��h�a�R�G��ym��m�F;����ae����׬5Z��4֘Av=�i��j`p�ϰ�v�������>����r�¿�h��b���'e0�F��Ӟ�	�F{����![KD^���&��"T�)FD#8{�� ��]�Z΅���A1RU(�l+*�"O��/��C�p�-���I;���y�bwm��<!!���P�qX3�;�Z�+rOP�Fk�M��R$51�4��KSB;(k!���u���jzȲ#�hS�'�/�Lr�m����o��D���m:�PT�~� �{��d���'�*��b,�-��X׀d7������FMׁ�5��Q��:��IY��ނ�5	���} �LK�{���;�%�U3��RWd�}׿���{spO�K�����;�	�o�]��q�7{1���1��w�fSvI�^Ľw��Sn�_���i��3d��5e���âs�i��Ak�|�{H��'�p]3>�����B�6��p�zz��L��+d�S��V���`@�[�v�8��0��3�5�h�t#ǏN���0�c#=��#�*>׈�C`}�ѓ�2a��A��j���2{me1�ߺ��o�F�!�i�=<���D�:�q�bh�t|,���2-u�Ř�1����DH�k��"���<�G���*�H	�T.� �9�ٍC��A��{������Y���=(�Z�d:���>^gz�s��[i�܎����i(PD}l�:}�wX�d��DcoXsچ٤=��`�L���JD�A+��w"�gA��wR��l���V*�X�y�h�D;�L�*�0��)L�P�� ����������j��7��/��/�g�y&F;6�ܮt���P&�]~���|��X𖦙7�m�����|x�: ~��>�����U
����a��=�U�e��@2�|�
{������������޷�n�{a�Clo����l؇�ch�u�d�4�F�UcP1�\|� o������eh�!&���q�����B��en�`XC�m�uy�{�+�n��FT�Β�����q�S���8!@�v�2*�;�*X�$6F�zlL��(�u����*��樓#�b*�1JoB���V��1���3�Y�o#'1���Z,l���y��-r�U���:YÙsj�0U"�0k��;�ZD�*p�F��	�>J�UƯ��.eX�#�7��� 4�?�4O:rd:�H�7/P�9�F�)9���L�z���p�HW:}����E�Xt��N�9��kF�B��`�?V9��Q�,��&N�'��4����^�LC�v�*Ñ��_��/�O�3�O���q�Ȳ"@U	�tr�`�^�C����V��_1�U5GԩۗF�k��KvԽ��+U��s
-��v'@ bv�zM�GK@#�g�ڿ}�n��m]����7�Ҿ��,��}��5����6���Y22�
�[x�.�rU��L��}�H���?��_x?����dz���r�Y�=88N����u�������8�<m-i�jGP��G��4��D
�z��:R�(�.��zwѭ�歬X]^ A���K�S~���l���Ɏq D2#��Rr��6����u�{��a��68�6-�lo�]zPy�<Z����_���[�PP��.�~U����5���8[�f�H����oP/����T��1���H�`���Ƣ�L�	��$�\A}�Z�u�ǏF �C]x�L�yl�A>1bc��,:濓�����s��#�/R�.n{I!+#�@�^�M��6\K6�d��	/~e��*#q	=K���<y.M;K�Y��M�BpS3���p�BW����u�k�jinɮF1�e!�4��0[���bZv��Ĉ`�����hL5|*������ג���5��æIr�ݝ0�YI�gC]e6��ǉVZ}a=В.��BC��ȝ�l'�sP�K?hI������㭿Śb|rݭ�(r�O�v���|����a���}�V9��&���R�����"B���.?��]#5��ܽ�h�2��m#�p��W�飇L��Ž��_�������H@>Rm5��p�T���g+Zm�0����g=�=>��O���F�W�S���>F�F��
�����)֎e��z�)�xT��xy����Y�����Bʦ�����{���j)e�G��0�D��8{C��uf�����	�:k=q��*�D) �V"B�}�W�e����Eh\u:�:�|��(�H�.ryj���<�%\L�M���ӆ����Wn��M^���60r��M�Q:��Rѵ@�f$Ԓ
Y\�F�O}Li���2Dc������Bx~�SO<���s�k<�H������`44iGZհV9G�+y�4ٗ���5�^ƿ�s��X��$��'[9�k_}�=⇰<z����Ƒ#��̊J8a��P8f���Վ��my��|��S���,ci�4� �5�0�$�4����һL*m������A�ך{6��%�{�^�:�"�e������1�O��'�`%��0��;Ic���({k8ݴ���2K�g]�{M�,�M�6��*��s��w�kw+��R����mZ�A'��vr�1x@8-����Fv!:?|�h(T_�(&H#n'�1_]�w��Y��~P������&^�<GŰ����L_�����ݜ~=���k��Ȼ٫^��>��_#�����k�p�&�u�� ��� D*d�,��6�P�E�� �t�p��=�	�D�}1�ƙ�*I/�#��J(S�q��[�S2����IjQ1��9=���mfjU����ZH�G������%��V^ј�Ly�>�ܝ>	ѫO~��6NQ�c..�&j�9�����h��S32~�c���H�Qˆ��_T8�R����t�D��Q`l�\%��Ijɀ�6z�'?���ٓȏ�
�s�F�a��1�D+��`��.����$�iIl";B
=�cjl"�2=��G�$.�1"�'��={�p&�p�&���SO�5���B����5\���9��0�>d�Au�x.:\�U׏<�i����~�\?��zm5��]2.�f�'�]f?l2P��^�9�T����%���&7us^OQ�מ��%�{�n�жc�s�9�l�}��O�"�U-����p=��W�\50~[聳���7߾@�E	��ވS������aM�]3�
B[c�n�\��,����u��F�t��9:;6\�x�������BT���u�|�,)	ۦx�\����+d�4Kj9W�|�5t�9s�ph�%&z�no�� ��hF4B��W��j��(�ZON�3�7?:F�w��&cYޕ��]-�?�;�!Z��c֝�|�m�S�����-&I��g�A2�s}h��z����c���_�+�kv3���4�b�<(˄��r@�I9��#�W��-7���n��(,<s��6�x�v8rκ�#��Ní�57..��������aS�]Zc���4�t���^?G J�P�Bv]1��m.�Ѿ��P;�)�i�=�0�����މ�U�k��F#����A'���r�:KN$!7�]c�6��7��e����t-ZT�K�Z_���f'�Y�J��"]�`��rՀU�gʩ���6M�S��74*0_��D�T+���L(j�Ө��ʯiޣQEEL
C/l�F2��Q�@N�����g�>�R�r�	�k�MY0Pg���ց��y�|:�j�xs����9�dz��<��Us:2��� l����cL.�XGV�(Z&B|��~׮^O7��m�nȊV�7=����8��#���#�-]7�̲���my%,���p�����х%��2�Z�l�E����?#9=`�;"b#4�q[d�̓�%e�``�ճܷ����VX[cT�X(\I�N's-�{�$ʶ�@l�>E�����H�� KBS<Vd��'):��x�.[bۮ>��s���,@�����l�a�=#�pr6@��6��[+i�4�H��"tP�`뫊�\o#�L2j&X��v�R��5c������3��c����y�&�q��ƽ��������'���#fI�M$����ν[u1?`�U#g�Qi38�H�\ϠqV8�)�R/%\�a�_�t3֓���˷9��1(��fv�s�Mf��������4OՍ�|�+Y}h���a��>��H��q��ǆF��̵�@ i���Ƨ�� ]0�p?ѷ'@��3���w�d�$o��w���㘂h�"PQg�6��is���7��'�V�"�o_Xڏ;��=
��2%Cϰ����9z��6望�l���}�x� I�����M�0�5`,:�0����G�h("� �#R��W;���ª89�5��k���F�t�y���k�����v2�%i���c�#�E�Ion���o��F_*N�pސ�$6��GEi4�Pe�I�஀�U̹~���
�"|�"ցPA���F�eT��&��Nh�󭩰����<U1I���k����+G>l��1"�!�Ah��3T������#Ҝo�F)���5�׌|�xί���]��Y��L�)���1��?�vԻ�����?Fi�@��k�E�.dv�5���B`���n\� �� J�Z�ar�ݣ�D>���A��e��J?8w5����'�M����%IED�iinàg87�F�s�Yx!� ����e��\��f��Fᐽb�v��Qb��|t
�5P��o�萩��̅�;g��<d)��K��\
4�6��������t��a��{��`�9;�1�_�9j�
$`gTg��yYOSd'��pڤ<��d�S'���s�ɧ�I���/�skw��6B^z����uѵ�[il����Z�a۲"�&N\�~U2�p�2IN�F%7��D/e��a�2����Z|G��k��N�ߓ��� /�G��mz]ܽ�T�wpO)�l�s�S�%��6�.Q�#'�e�o�KYQ
֞OC�{R�<l��
@D�0��2������6tZ$�"����X!�ա�dTGG���G���i��0���ΜI_��g贇C��{湧�c�!�nl����? 	��1��L���p2n��%���7=�м?ԣ;9 	����pDM��F�a����5 v��أ�8H=�	GF����.�=x(#tTQ��F�H���Z�8Vmh>��`�s���E#�*aia�!��m�cg�^�i2?=^�aD���i6�qX���րE#:�Qz��� $��G':����˷�׿�z�ޤ��{�<���TV�(6��i�5��yT���}ˌ��f�gE�6�KXӃ7�}؃��R�/�g�pŶ��������S+�9�p-sӀ!
� �"���=�=f'��hH�C����rc�B��$��pf)����Y����`�O�v5��������)G�$�xd�IH������:μZ� C�C�}x�Q�mH]o��vz�̉�Eg���;���}i������IJK��s�E��������t����9������wQd��%?),��{�ҙ����}!�RZ4r"�`�d8|jլ��î�ʩQ���e���>ؾ�T3Q.fT�� �`��9s�V?D�,��yP!�pv������]cɚΕ�fT����0����͙R���&g���wlߥ��%�c��^����l�Me��t���6����:���0L�������%�y����AŪ4S�Ϣh�N���W��J ]GN�f��.�������q!�m�[6E;pH��pga��	� �v{��!j�m�*Q�J�����l�:�$����G��%�e�D@B�6V�*��u(���rt��2��P�9�E�s{�����
l���B��׸�<�ΐ2tB��``����Th�OV7��5�#Z祃{'�E�%ŷ��$�h�5�N^��#@��.I����I�q6"�E[lo�z��	�n�Y��H���/s.�t��&i�������~k{�{�EE�,�vg�3�z�å��*bwY�et�@S<��R���hx��
D=�s;L`-�LqP���ٗI'4�U����#�|���Ci��*5��욮ctZ�RpS�u;m���X�h��U<MH`Dæ�lbЈno,K�4�(�!��/>h�牑\[��l���H���'{�����l�2#VPEW(^7�[0ZϾ�*;�"@�
U70�ۢ�ݑ�1fP�i.�����L���eC��)7ZW��x�x��Ml�4���AT�Yo�c��u�}����䕛�E1B�јf4�?�)sL�2}-j��Q�C�}�`�s�;m
8_�����y��ak�K�D�1��r��T�M��.��C������ʤ�8������ہ��A�~�"��q������V:s�%yi��*s�F	U������q��x����=�n���Di;�y�iQ����Y/��y���ʓ���yN+{�̸���P.�G^_�#Í9L�'#����
G�(H�pX��A3-"T��T�F�F£\�Q��>7c INb��#^�gee-MO��L#d����il���Ji4Wxn#*E</��䕄����N�"Z9�"2t+��e�+�>	�Z�yf�&r��@��>��1�lNC
�B��M{HhD%��{I,��3������53���#�5ʸ���r�c�k8_:%�u�6��!�@2?�y<on٦6:��̇���^J4���-׳�sdu���<���e<�la\�H� _�������d�P�O��z4'�����;�j��N��UJՆ���?q4��
�pi5-ݽ͑� �1&z����W�ɞ������}��q�4)T-�[Tc4p����%ZP70���A�:�����{���X�K�ܑ�tˤ���;w6��!m�:S!AD%���#�"vA��"�9�oCi�����D��cGA`���ϴ��VN�O�qe�V;-�Ay<��;���8Ԓ@�C�i�g�׈�T�[�6q���z�F�a����z�dsI*
C]�$��0�f�.�<r���D�ce:�l����w��c��<T�3~W�ij�kier_3��Dd�D���O��	ej��0G5�\#/�0��f� Gu)���X����>4Cx��G�G���ɹIy��������&��0���ڄ��������yY�6��X�j�������\�K?��/FY�5�+��	
������NT#���F����vUY�޹��Ǵ4��8�-�=_Fb�#�	KQj��zp��$*=p`�k�E$�a�����x��m�����-�A�`�<�񭓗4��S5�I� �C���{�^��4]_�����0��6� �MD��D����fD}�s��8�l��ߡ�����?�Cc�uW^C����n��K\ĉ�r�3�'��Ux2�%��o�D�Bڹ�N9sxaKxx<J�p�h�90 Q�OI<rtf�E�D�qޞ]N'���P<>"׼nco��j�e�t6�9P)�8O��*:���lT]hy-�NB(������ ��:�tU�]_>8#��k�nqw�����ge�9��N�;;��D�pҴ�:���EŇ�9�3�v��QG8xVa�Z�j��HS�����a��5H�-.SB@YC���1 X܇�?�!��Gȣc�<'�85�7D��Z׌��P��n�Lgy6���i��ڕk�2�,�ir�����{w���r�����NZ��[Q�"���땕�?�����!@���5 0-x�*�@P��	Q�:|��_�Vk�d˼s�v����0���.�\l�����T�p ��W�;�1��N*"�R� ������cf��O0��Dԡ/��v�11>Q��f�>���Ҡo՚S+k�}���Pe>[�:����E���W���<��M����E�� �R��2����4F�]B�F1�eآ���:�'?V-0A~�K��~�r��cQ��F��<+c�h�,��xz(����z���� �1���gLc
>�٬ȣ>5�3+>7��4l#��"3� Äa)gkWRV��dd��ђ@���� ff� u�B�6�`�E !�����x.5R
UO�/޻�n_}7��W��g?����O��v2}��oQ|/��Fq���k6��!ˍTl�5d��d�l�ns4���j��Lc��U��:�_�>s�ʟ����R7M��!5�;g?�z�sw�<���n/���z���cG�D���������g��:a�:c����,�����w_���qޜ�L9�{�������uS;Z���-�q��N���"<��:>�^��aP��!����2��!}�L`���#ߊ�&�1�w�k���Cc#�},�X8;""���!N���iແkmX4�5�u�N4a�����=�\�=£�I��W��/�V>�(�㒕���l�,�,�ܴ�W-���o�H'FGP�y/��y�Z8g}�U�@T��۔DYjjgƣsm��{���p���M�����1M5��&4�u"v�!�YG�ΐ竓�S��HX��rÒ@�n�U�"�q�B�K���T�7�*�p8�y�%��xpY�W���V"�π��A�h1K$z��7"E׽;Iڃ��g|��M�f���z�x����B�{�W13����uοwO�|���Z���YF^c���ZD����ʜ�t ��ܗ�oB��@�8��6��x��� ߵ�49s�F��&0�>� ��r��t�pO���/�1F�6^��V�S!�`� ���U���^�E`�3��u��UR7nܦ��IFE?���ƑK�鋿NE@�n���
�O�г
��l�Z{7��h}��*��"�1B���������i�=3l�P�h�����٫G��F*c��OE_'B�y-G��{*+RD�����°�$�ap�F�J�]�s��"����%�P�C�Y��J����w�8 cK|��kƤB�4'����PUŧ�'ndc�Bͬ�l"��W�2����0��0鉟�%�P��:��Ɂ]��9/C8<�(5�<�͐��e`���t�&Ց���XJ����ip����o��^yxv-�D8�L2�k�A.P��KG�Q�\��	���;�>��Td���(Q�:��.��&G�1���0w+�L�D�t��Vׁǝ e����t:u�4Uw�ŋ�D/���n��(��W^K�o�u ���<�z�p�vD��.�I�y���������7��T�g��M�WDvP4X"&���4_4!	�g�@\M�խ���H���d_���?|gT�ʡʁ��L{�o�GtS7�E�G$d�^",���<'�N4�tE8�2�Y���nd�=�jF�:WU���%o
F�����-�6��u'T��� �q(�W� ���ذ)�JB����r�lJ�CPӱ��� ���?Fh�h8�.?��;0���Hf%C�c��(��-�c���6���~��q����Q��q��NE�\�X-+S���`��gu��vj4R�����?tD3���U�岭�Q������<��h���e�w�r��b^`�3p6Xۛ��
i�N�΅k�j��2={�b:}��p��JY��	j�-_�;P-�2�7���|$��?�qy^O�@jE6�=�x�̧?Ǆ��N�$[M*,�\á�"�_�߅顙=S�8�߽A�d� EG<�.��K�M���w�T��e�$7�\�y�	�E�e,�;|"��`lh'w-� >����3K���s;P7�p	�w�r���4;a���֜Ħ"���e�v�W��2�7�'з90�ۀ�H	�0�6PZ?���2�yh����'G�t�q�T�OdN��\��pј���HD�gE/f���B�Fj�9�f��Y�u6�D�*���|��<|�s�|_ޚ�<y'B̥j�F��[j4Qh�~�ƌ���W���ε���+��x�6��dss^������W""������|�F����r�<ec��2�r�&hD��Sa�rͮe;Aze�rǝq�ч�{���pŉUF� N-��Dd�c$Ja�5)��'	%6ҕˌ�\%R��O���0lٽL�z񥏧��f�r�N��ݻw��!�Q�}����/>��Iw��vo>r��D������P��W�i�L}��U��G>Ɍ@�h��Y���k�5�ޚ=�(it�'�(nC�l^��������:f#���u Q��%�L����Rh����C�� ;C�ֹ�0���!�n�Q�hp��k[�1����f���qz18��P2_�H�Lsl��$�q�T��t;$Q잰�i��z���16��Q������2()" ���;_�-�����PQ����r��ƻ�f �vߣ)�XP� �)A�/�>�P殐޾�e��s�9F�ꑺ?�kK�jh�U)6ar"��tg�w��*�>��-P	D��Y.�7!����~L��xw����2�)�En
dD�E����M��5�����G�NS�D�����2��!�/�#�lTQ���$|��ie�&�C�_z����c�bބ��0�i6��̮���jS�۱o��UP��n83��4G4�����"���.����	��ҊAU4�a�K�K9�1;<x �qW��'~p������t6H��疧�A��F�
�v	(n�~�>C4��{�h�5�3���O>1�6�0����,6F�v_�m[N3<��]Bl9�Ȇ��w�;Ct�ikhT��1�Y]�hv»Dȯ6���!�����3th��䓶����.CP�[ιE�|��ʨ�e�@����M�#�H��U��aM�e� KY0��[�<`�Z�k>U6N(#�6
6��,�l&��u�G��er����b��_��g��?����_���v��Ѳ���D��Y2�-RX�����r%�\t�:�HL$��m������0�x���k_��2��K/�B6"���]��KW�����/�,$N���|��?������s��HkcT2�+�o�1�h�A�U�ٹ�l��v������Y��A85�U�#Fá�v	#��B8�9��ע�ݵ�@���|�6(�=��a�c($He�^6�ʓ&�
Ľ����W�N�9K*�eR�9z��viM8����,�N�Y��EW8/��т�˳���]�@�۷ɑ����4�\����M�x��-�'��낌���ӏ��4��9�Eo,L�W�}���D��0����
Χ��\���J[�F�{�y8﹄Ní�|uh�f��}),���;�k�qɎR�ו��8�D�[�������cф�M��ӿ	�2���=�0�PD�T+Ɂ�}�7_	o:��ϟ��� ��L�{���Y��3S{�ۙ1��\��Y�
�4�2�=q�i&��K�CJ���GON���Tk�ԏyu���S��[3���f]mw��9����ѧa�ċ ��VV�MiT8��h���􄜪}9tu5��:Ģ3�����Ԓygg�P$�2������t6H��F}ܤ����k�Gwc�O��"0�d-Y�[��O��"��2�@���4�-�9��ذ˛,��y�Uf(3pbַzYO}��J��d��s�ػ*�0�����z#`{LK�臬e����ݦiR� 筍kb؃\����aȵz��:^쇵�ٻ�=����\ë����T������$�қ��ɺ$�lB�L��y=D,�E��=`�
0�P�o���0�:Zk����~����_�b:ql4�i�n��6�Vl���ϳ�m�mY~�W�"�4���#�U6(O�h�X�@�2�����"7Qȶ������'oÌ�9��$=�[o��Ļ�8Y����4��޻7�/����p���V?��v��|ϳj��1�v�4-�9j���r<�%^][��	�<���]p'Jk�P��)�#1��\7�C8�]n�5�|�����G�0�!F.3P��_��)�����X��Ըw9��K���Ɏ�.��9=�����,k�伾�\�C�y���k�F�J�^g�]�Z��c��@%�zzV��0�T�M�<~&��C��!)����ŉ�tn�������[�[B'/F�nai%���u1��ʍ]�<�;ߑGzg��(kW4��k�+k�����~uv�����{��Rr|v�:�=����9����=)�#"j��g]��Ą�]rZ��C������M�F���ˑ> =Y]�?��~p��$A��I.d�p?G�K��ɱ�z�E��p�o��m󩋗.��t��>�&��:��>.18
��ʭ�����tk�;-m���q6��p^�^��?���U�r��??<'��QD�'�5,s�DuFAW6�(X�9<�C6ػR��MY�\�Cg�iY�����V��>�2{�19�i�R<ٻ4sp|��Z�M;+���G��'���7G	T���E��h�ej�/ߴ�f.l75��ҏ��;����t�Qgݔil.Ru�3ી��?TJ�f-��ّ�|�e�ֵIx�φBD����������+?÷*x�K�O��^{���`n��L4}�r��=��a�|cg�L+�s���7�{�aU<X;"u�1A��P�en�&�_�q�@�{_�e��o�GϜrZ�'��2���߇���:���,cN�H|η;�L�u����2����y�
&��'��[�&r]���	�kR�E��#i�p�V�D,{g�#ojd48t,���7碳�5�ѶW�h!fF�|�sDj簬нg:.&#>�,F��	�"��4���I�2J�\mt2��I�C5�6��Z�Q����dα�h&�M��X����S�\�����f+=\>ټ���;����g�_�ŝ�ee���z^wQ{�gu�N;)�g{�K�����r���H?���x�Qq���3!-��Ȋ������T�A�y��q���i���k��GO�����#�P��IH�7��&2#]NH����85�i��`�����D?6�/�k=������?ŋ���={\��ľuUgc��OŦ�t��D�r����&E�6���k�:!��9,":\:���&�lQ�z�>]���>���?����>�� :fvpB\=�;����56['U�5�ҝF�f�����Ϝ�����{w���M'{~s{�4�z`mb�X��D��ٻ�!�{�2W"�o%�m���z&��6��,�>��,;��fC.k�\n��? 	��M�]Cc�#w�]1��'�79����������`s���收1��)���̍��&��f���X��FGzcl�~���=�}�B�R+��w����!�$�{�!�����t�1Wg��a,z�3��?S��:q#+!<��8K�s�����@�R���3R#�؊�� M�+c"[+�l`E[�V=�5���T��F���� �&hD���I�K���u�6�PQyn:FA�˻�B�C�D�1#���LqdO&�hu���O2����+�捛(��8vXm~�FL��1-�<f����{+�:��lUBz?��P�Y��q���覂�=y.�1��ү��6��L(���2�d�0#}��ߌ�Q]��1����_IS�i,���|,o��۟��s�xuh~2�(ݩ$���	_n0cz�p�ZW�t�f6:}���;0���if��P�w�IT��ghN�Y<__�aCVL��c��F3��߸�c$(���^���]�| �Q�����i��K6�����T�����։��= 2�eS���$�t1�0�E8r<�� v'��p��3��!��XG:9�>��Z���Cц�3"c��
���s���ۘ*�x�l�+bd�����L��ؓ|I�t�'�<qB��8�N������s�n���X#�+GS������3b^�Us0��é��J����t͹��ۙ�^��G~>����G+�TF].J��8��V��bg�J����{|��{-�"q�}��{�ôpLf�Fҧ^�T:|`"���I���-�ۋT�D���)e:4���f��H,�~U��Y��"2 y�<�O����Z���]�[Qgz���Nz�:��X�5�������&��p�\{q�Y_��e��,���C�)�����]�����}��m�q�R�5q�>�1�y`]���hM,o��i�v�KP"�JH:����#4r޿o<���!".�쥜i��;W�����~�r��O�gm��K��`�6$	�[ϋ�Р�r�c���<
CtL65�Ad�hc���J!+QרFШk�����5����6`��CDm��ҏ�"��M�Yn�P�PC�j�m��o��A��QJt�&)G"G�hU��%b�,�p��Y�Dğ�ѱ:�����[EL��}�t6�+�92��\�ӷziqy�s�)��
Ghv>xv�3�ȵ�e�����ێq��,�'Tm�lx>��%t��[����9t ���+�����y��O~���ԯ|>�ݻ����{"Ǎ�F�o
����ƫ߂���p����ә��/�QX�'��?�X���t&à_�|9=��Ir��!�����7^M��(������I��W��P	�*Z��o{)1��M\Ѹu���b:4��f�|&Y�)��l��U��@YG����s`6;}<�#B�p��53�Ϟ�wa�ߠ��GN�C��e^m�J��wa緅o-A�p�1��L)��}?d5�*ျ��`ɔ��=���k�uj�,�&�R�:��b D�goL*���d_E~�g��7%�ѫpD�;��09*��!C���mfv�D
��N�4���al~�@��\q����{wn�A0��:m�E�Z� �9��TX���No�:T@��}��p_�#|Z�7�m��de��LTg�GԠC�!�Z�2�zP�&�f'��s���m�'0�q�8���}���Z�m�H�X�y��^��1�N���m?;�9��?ݳ�P�L(з�(�Xq-y�w����0��Ыݴ)��� �)'����U��|�)cOW����8��2cA��䧲��ԘV�!��I�vA^�^�� �{���OA�%X�4)�?0�Ϟ�Cg��k�=[��Y��*OGz�D�s��0�2�F��L?G��3��o~��Z+Ѡarr8��C��8�@�[q	4�&��Y���J�c��ˀ������$W�ln��jt� �$�h�%2i��r><r�U4jS����bw��&6� u�B��WG1Iޱ)���<�>�m
�r�6��k�kr ˊظ���&�`����&kH��*oXfm�� @��2+����Y��C�xB|�-�3���mn>kZI*��S����];9�0X� ���rL:c�D�#�[y��U<:�q^9Z��q����ϾU���Vz3�:�����0n/<�4p$9��A�/�6���4�$�ur�+���(�S�O��|�s�}HE�%���Nљ����~?Z���N{��SG�q�'�Z�;W���K���0�l��&��ߌ)V���8���o���H\����܁JI�P�x��L:s� }��F�߫�&]���a�v�k�_aJ��Y�_��K�yr�v���u{?MEΤ�Qg�w�{@��K���l�B"d
�k��/��Ȥ6��8ՃY^9v�f�/��lKk�0O��X���<R�=*�����Ǡ�3O��9R뼯S��Z��{���=��$��lr�<Q�E��;�p��M�����c���2���7�E���4���>,�ÈY{�kū^.yz��B��l���^z�����
.3q6�KQ�k�ܸ�O��T�ߓ��>���@A��F��+?�?z����S�D�b���CSp�@u2�C��o$�.m�Jdx#Cަ l%\��q����g�����O���p|T؆~S�h��q�
t(;k>���A��d7���"&[h�����p|NJ�p�C���Q����v<���.H�}���A�� �"4��>�2��$�IY�8��+���� ��$��?�<d�}(�i�n.�)t,��45�(�"�F�KݩZ���^D�P����؎,ʦ��5j,~��"���%Ym�F�vt
�3:y���vvw#s6hg8�Nm��WU��Ҍ�A] i�ƏA0��e�Npo���L��L�"����
�L�k�����AP�",��D�]X�hacx��NBVO��a(Ҽ��R֥�|D�����a���_ߧ���)�M���#}0D���،�H#>��i�� ��A�
�(���5
��Un(���s�թ]h"����W��M�<���*�����L�Pɏm�$��q"�P��nnC�i��#L��3��;�Ӯw��>h�׾�=zso ����󏦓����cy�����g���b�H�	s+KK��|�f/"���Z��� i?�;�u0�#�r��W��g�{6=��@���}#�\�s?vx?���� ��6M>�H�MO��{�ݨ��_�?�������/xe��ԘQ����p�z���`׆�l0��Y���R�~+�'�����m���E?!��`��,�Zc񆬄s���C�p���h��u�|Y�{�jq�ϻk���������GX�t.�b_��N�cD�sG��ßX_�5�#��8`�m��y?��FV���g!�7P����'"�
�p��3��*t����NA6��{���do!z*DE���ڬ+&)
=�&�fY�����N8s�Zg�9L���@T��@�X��<u�C�����y�=W��q��94������Wq��d���%�T�x�ڝ��#��B@)���@��0��I	��s��� @<R�`�S+ {p�Y�SZz�n�̫�T&�6���i�;��6��,�#�S�"�-��9Ň*Bg�t�q~����(w��B���Sȶ�̃�@�كD�ܓ��ai��Ju��R��*�@);[y��l�hroV�yb�~���i�~���;�����IT6�aQjt���p�V�"���bx�z���*#�MSe�X��f��˦��2Y�1}���],��� 5�[{�
Kj}�پ�l�N�p���(�ql_iu]��\�΂�D p��'��gTFA$s�n��+�ȳ�v�!��%�5���W���FF��[�*�_����N��d{�L��Z�P���!!eeyTϗ�m��}�J�v�oM`&��(.��W��{��Eo�6{�e�Ca}�Ԟ�t���t����vz�߇��wd%t�Q��o�}�$�� !a|ǐ�� i�`�m�Fi�O�����\�.��;���o�St|���(�Y��I���`��"=�'=M[کt�� ���hR;<`�܈>ܤ��?{�aK��Q�{>G�x��QYb��̞�J�����H^�|�9�p�ǿ���Ty��A`�A��џ��'�3��ȸVｋ�{�b���q��/��1�'[�p����+ rƳ���ka�#*��8h�v��1x>O̟�$���;?�?�Э���ڳ�K7漚=VnD�<�u�p�@؋b'kP���_�l���N�<�`H�:Ƭ�d2�t��edM�6��и��&c�DT�a�M��+ȸ����<�,��'ݻ���@����iehYÕ}��0�#�u�0�Fy�~:b�0�{Z�/�
�Kmܷ����-]mP��Ŭ�v]E�
?Y��bTW���:7:�2�Ȉ'F�ʠ ����Ed�z��h�@⦑���ׅ�
n���Y������F�F&"���A{ L�0ǲA+�#����	�I������l>��-�Q�ލB����z��P�A�����������.�b��0�@mc�3�-��F]M#0\�y���U���ı�t�:}��! ��?�n�74'HT9{��J���MI{��r���è2�'V*��yؖ�mn,��$��ڦ��D�3�14�Qà�����
ύ =�����#J�hݺжd4Ks`#c�������U(�g����^%,�%�ĭay^@��d�K�3���/�Ґ�R���<:P�:����az��U�9�o_yI�S�E[�BۍzY��k�s���pUA����5��Q\���M�=Ӥ"��[�d�hY:$2��ޤ��n�=���qj#�O۝.�OP�+3���|� �|���xX�Tl"� T�M��2�m�ק�YYZ�8><��.��FI4��K?�Ŵ�z��7K�9�f�&0���w����:��:p.�Ƀ7@	��A������.�� Ֆ�q�w�Thݟ��3��9r�X�ε�i�i:oi�HX2�萐�3�g<�lbd�7�����XVs@��F��.{��Y"as���b�U�W�W�OAZ������5t]v����,�L�|u���gr����8����p�>q}{�#�C�Ĭ:�Y��.,͑�ѐ��aw����9ɭr��"h3�Bגh��x�و�o�uep��67Wu�kF幚!� �!;��8�p�u��^	�<"|��93�!S>�?�1z��
�6�n|����[ A����:e��?�� ��P����kbf3����~by��L��nz�����HW�K#za�@.4��o�uw��]�/�reN�z#��ѾF��z��H������{=�9��-���!Cfɽ�F3�2�n����K�%؆#B������
3h���1Ɔh� �Q&.��_�AgJ������[;��l�L����H��z��b�W[�v��"�i��o��7���{�`'��cG`$o�ӏ�:3Z����E|u�'}�{�h�@4)�4c�a�l��B�@bð�O�ׂ����U����	�L��RU�X҃��:#!s˧��*}�."9qg�)�~�J8	#�*j�e��ǎr ��]�_�#�%��������oGF���ɪ�)�b4��(����jF��䒤�$���i�x�|�ǳ�@&�6���^fԢ c4�iёМ���ܣ����x"�;���w��=LO?�D�Y��V�ַ�G�c8��t�*���{�v��I��p�.Uw��%��{�4��q۠]h�Wei���~�f+��F�Ʌ߾7����8x��>~:�o2Z�֯2�㷿�C8��z�J�}���6h�{c1Dk�:��L�:7zV ���xf�B�]:KDB��KD�A��ܹ� ��]��n`�/�܇.08f��?i��=w!���!����?��QO�"<ʄ�/|�Ӯ `��i�|��<��c�,���w.�7'�=�]C�a��t"!��@'Ѕ�m��c�/�oF���a�"ES��X�F|� �[��p'��������Wk9���a%w��S����v�NI�����=&�]�p��q=���'(C�q6��~;��Dݠ��:N��a�����u�a\�_εߛ�S89w0����-G�}�w`���ՙt]C���-|-�/��:�׍6E�D�L4pny��o�r	�:�NST�A�����H�]&8����gi�t�5�7-�W"�蟜	�r�D�D�b/���Yg�z��U4����U��Pz���u�H@��Zv<"?����E�p�E,�Y<�u(�ևS��R�Mw�+!�	�_����[��ro*:F[[��ܐ*ΩVԃ��2�(�����#�p�U�����?��KQ�:w�,��h:vd����z.�����p|b�N�m�k������ŵt�v3ݞw�'��
1�x�6f�[��t��jqv�I"��� ǵ#l.�\wn����&������(':�<e��=Bl��Xv�<Wgoս*^�\�ZMC��
'��n����8�0�UC�N���6eG��@���%k�&�5c�9UZYA���x�+�ʫ�%��r^�a������6�Չ�܌6�0���y�w\T�11���?�����NG]��O?�^z�t�|�v,.��?�����D[�ҋ�?��;{�'�>!�w��q:�Nw�F�ۿ�?ŀ����C'�.d�y�][�"����0��?=�R�09�3�.��}�t���4��Yy"���� z���-������\��XZhn/p�}�{��$Ұyɱc����x$���^Т���D��S���]8�~p1��Ǳ�nݙ֧���������i�=�y��U&�-��}��P�|�4�i�ɹv�l-M$bB	���O3&lU���Up�En%�M�$���ôLV�n9��Ʈ�3�����F�ZaP:uВ�������\�w�F�:�fFJ��v�15C��ԑH�}p�F8k5��6?vvfo�!3�Ն;`^>�Y�A�זIk�����5�{\���:|�0��~��Aw��{�@$tIuݺ����aC��R�$�^�)B5Gr���1�3�s�D�r�&&��K�p\���w�)��vA�Vl��J����L�	GOlRn���hiIe-�5\�����wx������N���%ջ�$��L��_$g\/YSŏr
��C��.%��|��@"E�gb���W���U�Om�	8,V3�07�Rb������2��f{x��;#8�V�1�yǘ����1���l�������(]��uX�F���PZܐ���������nݣԫmH�gK�-��<WV�y��l�a��#h�S��ˑ�Ng��Cx��|������9��r ��ψZ�Q�-�'�.s}f,lK]�n���*��Mf-��I�B��Zd=���������/�,�GVN��*+��̤��=tx�묈|�oGO�
��$�Y.g-�O��c�c�B鴄��X*M��lb��A� bt�0�w2��z#?z,r�����ӝ[7ҋ�=��"ߋ����-����W�h������O��D���>BW�u�rHJ��p����W��jL_3��2վ��_��U��%���4E���%�t:)!���#F�j�̢�eV����`�׼8܎��uo+��W~/�w�c.��GOГz��=��J?Bx"a@����1��;����?�"���߭��t�&��t��.��$�i��t�@&L�Ds�Y�f#V=B�C�x�DǱ��;
���}�U���Q�r�*�F�� V[�b��*���3h�+��oTgh���1H��Y���eHf�|�޽;��7���3U�׮�� ��A�(�1D�"��1��=H���q�c��G�uF���8��i)sǞY��Ξ'(�;������G&v~h���y0~@=�g;L�
G�ja�m̺0��w�s�ߛ���,�
H����ӧ`��`��.=�#���e�~�x;-o����!����Mp.2��9׏NN<�I^S�f=�s�BNdl����JF=*g2����#=�w� ���49oT/z#��E1x�T\|&�r��nҒd<��b�����ԛ;c�����9��(#ٻG?9�ç��ZIo]&g[3�:��܏��Kts/]��L�r=ͭ�E<�-r������<{��wQ��˟��s��V��2���g<jy�.�朢	K�7��7Dd�r��_1�H���{������N��6ca��=�P���G�֫u�&.�rbSDUYɆ�ז�]�����\^�P����|c�ge��ZF<�S��C �\ͣ�����x�U�2clC�B����su䄉�Ǧ���(�A��w`:}��X��W_al�Uƕ>�N=�(���LG��Д��Ё�fT+ghA���O`�oG��g�|"��|�;���$���215��k4��|�m�{�=�Tc��Q�*9��qmsvuIH�s4��.uP��)��ӽ2�;�;���!�Ћ��(�e?��_��m]N�<'Ym��w�ʍ��k�s��w��3��~�!�1��{dO�z=OP��eX�0�(IE���ɐ�=F0v,S�1�&�ڽ_�{��B��:�r�����A<����Z���u�n���������:��D�NZ���A�;�'OF�!��X��k�15��"��ӧc�mo����jz��+�7���vY�2�}C8�:Y� :Q͜��p��b���\RVE�q�dG<�@�V��E`lܓ}�Q	ע��J'�c�uz��{O�}���@ڂ�"o�뉮{8F��8i;����A�γ��d�-�8��q�M�&�#���YƧ�A��nI5Ys�`��&��<��������{�-�MF��k�ㄇ�����YEϡ2>�O�'��Z����\)>g����?�Az|`ԣ�:3Ғҗ�@�؇�L�c����>�m���������C����0�b������CE�2u�M��`Eұh�n��Ǿ�ɦ1]�FD/b�@$�bstl�wK��Rm���Unz�SE�|�����z�18�����aZ�a7�}72<�܉.��P&����KS���W���;!��/�����99�*��Ȟvg����=��
���k~8>_p�e��>��v������Q��<6 �5�iD$��.F�Un4�N?rA�41���	m����r_x��K��s�1��ߩ�Hw:q�D��'_�П������(�1�3zy�շҟ|�;��Q`1%M��%?7�\Ow6nS�l�=��k]#"'�߻����@�*���W(��E2�\*�D߂p����<9�=�������;2E����O�yL79r����z�c�Pi��q��8����X?7GE�:�~�.e< ȋ�B��AO����e��j6(y�P�����S;rԕs��YH[G���0,������d磏���g���r3>�Z^XqjJ��w�]�r�UI�rb�TFGgϩgN�k��RF�.���:jM"��1}W����4�F���n��j}�pƵv}v��$�lУ�Se�;<��;0��r�[��p��6�;\Qy�X|ǱN7Ea��~�J�����UxX�c���6�����Q��2�\�._��M���K�}�\�U��j8�̛���T�s��^��*C����x�����3*7�/G�!��daf'�k�<�̉�qs�����]XX���0���c	�#��O�Z���`л0��]l�c"td`��z��S�?�)R�X�5f�I���9T�M���a-��N�nE�9JeQP�m8��2;Dh�����=�5pvd,iՈ����Z�����z�����؅����U6|��,���Goǹj)W['+��wB1�"?�sN=��{$�Ă���+w�D��9-s�:��#�9 aeӁO3K�s����U]�����|^�;9��>x� V�e��T�*�0����ʴI����e�ixQ���w�yV�Tٻ����"<�T�A�Wh�ڇ����^���>����Z�I����7ކ47�����}�#v6��r���4�y����W^���PA��O�	 E��5���j��MJ� �շ�`�9l���E��;V���tTp����:�p��T�_��g(�;LT����ۯ��:k�DGP�An|��EW@�VF�ȉNd=}�{����ch�Ҍ�� fņA_� �ʶA���	q܀�JU�sސ=0��p�S�y����S�r��j=U�6�!:���笸3��y�Y��1���mB����3���Ig1b5�μ��b9�ߧ�ߊ	T̌BR<	�!&��0^�}Q����:�����N�� �g��'L�/��N�;��W@1��,�����=�l�G�����`�ee�w�6��3� a�)�B�K�6*�s��7b`�|p�\�ѱ�#8g%]�v�~�4r�D:���c�+kd�VŐ@���Xi"J�>;o���k%�]�*���S��*_x�GF�᧕G�}��W��B��AB�9ɜ�xs|�����s1_�ȡ�8+��vA� zF�*�K7��U�����{�܄������C��y�����Fz؍�#�L�Ƚ�BpI�ǅb��#*��v4"�ګ��,�Ie�����bA��9B5���$6��Lk@�Q��k.������jE	7R�,�݀�9'TO��ig:L�����@z�-�N�f�=��lO�#R)�8��\ܒ�Ā�ܐ���{�9�������&׸h]r�\����]U?e[{f �Y��ʌ�DB�֝�ˮ^Y��>[������85���9d>C)���n\e���7�Ï *�^����O�lS�x.���+� �gYK����(��i�Z��p��\'im|Da�*����fA�~n4(��1���@?�#�����*��೪%��!D�f��W-}�� ��H���3L������R�o����Tjo�%��Q����*��cS�H5i�@k�m���s�' b6Q|"2�:'8>��^wJ� �+��1g���c?i���$�h
aJR�m�o�IÔumg]e�e���R)��?4�Y!w:�uT�e��]�Iվ	�?V�Qn�~}�{͙+݊ ��~�\!�<�z�˙'�Nئ����<�T���^����ٍ9���7ixt;"^�"�̺W�UT-�56y�_*yT�����bLj<���3�7_UE�_9�g����S�q=љ�����`l��Rtb��w��1ཬ9�� s��4��_����Ѿ�N�

�E����r �-�p��,�2Б�"������f�iaD���k���2�A�
LG��"x��sّa�ǀYt^3"�<w��m���ܼ�F�g1H����\�^ӊl�%��^��'E��w`�D�y��D?D�����6�+��<���(6���(E�Xfh̝�4�"Q�e�I��zn�|7� ���š�7W����G�0:��%Nؕ��.C��
jx���Z~�JFff.��j������#����^�$:{R�$�p;-c��$+լ[��+�"_V�0�1ؘΛ��7Pp}||�#���UJ�~�Ыt�v��e��0��&N��]�(��%\��X[[F�[�x/g��OP�.������Y!𐚊D%iŅqa��LO�>�����s9qЌ������Q�(y��~�Ԗ�#/��y�0�E�-��_���.o:*�]deXUu�Mt�˽�EO�:�'�{
�����?�ĉD�����W���w���f��=F{U; jX$�<j	���ko�|��-"�z:��.�=��=�}��W��^c}�ZE�8���h��z�o�!�!&�� d�ē�=���^!�aJ}����%r��0��z�Z�.2�n!�?��O3qk��R����8߽���|�|����a�4@�4���!:ު��Ó�ԇU��L��Z��:��H'���X9�<�NGC���u΃8*vb���"
s��SM?U%�UE�L܇<N�P�mR��C��'_�x:)ν:q�����\���2w�u��W�Z��e��c�����O=`��r�'l���gL�䎇:9��R�A�c�s��Ge�#�w�Ȗ��&a��K�u����z�)�².?a����8��L� ��6�m�{��{���D4���mrYo�/$�Z���MR�C���dnBv���������2��!(�j�N���e���Ι!O�����
I�`���)�84l~P�T��f�	U�,�j0@�1�|�~x}�hܻ{Z4br'|ɇ|�M����u��7/_e|�Q��Kn>IsI��1z�x�uGO������$6�T]p*L��c�.�M�RjU����xWRq06c�қ_�1��9�pO�$&��ػ�m��Oe���>[�0Φ|r��f����K��zoTrT�&~�y;ޯM2r�'�gE���l�_D]�kV�U�@x��<d'ō��������~"�)*
��9��g��]kN�����T�0m���5�}�א{�g��<X���'��C��o��oR~8��i���<s�Ӕ�����iﾙh���_�ٴ��1(f��@|z(���ϒ�勃WW��s��5�����K#=rpo�s�\�����rg��6D5[hv�s�v+�t�γа4�g�<R*��E.���}������@9�c9G�O}�3��'ǁ��0b��̠:0�o��?������1z�?��#UyR���;\Wo�؋�F�L����~��ڃ�DZ�t����[x��Q"�����}Ϝ�xl��P�9����עL�E针��hB>qo�>��������Jp/�1���b}���(h��J?�Qw�屫���uHe:!F�ƛ��N󘈘��N���\f	��1E#��{��S!�e�)c-�2ט���or���0n�Ͼ�zD�y��g�d�v�GE����1�E]�a ��>2r�7��H9�;)�%����v._FF*�M����Rb��i�=��=�#�>�v���V5�IY���W��N���\"��$��9�t�%z}T�x�����M�}��i��+"W�A�m` c3F��t��n
nQD�o=�7X~o��`�	���d=S!�ٽ���2�to��R�5J=oA�=Js�Q��V��w�R�I���!����d+<��L�z �A'���\ۜj��vix�)��n^+o0�R"¦q��Q��n&��m�����=�~�?�<6�C���v�7�=L��##Мc�SU��U�gD���=K/���22��5��5>�V sw�S�;+�e_i!v��ߕv��.���9O�6�hW�b�U�|�{*�:o@�5;��d:�';���4�p���_E,�/vf'2�0��:Vt�2�y"j� z�1E��^��D5�K:�܆�r��vb��;�g4:~yO�x��pxV!�&/nt�3܈�0=�3DgG��ƭk4~���a�v�/�����
t'�	��NPw��ϿH�j:���\(���at8�۾J_�e��u�Ɩ�Q���7�z4r��>��:y�<C~'��Q�H������1��ҥ��������ν�V�'Ϥ=�G]���bf�,���xz��gXd	1rO�\��M�q�f2�~,}�ܫ�3���~�MӐ�"�-���ٗ�L�	��L��A<ξ�A�x}���{�[��׿�o�ЧH��M%�7�u �j�(�[LU˨���Ԙ+ha_ｈ�#�Τ�\�.�$�aV�ѧ��,s�����Q�[�*�ؽ�t9'��X3���Ǟ8��x�D6��äh9�C�҅�OV���"��f4����� ǏReџΞ=O�M�Sj~�j�^��;Nx�q:��p��\ّIpվ���2�ɹ�<��=�EO�)�㾈���\�y˾`m	)w����8c�{pY�8�ΤXY��w�����G�3u�	(�&�<w�6�����i/e�Q�z�Ug���8�a�=�̯��Cu䫏uQy���_�Z��#b{[��z˺!沮O.�Xx��0��>��M7��g���O�+��!��UĔ����v��£���Ҍ�F̬�<V���"q� ��� K'XN�&�ue�\0F�14��25�2��W�8�
���ƊP6BL}�L��S�8CfC?�z���R��F��Ӽ�s���vʛ'� *���Zc�:G�Y��66���q�\�c<sj^�d�^Lw��Oލ�:Ƽ��$d��#�/�떍�4��)=OٵC�5'+��Ӷ�F��(���!���^_��J�J�a�g;E�i�s�������t\3M1��=~�P�E�_�cXI�t���۠��.�@��]"�4`�{(9s�N�����0�ֆ��]�z>���l5m,�M��ۿ�W�2��l����C]�a�F���{��p/�9�#N��S��ؓ}��XB��sr���>_x��������9i殹x���0���|��t������a�k�+i?��Ǟ|T
�HS�����t��Y:�O߄D8	j2̐�	j�u<��>7V���ܽ��9�pEkQﵭEM�X�o�ܞ藞SP�|�<�F�[5�lU�fX�hm�i��a˫4���u�i�KT���h�i�{�aF���Y���pax�(i�ҿ��c2�u;�T�"�#�FbV�
|�\�!$t��ѕ��4��Ng�r̟��'�k�x����-��������Ty�d9o��\G�0��5���ӂ��$�'��@0��}{銈,u�61b6��V�L��ƷM'9;��]��o7���Q����"��R��4"�7��C����\3�BʽXom;?�)�6%���z.�HTܛ�;��<T�B�K�Lv�z&�z Q��^�ϋnMG_����)����T~OF�2A�~��3�� �[b�i�]���q�7�х{�� �n��*%W-���Cd�wz׷j̀{5Sz�n"���hّKғy^K�r����܌ja廜�Ю�
N�Dr����gr��e���4Z��!��&6Xz���������+��+\�L��(8|��l�c�g딬��.e۫FN<�ad��U^mؼ�H\g�#�!d���|�I��"w�W�һ`����1ר9)��~�^��4p��޷o߉}�zn��5�,7����N��L�%*3��ԟ�o�FqF���T�]�M�՛W�+�~�aY��`������n�Ay�մ��,+�q|�ľ��g�A��8���5R�ְ3�3�R8�C���?�v R�c����F׷��qbRTUde���i`t��O�D�^K�����rm���̜t�A��W����?�����E���0��j|���v��W��t�#Np{.=KıB��2��ƨG�vȈ9�l��aZcMi��0���V�^��� ���a^��w�UGe���xUד�x�f.��\���^��N����bY��A�V��%v:z�No#�h�:��$#j�W*�ƿ|]΅ǎnp�1G�9��aSO�@�b� �G����h{;<2��6��=06�D�;�\%ne�F	��H��d$s�;w���1�<cT/]�2�^OҨ��k�+l����Q�X��`������V��A;u�"ts�}C3�I�K����y�Fs�Uk0w��с�B�;@��M�_�Be���M��} .�v��6�ݻ�:����،�>���9���c��*�nm�!)I����ʂ��d��y:9��r:ݔ��oP�Fi�h���_��p�\[�@��^��}d�'�x�5k�u>TU�Ik;��\�:p�|?��)ҡ�!��m��>���C�?:v��3�@Vԕ��%w���aγ�OF?��b:Pp7�p�W0�9_Vh,3^,ܜ�	D�Y�*����VT�BCAt��m,�]lP�U�����2�ݏ�>����q���UN/�E�m��r9��(�.�������o�`^T�~��mY�v�y���-s�*Ԫ����ݎ[ű�$6�p�"�-�f��"��%��g������#�9��:o�v:56=��ݲ�Py��F=�nA�@�lA�o^����׾G�mO4��x�YF�j#.�֏S�"W�L�F����"��)Ubf���d��"����`�����~"��ܩ��[o�{���W������G��Q�1	AU��s5񛪈ҿ��s�YAi���Z�����J����~��`��4|+��o�)��'q���L�1�w��)��u�Ht3�U������1�O�!:����i��;��`y��ōk���Z�=��9�����VV��=�XN��z���(STũ��r��N.!��*gV�1T'��i�Nw4��gGT�-:�5���,5t�i2	M��r&y�-#�����|�e�a�������g��m�o߾��x� x|���x%��x<G��i�$� ���2��*������'�y��tz���A�He@��Y�Zx���2F��wD�Az$�M���B�Rk�0�+�8�D��ip��	s�7q�MMeҠ����u��Ȉ��#Jg����qvGA~N�<IJ��{��Co����bOLl�y�.�hG�,�auD����࿄!6�s�s�N�0|>��R��5�x���1P��`91�j�����Z/Q����B)�>��1�zf�ğL��] Z�Xu ����0ʬ��A}<4����=ֶ,�d+O1"L�ܬ|\���'y��^�s^u<Q�Jt<�Ji�W��>��Ex����A;�r�&ǥ����v�r�F�� 	�!:�5�@#&��aFw�~q���+%kE�<Ɨ�AI�	;������r#�|����!������h��Fj���yɡ�Sn��|�}�g!��2��_�x)ݡ�:9m�k�C��n�i�e�l��^~�&�P��dUO���Ї|�(��.ڵAI�6��'_�z�����)�sD������ݝg��
�|�ȟcحrDaF�J��z���۩���tg~�{���;�+�d5������Ì����#�NyM8V�֨��/���P�\�����t�����@�0��o}�[1(�5o�O}�S�I:�E-2�W�thd�(b���4����=���֭t��Cm{�6���;�������R�iQ���fz��7 %����G�o�
܄W�5��v�����M	�~��)���ʱ����Ga�-�]ű�A�f��鞸�9����p`b��:�EB�Q&���/׍{�cu��e���e� �?oC����[U ��g@9 ����q�y���C����h�kt�T�w�Q˽"J���8u�T����v��`Ȼ�5(Ά�ꢪl�	�#b�,rR��O%�Ÿ�j��%q�������_��ݼy�gv�:�"���>�qtC����-Ċ�X�������@�,�?p(ƞ�q�LL�q����=��R��{8��_#��>����=�!��{4��%���<�.G���r��+~:v9&6O�d�T�5���>�1p��Z��qo��Y�(C���p�n߼�=s�* +�q��Sʺ�A����G4���} �����zsd{�5��޷�|�V�aHd�g8.TQ�����\�QAE�w8��#z�Е
�u@Lya����.`��3ѝq�전>B��\��H61��t~�R��s��;���5�l�ةw�܇!H��(d�f�s�Jиg�2	$"P��弝LV_������%�F8G1Fy���۾��,�~�4�H��6�O,W"���(���Q�K!j^U��ёp�o G���K����(��/s�{����U �{�΍��P�f�,�I=���Ŷ������u��u�r��j�NR(��A����qZ O�&�/~��4��>gڿ��;��D~)�о���G6>2�u�$����r+�[4��mm�
������'N�Z�D�k_��{�6���F^�����*���A����~�k�FIΥ;(y��z�V7�D�<}8������H��_���,�sm]0�q�������O}2}��[����c�ƹ��&�K��3�r�bz��m=��\<s����sl3�r��ͮJ��k����7��#`6�y���T��8P}B�U���a���ltɑ0w�~׶�QD�D��i�+��:�F6�=���N���s|��4��=~�h|pb��2\��;9p���H+ؒx��Gi�j/������e�IwVh,1��W^#�s�>O�� &�  @߿z�%�r�E�<cxWWX���:�4jqo��c��Q<�W4�1�䵍��Q������V _�!_���L�o��0��pY�Ni4�721�1���>;{�lZ�w;}�/��g~�i2�3��@<ۅ῞��!	�[�����:�a�ÜD_W�J�u�Gu��J?�U�&F4�S����Bh��D��^a��>��Y�RNG)�,M]B�����Ξ+�h�O�9U�;�Ý���~P���t�0��z1LyZW^�y��R��Zbmi�ss�
�*��X`�T3��s��s���y[�����To�����a�6� `��h�R͜��ߕqvJ��p_�g���q��Q�^q�$�Ԇ���mw7cH�4c�8��k�P�tB�Bn������b��%�H��R�9J��4�*��(���F�����Wc.Ԯ"�3�N��FG���*�W��U�v3�0m҆U��Qo�?�s!�EJR��]��)5R66�X���ܺP���T��wL�����'�Dc�e��m]� ��l��wD#�Ӈ2�(�-#�1��.�O��L�obh���{<=�{�y�_��o�*���P�Y���0τ��S���Q���K�^cr�ݯd/ۀG�A�f��L�r2R�V����9��ˠ᡼!%:d���b�{h�W��e�*�>������˫�1t�ֽ�t����?�7=��)��D�sN�Wg��O|�}���R&��B�m��a�<k���Z���:<N��9e�?�����/�wY�N�N��d_���[��7r5�y�㸹ǁ�u�c	��6`��TG�q�%܃N^G��#���
���rg�B�|�.�������KW��7�#�� ���k���v����9u���7�*�q������ud����s�3�k8k�������X~������$�p��?�K���͕�쉼u�χ�/���sI���\(�s�8-����8��^p]�~(�]G`��;�1r���Pj���Y!�S�|�Bb����Wz@�~V>Sv�ׅ�="�7Dֽվ��f�����W�B�ބ�rCx`0n=�J��=T���8	�;oE:Y!=���Ơs�v[u!��nN�d{�s���UD�`L�A� h��1�ܼF�z���_8x*��Sv�l��u6]�����X�kHr��:�4���d�p386`�L��	X�����ߟ�B:�Tb�x:�6ŀq����R���t�#sڈ��`��W��f��@�疙9��EW]E�ѣ>�Ϡ(�G�d/��.@�$4{�ˆ^ �Q�h���c�����yB���-���]�m�n�7ڐql�5�FLAH2B�����;i�!�^��D�^�~.a��M��oI���F�J�KKx��a"�IF�.m8"���瘔5Չƛ�+igdb�i|��E����N�,�:�=ޭ���T��}��f����(��R�v��8"k˞j[s����0"�hʽ|��q����v�zI���_}����uF���ޤLO��#����Z�^���ι���}7R��ƶx�A
�,#TW�G��n`�q�~��E΅��{��a6s$�ݢ�o���ƽ��^h"̽���1V=����Mk ��W�/П�繺CC�w����- Q��0$��L����@f��2G��GNEU�0��~�m��o}땪�RU������]H���Q�Đ��K���L�N�n��R�E����;T[�u�%�����Z�b歍�={���7���J�"tZM�,c��B��w� )�)��H佽�؛샚�hN�!u;˶�8��:D��$龱W�U$"��Ȝ�N�!t�"r0��c*B�hG��Bg��3�r-l�ZR+��mЦ�_�~:��I�H{�y��.`'���;���[�hdu��ߟS#��*8���s��\��0��������&;��p ��|�Y��誟*m�P M��|ti�5��Q���z��0H.}�~J�6�����ͭ�16!61{�>bL%"�Xe.*����Z�MP�D�l)�c�C;w�#�[�6�ϡLʙ��t��F+����&����b�Z�eF�1N3�����N���'�/_J��*j#��P�vF�F�Swʦ6'��ly��1Ց�$�P�Q�A���	D'�$a�rI�Fh%21�l�YX�C����U�[o.t��{d�˼�4�1�nr�d!	J���Їu�4c�s,��m)�{��t��T�'�wӣ'�{���/<e7�w6]���g?�I�?�z'����&��� �>r0����+o�M\	��nh-��/�җ���@�z��(�:�b4E�a,<,�1�]�k@h4�7�K��VwHq�KU|*������_���@�1������|��my.�X��'N�"�M�Xk$]8w�c�� ��v��(1�m��SGN2`7Xn�]J��o�Q�j�s����15��8�z2%��,�}���t#Ƞ��>������r�i�k��� H�����_������d��&�[L����!+Z��,p#kj�W��_�W�b��K/dh�{���o���?�/"���Fp_f?�Q�(#l1}�3R���7߁}~!]ۼ{�9�O����K���^���������	62�.Bg�"~ s�k�*�o���y�����1.��"���7�*�f;3�]�̙�w��x}F�����}�����{�W�/Goź�=�@���[}�S�;oaۙ��zq��H)�][���bE����r�}���>�_���;�O�O�g/�eV���mP��`F�L�I���r�W�{':��[Q���C��S����e�<� �Fu��-��:D����>����οh]�K��*����{�4J�U0R0"#��A�F'Ӟ�T􊸄�������t6a�&����F3s/�IwX���4lq��ш��N��J7W�?Ls��\T�N�yf(��+c6�cpUFl&�f#P�������-ꞷP�}���N�G�,��+*RHo� �|d�#��pݢfya�u6�i�U�g�"-qst�g��7�-�w4d�Ǿ%oY���������㘟q��(d/�9?�۷`�Z[-\xY���cR�
�s��(�Y��;�k��F��Q��J���{�3z׸�6��Ds�(�1"뀾Q>W�m�t����%�3ju�f)F���[0��hr�\�w�|�hMp.��ޚ��i�r��ݺql.=v��������=��Y�S%Z���L�j�b��sS�,׌���H(uv��U-:\M����D�C(�}����}�u3�޿L� �e�Gg���~`Rr�������T,Ҥ����sms9zD�`^[V �J���A�K��k��;>�D�4�	'�{0 )O�Ns5��7"�?�ǁ����8�g��뷙5�à�aCU�&�ڒÉ�	�O ���#���w���������N���sW��>s�t�C�C����~�Y7�����}M{2��n3,giy;���p�W)a޿E��.�>��6i��6dɨ��Xc��_A��$E-�k�r8�h	x� 2C�*���"`�k#Ĝ�nw�t�-�M���+Y�nv�<���]�Y{F�~�id��������0�w�6����kئlԡ4�� ��O��i��8�i��7�x�4��4J��C��`�qFYU	�|N�T���42�ѹ*2�x~.;"�b���&4�C���c�Q����N��o�L.�X<>��!��^��cjѲz9n<�Q�Cc��J�t����7�n���$���m������hT��H*o2�d	:�����qF	�1�10/�XX������S;0u�BnӃ
��^�*���DL�I<6��nu��jy67��;d���d�8���sΞ��N{%L�n�sf��,�$b8=r_y�Z�[��A�lAL3����;G���Q�؅c��ߛ�]cn�a>3V���!�k`��ڐQ���(�c��Z�񝷧'�ϫ��v�1$��K^�ƍ����(x�M�%ʙ�B��IG0����K�>�,p�X�G�<�V(͙�&ơ"�H ���"���ppT�ܛ��B^�I�h"��0���^Φ;�<Ɍr�A�qm�R��֮�(>�;�Ǡ���+�џ��1�ͨq��>��t�Ң���:z�<�8�����*�D7(Q#eC��Q�QyW�t|ns�4��q��>x -��$-ɗ$�__�&�2nL��������ԏ37�3H��;LΛk��ܐ���a�9���Dz��' ꑣ�fr�鐺�K�	�a��l����Gy2���O��Y�|��)�D��Zԋ��@F���e�?�L���G���VFM��Ҭܝ�}��q^�Y����O�_]�@�FS�^�1��=�h� e|���XA�5ʜ���}�W��b�򟥙.�y{��D��1?�@�H��%pի^A'>:ʹ���#��c'���#��Y�m����D�~б�wJ�&d}�Ϩ#N�㻧��9Ώ��EΣ���[��\��BW��Bz'P�wp��|�����A��9�� ez^7�Μ!ec�"����"jw���eԐ�4�}% ^�$���Iv���k�N�Є�φ>TḎ�Y�<��-�M,�3���*<��a￞�N�4=�Dd"�+�Wu����N����RK�jiwIQ\�
):Ё�Б�CA��`��[�r8;~�̴7U]�]�<
Hd"3����~�7��F���PY��g~�5�����^'(�%���|\f>r�;��F��ٵ�؃������ƍ啙0(�3��E�tT��|p��܄�j�Z�����欢@k�>��K�dAF7�97�Y�%:�9�s^\ղU��4�~UvIzs#�J�\�Ŝ%ȩ���N.C8��Q^��n�H�!�y�T��T����>�\�ש`2<�O��p�NaF5<gP˜���Bx��YB҆5bfW(Ց|�2������JqԘ�G9(�+X���q�on��v���@8j��h��Y���D9����K�n�5<��� ��=���KQw�~�g�P���>���_�J�w�ys�C���������¾q�9��thң�BZJ�а���Es�3O?=��Ю9�������v���!7X�4��g�@f�q�
Up��۔�T�$�f+~��ÛG��E�ԟ�|rx���az����е�����ps�
uʴ����`�݂��|/�_�[�=�n�9L־�R�y���e{A��4�
��p��eD���@�kX	�\O��6 �u��x�eK��g�}p���I�ީ�S� ]��ͺd�.�v�L$*�|�6 �S����q��~�i/R&�U*\���(�]�ڰ�Q�EzWQ�a��XU斲9x����<f�~�;ޓ��k�4W�;
}��Q�@ćcM�0���q�.0E�d����x�{ɉ��X�W��M'�lT&|����bIS�F�@���B�{��n	�{;����~�j��:��QP(g�ؖ1^�����?I�q���B�������(�Mj�I!<��/R޹�F<�{7��34��FV=zγm{�`_�_��T(�y4�'�)-��Vc`�<��(h��||�<J�v���}ָd�+���V�|��y6M��12���K��t���D�6�Ñ�.�w�&٫B�������2���k�~��7O?s���Ք2vS8��N�Z�g1օQe������ʱ�g<XZ�|�H��o�Za�딭U��.�,,bU��ϋ�b=T��˾-�r�xZ�S�/�e�����9�LP�!�� 5�=z����r7W'���&Q2Z��w%��c0���~@���+�|�w�����؊Q�m�ok��a��5�0LyC�E*C�~ӭ���J
��r�)��2�$�����<<|�k_~����#�h����9:��e3���|>��zj�m�{��E t�w#�9h�u���9B�6���z�ס����h
� n�+�B�۷|���JD�1iZ��q��>�8YB}��z�ں�p>aK�ȏ�ﴷ�k��'>1<��8�d�N��7�
�[30�i��)�bv��	��	����g�6�D�0��+��`6n.�lf��Ƞ��ʶX�6�0/N3�z��N�
a�
�u���m;��h����3Dv lK�4�&�g��^��^�!s�*�� �������_|�TD�!M�#��/рR
~AǫT�z���&߭g�:����Ɉ��`�1�e��	�O�M�zJ����P���g����Шb�뢸�:�]���
�������ծ~�rk9�d4|�J�l��#�n�|�֍�)��"R1E�,PsI:c
j��B���(���T�Q��q4
<�3�w��wϺ�Iń��J�A�_�n_�o�li���x�ﱦMH�� �J��t�̲>w 8���dD�`#4�%���d�_���lG��dUqD���!9�d3�%������-�P]�+�5:u�2?xe��q��b�,�Y2��9��7��;�J�Q�������Y-���������}`�+G�x�܅���&��'T���� a\�Tt�����Xҵ���"X�
Z^�m�,2?k��Ŕ���Rj3&;��n�FS�k���y���B��@s�jcT��[�j�Tv�Λ����b��&
�v�n�y��Y�:	 �p�
^�2���o#x��K(n�d�~ X�鵌�H�1^�D n2.�
��m��qL�&���sl���Lk	b��SbrЗಥ��zVU��w�p4�=�y;^(FBp�põ�'��z�R�f�eeW;��D��gO=5�c`��]�]n��C�J�x��3\���ԗ�:��y�?�2��dZ�1�kF�w�ߨ���Tw��@@^<�@�&Bt�8k`e�@NOe�U�ч���[i~2	�ε9�J�1�)�E���]{����6�}f�XR#�E�hH����$(�mÆ�;�q��Ls�m�6��O�g���V�f��wNCT2_���:�����~�����v�\8��;�8��ȁJ��8)�-���Fֱ-P]ɩ��x��Ž`�9���v�LԮ����?�O������o��E��VX�R��u�^��8	㐙��~m�b;�8ѵ��N�6�^:���?{J%N��8ƇD.*�ԥ�`7�Uk5k�cAl4�����x�+�c*�x̍�)�����"-_���Ո�������c��:
@C[�R�����n���K~�d��D�M�)־O���W�'�s�N ڻ��ä����{]�������?�'����I�i��<z8)�*M� i�^X"Rr�H�%���FC "Ax��·���D���^�k��#���5�S�څdX��*.M׌ �̴�ёwV�po1#J����t��-Ґ����Ż�ш	~��`b8�	��c���ZF`E��}!W����*��y����������O~a��]E��vZn�ƑTy�8��c��c�LO5�.�Zd.L�F��|�,?�>�A��֭G� !ͬ���:������hZ�wPp�Ϋ�����-���9����L\{u���]�y�V�u��%S�� ,���<�==�
����رɌf,���&;u���2=���\��m�нvcs�����;0��6�Q�·��XכһË�[|ۮ�����B�0<�����*8S��<t�=A�����-��tj�7���Q���
����'�R�n�E��_�o��,!4�i��e���8��[�p�O����}��%4�O�g��M	�"��֕rk;e7dp�@�X��V�y3���xف�2C�;�N2�;b',#2���-��
��1^�.����E>I���G�f�3�{`���<�p���R�=i�����&�._�1�2�f�E�!���m�F�8sb�v�h�}�3,<�
����'-� E�$��%���S���H�yZ�J�>]R�w��,�w�<���c�7�G�W4����0~�$�~h�%9"�mi��3�#��g�J]{�f;�	�k4k���C�|���'2�I��ly���\�Q��m �M�1^8�:���@Hyq��To�%����v���2fU�c��_y���F:F��@8#d��w�U�8�DFDƔW�:�ڊQ�)�Liio�4FUƞុ��ٞ��ַ�4L!{dA���:c�\d�8�z�Dl:�N���=ua8��%�^��i�p|�u�wX �֜ ����\���I�C��5���`��a ���}�y�x�&޵W^QNX�Wk�c U�� c<��%}���T�<6��7��'�Rb:%�FX��`E��52'n!�
�x�>�V)t��#��c��g����8O�r���V ���ڮ�B�buǕm�p�Y��a�W�]B�[����r�2 �M��B��@�ZJ��.Ű_NW�8�(�p\]@Y��XRѸ`Y�Z�IQ�5t�Z���I2�y*aTr��1&$�H��ROE��PEzji7��c�	�����LT���*���ɥһ�n(U�{H�β�bh�\$�w�Y%���$��ң��;�����{ �J̑�'<��@덳�6Jx���/>��':���p@��L��c����<�[(�1=w�<�gsk޹á��Z�Ks'�o�O����P&W@�K���$gj�F&؂dM~x�K̽mu9*��fm��Lx�e�nBO�9A(�����Q�;i��O=1>�;�N� @��78\<wq���A��a��.�'�~{���� �x��&���?�������+.��P�� �׮��wT�����`�\�K�w�����.�bVb��]��9/�C?�r�!��Է���~+F^M���Qk��Ͻ/�}�	���n�\�^\&2a��1@��ɯ�5C���X\��W���x��'�O��F�ʯ���5$���2^�aۊU><K��Ǣ�w�1�r���Ly�}�:\Kw4D��h�pLꕪ����k����zԦL)�r����6l����%r�D%���s*<���#�t�����E�d �XP����%�>�����I;����s�u�ԃQ�-��q�F�0��1�R{"M�"x��0?T^,
�����لe��.�k��Zv0앫�e�c�{��ks\L���p~�f�G#?i�ȍ��yQ'٤T�~�B_��JGȵ�D��}���0�/��6�lɫWn([H"��nc�Nccl��[���y�%��Ƕ�3�_y�����~����]����O��-�լv7K靮CK1�:����G�g����%�W=��j)3܈�2g&zSkv	��X�z,*-��<
��+E^f��׫+�5��@	~����0���*-<צ*����}q+��-�w��+7lj�Oᚐ}ج�5��1zPe!+Nʤ�-�9�#,�}�;�U�� ~�0��M�bO�ڋ�* �27����{z߆�7n!�ņ��L�$��'��%�%�(9p{��@hNH�Bn�p��'�[��o�]�����fix����f�5��-��׹��P�T�8&H��&��~d�ZH�� 6��F��ܨ��Ry�kϽV��)���]#=�RƜ�E��8�Ǹ�0�D>�^�&=�ُ=2���X~�:��ɻc\|�+_��<�Z��?}8�i7ф�u��cPt�#��ɑ�|v� Q��\��ћ�����o}�ۑ�W�x�1I.�0j����S���!�'�}��j�I�$6�W_�FO�I�I�dSP�
��D���]��)(t��rҘ ]$� \ �\�r/ZFI���������[O�"s��x�����R0#�(]��6�%�*%���$��0��mp��a~(�Z&���m����L�Գ��c�i����Ch�{�0|�j#�]��Vx��m�)3E�`l��a:�:ߔ�73.�p҅��Iz�d�Mk�Y�}���+_��p�=D.\+J���FGa�)��x��)X����f���f���!�7�r�̕Ke5�{v���Ҵ*�W�qIu�i����!J�(��x�A�`q\�?y���+SLڢq)J�7�`��S�~t��_x�5�;�OS�_��
�{�H�q���A�J��ߢ����<t����_�����N����GLI�D�R+���Va�BC\��Bw�ּ���]	�߁)����V�H�\e(�u�P�z�-�%��6j������k��P��0P��!u^D�h;v����<�ތ��^��b�x�mg��o[ϓ�U�Z �p�\|�i��<�PP�}��A��,��Wv���q%zj�7xm�0,�}�ӟz���ގ���n������ �!�v��e=��-йN"ף�n��Zw�2���(�D��?��'��Ƶ!�BӒ�I��D�O�?I{�9�������c�/�s���f0�(�J�͒� z��5��;w���g?q�����c��L�hT>y5A�y�5��$�C2�|ψ�mČ�	'5A�o����3��N)�Jғ�������a�N�M��p���-�����(i��۷��ӱ'��m�6��l':aG6��pϮ�i.C���Umt���Ȯ~خ����p��ùc�������e�W�����D�KD����Fm���Yd�^��4��Nb�XC���x�x�[�a��m]�L��rr�s��w�v�&��m�u�p��2!b�ph�+�q�d1)Wm�l�a�2���B���N�m;�O<���ڊvZ~<iA���1��
\ov(u�w�X8��	��V��Pm���T*��> ���<W1,�s����hqJ[_ז�O��jW��Z�B�Z�[\���[ ���։bg��pΞL�9��5YND���^dYK�i�濍8����0��geLg�3u�J�ƾ��-��,/�(�
�Rk�jP�b�l����ޠ�dR9�翎����t��0֯��p�����c��.̽{շ��p��f�Qj�f	C۰���[�зl����w��k�w_~���$N��l�U���%˺<�0"��V�	aC����V�YU�1d�<�N�Ŵ�XQ����0��&w�P�D���Y]��,�p$ǳU	��뮞Q0h���X�c�k6���_ee�0W۾�H�(�2�.h�RD�x����u��M���~R���yE��uF6t�a�Q�	!O�2F�(EXM�W�����a�4t�/���V���=����?�j�
�OB|xI�7oC�/S:�)eb�jl�4k�1\�%����G<Be�2�q�W)�Zo�6vٻ�0���gO��0��8�P���?s��u8��:ӿ��"��9b�IGx����:����?L��4���u���9T��f4E��;,O�&�J�>5S�ݔ�P�.�͠�"%��o�'h�Ǟ>����/�J���TG�ݯ}�K���\��7a����Dr�S��.y�s���:�w�(���v;~�V�G��<����꼝�!r�OS����[#:�^�u؄C�_<�q\��=l���wE��!h�2[	��zܖ�i��� ��>i��:D Ԭ�� �ÆV����@�u�dp�`z�l����p׽���?:�ѷ^"C���f��nlD��(=uC�2ѻ7�S�,��,���TK|�}�a��WJ�0����N�MˈD�&UL��P��x��{���"�g�QD/fm��~���S���Q�c�#ytx�����������I����B ʠ�d�>f��+�%.��E�q��2�?�Iq�E�V$�A�L�)��.�D�b�G�3S����?]�k�EG��<��M$A�կ�9&�x�r�����YG���K��4Q�H��%�������=G)��ĝ�O���w�и����EW��w4K�3�R�{���x�{�|���G��� �InZe��ٽ��5Ž�s��y�wֲǨ�U_�U*��
�o�R�ň�*KH
ei
GJ�D���X�k�O���/�����ԮL��S�{��5u��nk3�͚�4��U����_6��\�2o��x��c������q]R�������{e���+�&-��9��q�ׄ��"*k����F�v�4��$�|彄�S�Ns׎�����?��%C~v�j�������h8r�����(�q)<���F��/������<�|�&$SX��U����CI���7��h�-v��>�9��%r�o�x������?{f��W??�s�]����3m�̋��?���{�Mr���m*«E5���F��<i����>�&m�a+�b��ukC�RBB�g��~��/��}����cg��|c����[�;�ޢ�����W py �>�����W_(o^��n1 rw_@�|���"U ۩8x���<j�(&s�7{!mI���xſ%;O�9�!(-+��)n�u��%5q���VR0�8�aX���gO �˽tB۽�s�Ϟ��"E#�����4�y��=l=��%h)��"0�I|��6�a��l�pN/�J �.�3Ģ"&à� s������Sy�t�.�|�*��0ȯ��H׼�(%"oi�J�A���?�2�3@�%�{����Ç 7�X��p���˴Q��P�����B���V��R��
{(���J�X�1����#�-M�W":������҅k2�7j�g��&��Y����;y�"��e�2���Bq���q����uu�5YX��B�wR1�W�YƉ�B���֩4��$ұ�$sc�@இ��ި�u�r�Qƹ��po��3�k�Þ��U�{wm9���?�������;R$�ۍ�̏W~���jG+,�{_�e�zy�	�6����j�r�}Y�1ݬ7Uv�����	(��[H���:)p
<g�iҚ$���Gf57C�k^S�#��0x���!G���1�sݖ	
��M<��w�G�K�Q/z�3�M?��K ��s�3�`a#�3�����R:��!#��g~��_���XƽlD��s��!�;���c�B*��`F�z�ό�}�ci}zLj[!ZٶmԔ/�` P��a~^y����{� ~�S�/r���QH�ڥ�=w�B����e���,�kMX>2\:׳^'c��/~ƶϣ$ls�n8����Os�i�f�9_��?�좘��⪬�{���m�7"���'�D���V6�]��)
~�o�wf8z���*���^#n�&#�҅m^�������/e�����9X�^�zI7���������;qb8��4as�l>v��������K��z��$��e	͆mZ2N��3��,��
}��<9U{ �~�V)�5d��z����CQ=���o��o�?�di�{�^�#"��h��q=Jr��q���p��� �����KKj�~?��ہ�4�,�0��I���oL.�ߊـ���(3��NT(3S+�V�W�֬�:�k�&]���#n�WSf��{�H@�и=����/y��̺`�v����/�w�F(�]#L����w��%�5�c0r��,�*�5J�%E�]k�Y����-T$$����)�O���;�W��5Gc�	o6�jL?)O=?qz����_o
=NA��0���{�y��1Z��]���%�)P��a��ņ���c5O^CZ,�<^��������ڰ�ͮ��1�x�#%:A��߁�2�w�㱇�g�x��g����I9U<���s���p���5�Y�a�Ҋo���D(�n�D��k��c-���dE�w-A��J�N��1�7c���OJ�������]&e9�)˙��[���4�n��zфI�,m���4�1) �qC�l�����[u��C�}<�$Q���<%B��]���ᓟ�ܰ�/�ia�(�ؓ��m��wJ!k谾Ma� x'a�250C�Q�b:��Q���h`9��۷w �߆�� ��V����7�%�l�T���xQ��̅^ ?|  �^ji׏�Y3[���nS+~c;��_L����K�W�f��"͘=���A���Ͻ@TPʒ�%Qė.�^z���9�O~�b�,��$�n����a����Ry�z+ˤ�Zܤl7?Í^�(4��Q��3y�UD��_��%���w �}XU��n�p���p�<쮝	�26���/e
]�"FM����?:a�}��í7iȂR���Y���O���V����.,�N����6��OS븧P؋\�d9r�/��fHl�&��1���o��'��U���W/�?>9��֫ÛP��Zw=`3p$   IDAT ��sg�W@L\���שHI����GR�=�(q�e�`]�f�ӻvS�G�|����%j�W��H� <�&�c3F�QV+{�4\lz�r2�y�.\EIHH���Ű�J/_��h_h��C���-Q�D����s�6
�:|h_�yS����ktE\�f��zɇ�������p�,� ��n�<���N?���kF}�$ʽC�h�"v���E\E����Q(<wu�U���uu�a1�WO��,��~N� �}����!�}#�E��T��	qT���~���!�Ns�]$�˂��֭���~!��됏S�O>{���1���Dy��`Xo�`o��L����رuәO=y���_�z��.�!��M�#��4��^�9*:J��p��5�\u-�����%���Եqr����"����a�u��z+�o;1L��p�g4��k�߷�f���-]��2��ɵ&/�񻐚�C�O�y����� ;��#��	"�)�w�>IXj�*���>�R(���X��'�dNQ����o��ɒ���N���ƾup�I2�	J�P@v���[zQ��L���.f��P$S!�XG�}3 .�Ֆ��x��@D:G3����{(���Ո9�iǦL��s�]��~�>,���_��㝆8��u�'��ƅ�����2���w89P�E�^<:�-� d����C�_���c� d���7�S���E�4x[�z^JŁB5kb�e��hS	�9Q����zs�+�G���-�3�#�-s��= �1<�1�jv�}�5��1@;��N�B�(�����e8z�I��g>�����4�X�i��.�X��g�NtK��.�t�ˆ��v������7|�k_L�ȵ�X�D��(����}ï}�K)ۊp��ˍ�,aI�3�x�u�FB4��W>W���L�<p�R�Y�SD{6�ʄ�%@?��7���^��v�wΞ$�����o�9n�zy�:�r����/
C9Yb%��{F�]��F��Vߔ���м��i���>o��=f��b�S��r^:OKң�R�~6��K��$G|S�ԩ3�(cؐ�غ�ѫk���]�DK� ����LYY����)y�#������@Ύ͕5�S��5P
�=�w pS�~4>�m��y0ߡ��s�Oc�})!��}s�^�ޔ��9�������e"(�]t�څ�2GqF��LR\`�X!�*J<ӚXc�	�vK՛C�!Me�v
�[�/Wqn�
vv�3�s���M�J���u^�;����gXf+�֑��=w���o��KO3�����.�{X�gnҸ+�rU�ٔp�[��n�}}1�3�e��Ϧ�!%[��RSC�y�Y 5�D��S7)*�M�a�B�V`�5���$A1��U��Psj^��z��	��Pg�!a�(�Q	]�Ra�s�E&)��kž�\��a��|�S�L��	���g6�?��%����5�^sjfʜ��b�n�粘Y�q��w3j
~�I��aa-o�x%l�=�^�u�� �}O����E��^�
��;�E �Ea	tQ�o�]��Ӥe���xtR��g���ߖ��Ǐ#�~Iu�e�C=0a���}P�.�+�3������a���a�P�8�&���.��>�3 �g�tv�4���p�R���j���kU�W���/��ʩ7�o��!]C��q� �	� ���D�e4�"BO�G�<$�˩`@^~�C� ˗��Z��zJw2����w(���A"�|�u�*,p׮<�;%Y�� �nP5p�p��y� z�(3���݈�߶g˰��^<�}H�5=4�{��ݤCLsT�9덥��B�S��gݱ\E� �S��;�4v 㬰V}t�f�T�Ft,s����MM��=�=�%�ћuo�r(ίwm�Pǆz�1�܂��_!��@����$�	W�%�(�%���3�g�\�S^�v{=�G6o @�r���m���ڿ��3���0����t���*��|��!�q�L�[6���h��S^KU�p|tye�j�-9��+�ޝ�ȟ�%-�V��U)8���X��w�=����������Ż�h)��$�M���X�R `S���L�'0�&Ѩ�qN���X��A�}׃�Ҏ��bL�MCvc��N���S�S4�_!�b.�ֳ�_�^�^>j*���=OdpE��sy����y�����f��q�,��&����@�+���"$��e���������K�}a~��tr��D���圜�!P�pܧ�\�Mq����QZ�Vv&����Z}��t3զ���B^�ҵ���Q����5�n�W���lFØf[��	[ī͢�+��r(�(v�=>7)�Ǧ4��
�i��(�4��#xƳt)CH�=�k7�bl�M�N����>�ȣåk��}`-�C�[ o�^PP�Bɰ_Rd�^��Ԯ�s[��קj��
l�jyF�-(_o���Fw/{������\��z��Ȍ>�ƶ���ˌ'������ߊ�sp��t���������!�R��?}щ��aɟ�y����>?������3������C����jQ�C�UJ�n�'��8ky����k��x��w��� tS2�]��%�QV�����MWs��i��g����)B�A�kt��o΂!=�e~0RTl
s�3�߲�������w�G�/3^��F]�g!I�a��O�1���&Dy�����w�	���!L��庶�-MX�ߵ-k�P���}ix���׿��a���Q�B�v#,),�~	ı����qu�J����q�4M�,ˤ'+�y#&��W�g�̏�����5��^M��p�ܠ���w��4�n(︩:�M>{։Խ�B�y+9ߔ�aL�/ʧN�IҟbR�s���xQR"��h�}Ɬ�N�$��=��m{��)<ދ쩭܇��}�ꆅ��so�Э��쥌����Pi�5y�z��H9A�+�%@EdD�Q��v��.��&K.���,H�y.I���*4ܛ���'�޿���ZJ%����!�Iw9&�.&� �OR�'���H�T�:�K�j�rxb �4�Jvi�o�Ny��?���1_�B0I��"'�UvIQ=�a9�v.^G��&G⸭��������:y�FiН���:�� ��,�u B7Q���kM0�����dB����+� D����/�f����Ͼ����჻�ڶe���k����|�Y�Y�|1¬��K-��b������ب%Y?���:(��� Q5 �lY��Zzx��&W�V#_%�&+5��ZB������ZZ�*�7L�MKī�׸������*-QAx	>��3C��~�)�0��g�ҙ��~�7~}��'?3�M���?�%߷��������JjcJE�D�δIHVȣj�+�h4�'�rB�MIHf7��G�=\V�r�9�/�vlx�$%*ze�ъ� �=�����*m�w?m Q�����
'u��[�m5w��-��?��?E!��瓠��s�F�ʹ�\�Ar��J��V�[�.G���K��g#@�c����pe�S-�IP�y��Q8(W9�7m߭X�ב��G*@C�x 8m�⨨8�"��fg�ۆ-c`�*�OJy����U��u�~���a֓En���s|v�I#E�k��/�>�w���O=	z{wJ�ާ�t�70�j�v&����t[�V��}d��Pqz��yǍk�*aRk�mt��·���h��}O�a���s�'IL/�4�SY�G�ʬ��84U��X���]�z�f����w^SI�$�o%��G]宁gT�p�5"H�C��Q,s�c���)����¥�wm�wH�=GD�hɲ�!]a�K�G��rͨ�
x�fOڹ�u;Ѕ�^/?.Cɢ.��L<�R�Պ�=�_JFm���w~�H�|���F���N�:����L}P�R*H��%]!�`�E{V�FS�Yl	����j�UT��=�h���Q=�F��%���á8��Ð�<0m���^���%o���I���*�C�)��͒�g����ȣ����~]����ggΜ9���G��w�;��0���[A�'���2�^��K��O�����B��ҁ����7���uǮ}����z��g��^��JE^�Qy�U��|�ۮ��s��*�Z�Q��FmSb�TyQF�Ik��
�z/a�&L�'Ne�{��Q���d�T����"�L�eI��9���T�CKڒk�> ������"��V��!*�x��	��+�_����-�YM^}����?J���h��y/��-��Q�������ס ��]��6�1�d����9���}�<)0�9~��9(IסP���?��0�n�<���	�ʾ�Si�zk�Z&��EU0�P�i�r���pZ?��(z�P����������ީ��׶�'��硿�x��mx��8��MԺZe�o��@޴��-���XBG���ـr���
��J9�ETt��4����+p�V����e6��D��M-���eD),���M������TET�W�[Ě(�ϜuX�4�l\=��:���(QQ�z��p,�����~j��ٿ��9؆kW�%�:0L�x�_�b��q����DE-�E%������L.�֏�[�KC���3q�~bx
�)��\g�T
�5���������fW!������*�5n��?��Ea���q�:��Q�����^��d���*j7�n��+�y��S�� ��`P��|;������4����5�*��!KX�w �`����FH��f
$*�~��5���ipV�ըb��x�h$��M@a�A������8�.]:�:�+���g�Rr
 �c��O�%2v  _��0)�2�zym�%�#s_t��=ȝ�G�4�w��?���vqn�I�H�5m~��M��cvX�YX98��!qg?�H�2��o����O������M�lCf���ʱHxK�P���&�5?~bx�w��w��K����������^=1�B��ށ�a-��)�Z*Z��a�����^eg��?��|���6���\ˢ:�94=|Q%�O+�𼻕��Y����
���h��i���q���"�=�0*h�ɍ��k�(�<��@�u���\�}0�݆bs���[g��t��3i5-p9�}��7�W`esL��'$��1��иz5�p	�4˝y��l�QR�6��1��=�Ǣ^�l�����s_���Ly���)�E��� ol�4�����x&֏?�t��{���zX�.&�.��yʵ.#D�?9��fx�╋x�(h��' SQ ���+�ߢ��p�#�u����y��e:�� hs
��4h�M�\_�Z�.�i�L	Hm���lԧv7+p���x����5I� ���1s�G��*�W"6��XVS�<�&�r��v��t�T�(`1����=8C��0s�u�BL��Hs##��ٍ�l� pr�|pRx����N����u`�v��`=;OZ�����gZZ:&�M[��;aw5Uc%^��DՃ˘�xd�a=�Z7�Ʃ�� #�i��{ډ�d4�j	����S�yH�����ϕ���A������:ɕl�Xe�7b�x�brR�ǜz�@����#�]Z����C��F,����AX�~����X�{Ħ*0ĭ���M{$F�n*:�C�y⢦�ϖ�o���eZ]q�#�zİ��+G��%V��҈Q�z��ƹi}x�H�87����V`��#�脚��]�V�()������O�E>�qSUE���p�)���[�Uhf�t#6���w�t�4�j.a8�h���q�5M#{�Ƹ��F��y���qw��H��$N���˟�Kߓ0e�Ͳa����`���8�m�9�1��իsc����?��//8rd�ʆ7�����%�'j�Fb*�lH^�Xÿ.�"7���
�<(���КMu��X����aǛ��G�'��煐�Nu%>�@4o$�X�IՁ
݋�]��}�@d�ғ)O.����rb��K��i*����9?=<3Ӈ�SL㍢;�%:�i���کKo�{�@���}��a=1���ئ����3W��|����
$#�=fd�KƘc/�/�kq�5�����|��+�P2����I��N��)�Z0��G����pmx���ၻ��m�$jq�w��'��m�zʓ�06�K?���������[�3��w8��α�c��BJ�^}���_���߰$��U?`Z�{�K��?2����õö}���H�_���w2,���7�d׳�Ab�	�rME��g���6{|�0��+��(�|�<k��݆��`�`|�"ѕ�aˆ�Y�z{��	�TҘ|;��;{)���h������g �%-�yB�7�X&0���ݧ��vq}�v�Q������瀢���(^���r7�n��u眧v<�Fj]��.�x��&��S
?u�*Q[`�	(�s)��1����Cc"���@�4)����^�͂�gM�g�R#ʗ��� F������MR����i�k�Gc4��8�6j�ǝK�
�v�(6s�+�Z1�&0� ^Z9Ri�n�t9e>ηQ�	��@	n���y5ũ�X�f����u oL�D���c�TT������\C���M�D�8��K�Vj)<(�q��,F��=����OzcF��w��8K:�{��S�v�؅��X���?�1�	쿆���7�:B�[!��6Ǚ��@�h#r`'�4n�y�ell�BX1��:�ە��#�ޑ
�|��+W�����Fk�u%�7S�g�k�;�e�*���� 	�]�����7�?�%8T�0E��WCI[~��S!ބA̾Ֆ��a��vQ�6��@������+x|7�ӕxb'<ͩc��*j�i��v��c\�7*� ��ZK���r��-����٧ W9S�f�i�T�����)���QɋEl���v���k4do����/,�0�����-���K����^��PSl����K�\AP��K%J����>4R�6Jƭ]C$v��\���K�;��<�0��9�W��?ǂS`���\`.��֓��G#���
�/_��'oE�l ʰ9\C���6�w������@���Ȟ8y�\�g��g��ǟ��ߠ��������<ш�B�d�̟�Ռ.g_��g�3s?�N`<Qs���%m+V�-�6?v7��6R�Gͮw&�����dK�k0�8�m�����9kՈ��@ ��7�P�J����W>�E�4��R�r�{�H>r���[�AD� �8��:x/=�w�N���c�""s�����^j���KxY���R�!	ھ��1<zs�̉{,���3o;�4��GaSa��p�����)e����*|u�"@*{�k<��V� �|WJ�*/<@�9a�I2њ2�Y*oհX-Em�<8� �v�u��=])�� ����o&q{����}�Mj�E)���-\���D�d�xp��H�m��|(��ua�o$"b�}�X��˓��T��.����īL��z��v����k�y-2
�@���w�h]_ZEg�W�?^�W,��{vo�[��ƞ/�k97��7���p1{v#�� �i������x��?ל�er=�Y���\�r��D0����{v�[7|���sL���~���W�&�^� $�ug?�H�~�ԩ#'O�|�H	Z�g�}�k�\�n�s�K�IJȓk�6�6��<����+ִ���ʭ�{�&- Il�EBD�(�śsxy�@\'$R�&
��XS=��[���%c�;�E��$��4p�������Z�s4���5OKp�x)��WAf��\��2��xM��n�̳�F�e�bU'�[�\n��Jql7�����J��S���KM`� �������b�����
Ԧs4�0�+�ױ�4̰�5�цʧ��yB���T��Rꞡs��Z�]���F�	9�Ζ\��*�m;���_^y��S?�MZ6 �[��(3�&ϼg��?98xdx��W��������tl��?�6ㇵ/�6^��
䓟�7T�������_O?�<as��o��0�#�>1<�'i��8y��a;(�6Rw����a�#wSK|	0�ld֒@E�!;q*�Xza���[���0{~�Da3uT���0��4Ѡ�z�T��A��r�m���f=���qHtf@J��:���������$o�>�Y�BD��W_�P;9���Cۜ(��}[��3��/���0|�;�a��°�mx��	��a�!ް�3_��D�l����w�f ���xSU
֍��\E)��P�p�bK��Rajy��i���h�0��|V��2"��*R{�4���u=K�E9�Vl$Ǡ p����{7ǟ4� ���@���gs0�V���-�#�jS�4�߫&+�����C������f�=�j�ltG^�TwW���N��:�:޺���&��#�+�z)�b�@)p�aq"�`�h�YQ^�L�t�\U��C��~§|��$��6�zj�@�D��b���F)�ܽ�����lX�:<��Z�!Z�x-"gM�1:u�-ڙ�;{8<�1rɮxa��K��O}���U��t�A:�8��ݘ�ٹ#��������I+��O�}�cOgE�)�Z��0���J��^�Y�r,���az�aRy��� +ih��VN/�I�h^,����"�3�ۻy�N�3
������R.D�,�V��Z�a��0y����}I�����uLM��ܼ%��dֹ�mEY��1��8�}��{�2���d*��e�I,/���?<>~/����1/�cv��"u'���x}w�;�H��l����*�1��o��2<��e�ȥ����+Ϧn �[�y��+��� ����1x�7 �D����Bk	��m�l�R��r�E޿�k�@�ior}[�������={@�~Э�
vD ڿy���ã�?>9�o�s��e�;�?�$u�0�!�o���۱��Or�7�_v���������!D:#rnu��AY��-AZ�^f��1�)VÖM�v1�i̼9�����q�(�~�K�n����7o�����H��F��9�3' *�t��E�V�` �9Ble{��n7���/��E~�����X�4<���ý�>8��|��&
�j{��U�SC��S^���U�rd?VɢUU3o�Jo�P}�k�ʍf��C,½W������(I!�et�Q)�2���kz�r�e-
�2����x�B�=L���R�֪�M}z����[Qyxe�Z���g��c���g�Lm�5�%H5��>+N�D%�3�-�]�'�v���-���G1W�M��y���0������.J�v#��,�������h֚����U�2�6�W���z�y�Y���*'� �`�H��{�6�� �(s�M3���t�#�~��0	6F#6��ѱ�TZ�N�Bރ���r��q���C��Ko��2|�3������9�L:�$2�f����8�n�o}�[��A�_^��X��(�<�z��E��z�*$�Hy�.P���Sh{�fO�AY� ]���p�����V��`^���������˽B=	�!X�B�)�E�P�T1�L&����k�
d��L�*2�AJ���O��|����P����+�����������p����ٓ�-x]��W����_{��h��H�^��vj���z�8��`	oE=��iȴo �6�N����}�;�^���8V˝�97��R�FTz��8�����\)1���P���z��P�2���%	ḗ6��Y�v�x���C��#��M���`���u�@z��!��/�K�,?F�$?�n��'?����o|*�Y��]��3��=���{`�]8�#Q���?(_���(��n&���YG�b���%X<#��#mL�5E��%������4�'�ӷY��>V���w_}���9|��?�`r�(�R Nӡk����
-�|����oE%h��,|��vh{�8�~#8B�{ȋ�ݵ���ѩ�T=l�0(^�����u1AM�}�e� ��جE���T�,'R����*hhS� Ī�-u{��+��27�?Rѝ~��ձ�J�E	������f3:����X~�?z�^#@iS�x�[���|��gYثƇ׬7��ZU���O'R5�an%�a�u	 �����5��,Է��������:�L��H����R�f$�Vz�f�^]s9�e|�,f�IZ���?P�>͞�c{B=�����i}G��|ט��|-)PC�R�{������O�����wŎi�@-6�5��/��c�� HSeas�%��H����s���N0<S�dY'���8F�E��]���q
���an��.��Օ�����X-ބ�0�W�2�c���7gABzq�&�{�����^�E�j��ўoʂ^^�:���K-��!��Mc���Z�|$H�\��t&,����Vw��b�1S�{���)B��Kt�EX1NE6��K՘(�H:�����A��n�@�w��+�Gu#I����w���g>���y��~���D���&����B�*u=����e�T�8C>d��K�'��	,L��j�R���o�)$���a77�|�O����#�d3�]�}�ʟ�ٟ������2��K���>����j�5潯���M���µkW�9���!�Y��h��2
A:;Pdy� ����Sǆ�}�Gx��0���W.۶n8����ǿ ��hޛ��q�TX.�H��C���D�G��Q�+��9��� ��f�Vk�Qҹ��%�#�b+�I;�ɰ%"�҅�Ʌˌ���ު�����t�z��qx��'� �w�J_n���ٽ{���{�)L��fTqæ��&hUJ��Ш�DK�Y:��Z+�כ��@���_<|�Q:f��JPy"����p�K6�_)��0�5���������%؉<p6o��%����׹���!�p�3KM0�
��k7:���5�P�i�,c��uվ�7)*����J*+8��Kz����M��S���oʥ���rhL�.�
/z�ɨ����tS����Ys��ʊJ��/��U������X���rn�^���Y9���m���6�/�sߛL��4 ����-��m�L�D�؍1���dL�/sź��E�i��%��sϾ0\C�ݼ��)t�f��p��W�N��N�_�6�z�v�ǲ�m�RT%8F��d1
@Z���N@�C��<��
*��+ ��Ʋ+�,s8�Fe��u��֠��{���oi-������ ���cK�e�s0;�U%r��Y~�c���wNʞ�/��]��>�$�,Z)jK7�����!��%d���B���=Zk!2� {��
�K}^��#�w��1�ع��!�	��M0�i[}�����M�]�=�֞3ɷek��\��yqL�k�֏{�1s6�X/��(=)����T�?�;~��� �.�^sk<�����k����o���5����4���8\<w6�Y9����lۼ5���#o����֛o�}�I�~^�Y��s���j���O��?pee��7��~w���ߢ3���e�jo�;O����ې�,P�n¾I�t㪍����B�>s�Fi$9��(@ْ���Y(ry��D) Tѐ��*V	N�>}��ik���9@�=utx���Y3c���q�rܟ��'ׇg�{
��/�u���}e�C��}򙆹w���ߑ������F@u�]GH�Ѓe����
Wp�X�~��D>V�,���V�.�=�V)o#h��ve�Asz�v��;.#���VO^!�R��5�*�ev���s�*�|��#Q���s.��7!	�\B�ݨ(@^u?sYW)��H��}����*��[C�;^�?`(;2�Ej�ZY�)����Zk`3�cٚ _SEa�[uh<�^y��̀Lz�jR_	���l�x����ｵcf+^4�b�T��x��Jw6E�j�)"�!��I���H���%�[M!��A����tu�PQ�p�P��"�_:2���@�ۺ��-�jkc�'�}FD�M4��Ϩ��1��硳�& )8�l�rΆn4�2#�P9�� +����f���N|�A�����Z����5�/����c�G��[�3*�l(�"�<�c�Q��Z��
�y���'y,ȐW@y�����}gq�x�89�5̃Z c��+��j�+�'�h9�E7u���&��J�S��&�R�\�B�?s��qΛ�H�
;a�e�c�Q<����rs�Q�H�����Q&��L��N���K����*��&L��#,j.���n�S;�l޼���թ����+y��dx���1<d�CQH�b�����!1c�I%`�E�X����N��B�C䌽��Z�������{÷��� ��_�,�:����_f>��O������n�Ќ.M��frFx&�	9�,L���I}�JV(����*:�.c`w��>;�I[����E*�;
�G�`6`�,Q
D=8�w��i �����[a�ӈڈ�mH��Gxax�����H�M$������/h�r����ch�K���q��hﺧ�ʹ��;�M���C���<����:aޏ�ջ'T/7�)�
o��,�z��)k��O/��V�r÷���8���{��&/95�A����;��W�t�[�=|K#Ğp,�2�3�E�����lޏ�װ(��I2����$q,�0��≶��;��퐳�Vz6{�sf})�HU�Q��i�����;VT�)���zV�r_�m�5�|�xД{��\�9Y�;�-��5�qͦ����;�&]͘�Ik��X;wFO=��:	5��Ҡ��3���m���b�)\	���II�������|������#�.qx,��{`��B�����KȆ;����:�mP�=�ܬج�Z�k��B(�4���\f���i�g�i1Sn3��>�^�z@tn<��aF�{Nar���u�.��/ٸAʰW+'gs�F��1&��C�TaC�n�p6:��3.���L���~�B�s�Bh�ܪD1��$O�aC�J*f���Sm�״���	N�����`�������-'H�h�H�Q��ڴe;�Q6䖝��\;6�d�����9�$'���(�|����"d��$5�����e<���Y���s�s�����}������ӄ�(���tnnx��W	�����?��&�.ԯ��?~ix�w�	O������ �J�|�`��!�|��������ȼ�2������o/F�Eh���	<ѷQ���|���a?!�'{hx	p޷��x���x}�k_^��������!�g�PP_�i/TJD�lx��Ѵ��A��<(�D�<���f7�Z�y�҄U�;�����`>�z���+�0?����kg0�v ,���޿�����-�?Ex��a=�7o�J�����׿}lx��3����IJ��1���t#��2|��-��CJv� �{�!j��ʺ����l�z/�*0��.�i��h^���+҄�y�g]���\F��>�e*]�����U�w�v���qy��m��=�����_���0��ɽ��!��iŔX��*�g�L�I�|T�:��ngDo��*��,���cO(7LA ����L�-����
�7���2�43Ҡa�do5�X9���*>����.��1�#�w*�����c�Δ�
���(��(y�x�S�����u#/�H���;1u'�U@�6ne,6���}̋��$goy���D�\"�IO{֛�8�K:v1�����l	`�[C�����0;�%%��|N���VB���q
n#�"|�ee��T��s��n�o�4N��}�(,d�BA��B��7�?�gΖ�h���.��$Jgލi�**�S�;fH>��*QQI���JS����W�6�һ�s�� �;6Ӱ�~��� ��t�O�}�� ��S���5"B���{��d�����e1�6�/�{9�
T�?���҇��`Y����G���I8�}(˴���]�	y]�4����6}Y���~��5R��y�gZ�][�O�gi7��I�5��e����zp���'O�<�}��D�~�� ~aN����hs�h|��:��y����W>�	�{�ϟ~*|��P��C�z�_Ʃo~����3�������׿J��j��×�u�t���OS�n��[i�"���+��'ՠ�oC��v#\�n�����*S�V��a)�F%oEr;�i11ů��j���[i�J
��U�C����p��4�/,��8�>>ǜ\w�P<��~�3��=BNCQ��&�o��:q����/_^{��1;���'>9L������<|���&�����;��u\
�E#��ඡ
�B�F}k��؁m	Is/��C�*����[Ei刏B�WT*Qb�%f�h�4��Ϻ���<Vg��A��s>��5�G��{�}��lͻMN8�2؋;��ι~�f� 4��g�P�h��K>W��*(�t���7i�Sv��M��F���N�<Vs��f�M۽.�ȋ�߲���@v]���`��C���QR^�X������|�S䵷��x�Ց��YS���4�@�f�HsD�^y�d�-�����L�����h�w�>�޿�)xD�� Yv�ȡ#�,)7���J�-r0k���N��4沝��TJ�7��!c1ޗX��Ww�_�<�͔*�*K��E�%����OV�ц��#
�l#��� T�#��ɔ�n�H+(���n�e.�+������ G�T
� @1dS)�)������>���r��/ek���@����sj&o���j��-/�+��f(�Rи`��=�^�S�1�W��|��7J�f����8�T�#$~�6���D� ��qi�� �&����l�#�����(#�
^�)MKhl�1��!���o=;\#ל|j�w�xyç8fRֹ��'G�k�]X�[�>�uj6�ܰs���O>1|	������?��!���DAI�aLۗ�/������~��p󔶐���&�ٳ{/����>7�_��=�Cy	P�b�����q��˛f���n<���&�vָ���;����Nb�RY�~�#@��2r��a����G�R��'��/��
Į\h~FzW��G#'Dl4H+�A8rÖ|r�6S9����OcpyXtDS�x5���g]v���9�{�$nM�.��⇯s�*�'�)��uHe�Q�{��k��U1XX��x<ɋ�'#�(J�r��i.�[\��*$^{�{�U;^��]ڌ|:mu�m�T5D�S�֍Võ�=��yG�w��=���=g��yM#eP=T_)����~-Ui*K�vUBW�#?����9�ԭY0 �{����M���B/���D�zrƽ����7*��������7e��bP�0�qf���B�B�!�,-á��4���Lc�-��C�	\
�<4�����}��
��K�c���apY�D�^���w��Y�^m>36�9u�ʹ?~�RFJqSx��o"%6�!2������;����f��~�s7Zk[�j���4�,���8F�7:v'�/Ys��8]@JyS��<�Q�,H�ۿ�\����YңY���&r�	����#
���|�£�}��*��*@DJk!ZRȤd,Q�*�����"�'}�4MHT�+��ޒ�Mo�����: �;Գ��%0Ap����m�o���g|���BWc�R2r��?�5����ʖ�J��F�)ޣ���Ux<�8�G˻��}
�Ǉ�߆}o��"�ۻq���?5��'p��/��^y�h��\Ǥ��`� g-����5������_�M��p��O<����3/����3̓�Dy�dӪ8=���'?	(�������?��H4�x!`$n��/|���D��=��*_�	M��pFs����/�a����K0I���W^O��M;Q�S}���g��k�` vC�b�{�3�=��%��5� 4Ȱ}b|��]���r�c^���KYPи�`�\��B�"@� �m���z��.5c���??{��̰�0u�m��EVKM��FoX� ��
^�x�唧}�49������%l�;%�$��t"p�Kaj����Z�5�Df�hzs�����uݮ庽�^:V��jD�y��1���d�,�����X�ʯW��iT�=z�Q�1�/e_���纛U ]k�2���y}�d��yN��x�8˒�P޾{@�Jq4vY�8fW��j'�˪E��;x]���^?+���U��)�f@���Hd�7�(wٝ��3��������1��ˤ����CN�〔�km��,RW�� ���k 8�,�vd�:��r�W�4�#����W��)�$���� �F�ڏa�)p3�8V�6�x�-	p<��`F6���#ֲ�&��r�0rk¹���|�Q
�M��G?��,V�����V������hÅ���L�^,P�`��[���e�*`��L�Yeq��ꐕ\Yl=�[�7�Z>���d��]�]�v��+��9W����dfj��Ά�����+^�m���zhOm����%�o���{Q�����E�{}��a��yJƮ\�?4�`�l��U W�k*48�V:��M\������������_�2�.e���M	́X�n[�n׻+����<C�nF1S p;������O}�zqx���	�/��~����ç7a�+ઑ��6 d�]�0���!ex� �Js������n���3���dO����I��v��4���/����{��<���O�����!B�[	G?��G�9Q�O���[���7Ŕ/I��Z�f�J@ #Q[��Py�bD��۴�
bY0d��.g]��׻��-�}���[�����rO�5{�G��q�r�p��Aal��M�T�N�e2!�Jr$�IL�z�0�����9TZ�,��d�3��V�(�W!������cG��1c�q��{di�3����{޻ל�ptO�i���,t]9�Z �|נ͌T()��{�}?�Q�v���[}��GB���u��~n��̬ܽ^2�o�T;��%ru�a���e��5I���ܱ�h5*B�f�ٟ��ȇ82��Onwɓ�1e�t�\T�)�j���N(as{k�ȫ�p�}�O��g��_��p>�����0$V����0��j!{�X�l������ѵ4��l�Ȳ4���D���HS~��|��oڴ%�OβOg!O�M��F�w�$ߟ+.���H6���c���W�PɞCc�CcD�����������O6�8���LW�[��^��Rh%>|��|�Mn��6�����,�Iȭ�a�V*2�t��j�$����vd��^�Ql��h���]K'�ڣ�G�l����YU�����{n��[��p:d��*^Zh�����ߞ�����Kn�����S�~�l,�m�9�P6���L�?�ϦәD�o �d*ہ}��Ki�x/dQ(\��>K����DT�D��C�x'�5������}L�j?I����?�]� ��A�g�9��w�����Hd��2�Ԡ���2˲L�m��ݽ�����y>��!����!����r6�������N����	�x�)�H8�p�e괏2{���� h��Ƒ������0 'FJ�4R!�ܭ�w�a|(f�"^$�0K� [)�R���R%�#�L�b�p�"Q�׋���K/?p���y-��R�o+�����m�bZ~ @rT�����@�8;3I���x��`/��s�ɿ�]V�)�*]�4Ft����,&�b/C�{��Z+=��7Z�֑𣯅��s5�|������Y�^��D� �w�=�<�����n���8J��TB�_3Ҙ�nxS@�K�A� U[ Mf�H��	1)�,�P���c��M���W��F�E�P��H�e��oFs�[i�9�U�ՅLˑGV4i��r%���#�6�tM���/�f
f��4ڀ@i���_�Ѽ-�YZ��(�#d{��B`��d7�S��b��j�{��H�á|-�/FZ��rz��=�E�;���ߊ�p�Tur���HlAm).����;�q�y���>��F(�� d�<�nE�NK�Fk
=��'Xko���,e*r�Z�m��"����Je�w�����nm�x��{��L��4�&a��ΑQ�k+�_ @���,���r��3�	>�X��pC�Z�uWX~U���إ���W��A���,��a@��S�w~�\��q+=�������:!Ϋ�$b�Bmۻm�����@���8�>��SO��ng�(y�8\#�o�7g��T���WX��l�}Ζ��_&��kJ�1P�\�����F\��:(d�%�sM����kxBzG��������S����y3s��~���(�z�P3�5��o�Σ�o��������}�5�(p�+c�o bq�<HN��T��z	��e+FK�֣c3߆��θ����'�u�R�f*E�*ذs��fH"T��д�sK���V��9Zs�\]�^IB�K���~���Хh4����6���y-�N��A�G��h�7BT@�y��M�����4���AџV�Tŉж�ӛ�Q�Q��k�k͌���1��Z��w�(���W��AM��y���8V3 z���1G[�f�DqW� �y���M��g��k-������F/4g!�Z�q>}R���k��M��Wࠨ5]�-ͷ��w�D��0���.ӡL�Vg�B���n3���7۾�d�h�G�zW_�]�-i����/� ����\�e�bD& �MY�H٫&�F��^�c4�{�5�J���
H����JX�q�$�XL�F�ăhlIh�ꭽ���h�w�c�|�F����E1�n�W�IVI���r�<�����Չ�kz�g���V7�/
�5�*�qU�>��,!Q�����^���Œ1�����`��Z(�V�1�b/AW®tp=W�������P�7���W��v�,�n`�����u,Z�)�j:Q- �����t*�z�y�no=Y���V��B�668J�J�{�@�������yrŷ�w_��8�y�°o�V:��;��ß�8<���Æ7OR�}a�"%G���)��_*��AUT����#���$
}o�uq��+U`��{�@]7\N�8�1� _$��"����OϿ���6%p�xG���A=w��}-/��a��}���[�>�n�I����c������tx���4*Am��K)����t�7�����P��I�?׭"R΁�`v��׬���鑴2���/��EDs��R�ոEF�.&#9l��\i?��2f��1�k[�>l|�w3�o(�+����uޤ�d�&>��P�e���I��+ݨ�2��~p-��Y�]�n��+�5"�bZS���^6���Bm�*��Z	Z��U%�k�r׵_k�:�=��=�C��T����f;_|��xӉ��q�v���ȃc#;�	�(1XP�6x
q����T����T4��4X3n倗��tq��p٠�0<'0(g)oF���07Q_,�.=�U�s��}�Q
�	��t%�Y�s�*W#FP`䏴ՙS�42=V���-{~ɴ8�k����B�iRVz��z�[Eb�A��A���:���=̽	Pv���#�|��F�4b%��m��Z']�_K\�y�`D{|h�?�(�A�p�¾����J(����U�וe�hZ��nĳrsIo�7ls�ڂo�0�$��)�ڐz�E=�����WBYmA7�]�YRH��R^��C	��
p0�FEF���]`}������k��[j9��W��(󤫛�}��ckxK.z:��:�����@�z�Y�c+����sP���?�~�F��oP�{�wO>CD�<@:��#/��e�Ǵ>{^�u��A�H�R� �����0� o) ���,�FF>��:���0�K���5�}�.���s熟��-j��&m
��G �|����<|�;?޿���H�Ǭ~�����=�������䖆{���w�O;^|��A�+x���kdJ77mH���?=&<�m[��Iى�fl���&c�1��1�N���"�+ox����ɡkTVT`TL9�1�;���?;�ri5�ˋ����ֻ �_���3�o��ǳY�q'� $/ꞱQ�� Qj�uv�F� Mq����*5�5sՌq��c�� ��"���hSކB�Zc\b��y�M�3�Fo�(��騇������
�P]Ft�A��!:�Nb@��0���Q����+�����;�-�v�n��D&�b���c��x�7C|A�8&_�+�w��Cw-��߰�ְ�>�Da�k��_����4P_Uy����پ�+B�oZ�����^���Li��Lo�����,)Q���5b�'"7��E�卶r��br�_^_�����`.�!�S��9"Fc7���q�xЩ[̚:+���~��>��Z�B(��p�{`���b�]�eQ�ps����7�0OSB����S�mPJ�0su�*v-�n~�o�^NS sh"V�����r���{�̬��u��� X��skzkB�E.?`x���t+h�ս�
�l6�OE_���"�"�ۜ& -B�Q�[�Hoī=��Y��}��n�(y��7m�3����xi[���<���e����O�1?�Gw3�����Z�|h����.���Ru��H���X ?���K#�5!9м{{A�O�5�U��_���8����u�S���L8X�vmx���C�������ej�	0�a���?����6P�/Ѧu�?.�6���\�"s�l�P���Њ�6C}���č�6�g	�������3���-��F.HJ�m���0��1�.F�9H6�$�qb�R�i%�rM�#��՚�
&�chi^>��'�o|����֤o�y���i>��/�)8;�ɀ��P*x���۸k�(@r����ֱ�6m�B�:NK�-�=�qK"T
�x�}�y�zkͰ� r�}��>|�{�#K� �H�댏�.�{J�����Z7��
�%OAH��7��4�Ka��]�F��89^�	�3u ��7;��*�����t�6c��~�Ţ��;*_L�I�k?t+;D�+�4		Us���m0�h)m��&�`�J�d>8����������jAJE�`i�(j�O�)�N"�H���QĒ��{�7I�#(8�)�fd�as��%��TZ�����d&z�r�#������NOɵ:w��|2�Ӹ�Us��>�{����WW{��O��L�И�p�g"7ȡ��|Y�|�?�(�����w�^"jջ�/緹��[ُu5����ݤW4�PS�<�G4k:�Cڦ�=�Z�������
ǜ3j����\�.μ��)�%�)��P��(a��H7k�r��ꑚ;�L��c4De�ɱ)��y6E��|�k6�(�M�ӕ�L�	*��5�?��φ�|���w�X�tk�p+�q�\�o�{.�BnY�eYS�WDK�D������M �I�Ys=A�BW_+p� Ebz]9�-�f���Ǜ�J������Gh��5J�"��-j�W(��K�O~��c�.��[�(6����O=>��Ɖ�,�>�����̟��O鋾}x�����)5���Jr�Ǉ�jr� t��Y�7����	P��'{;�B��Ĺ���>�ܳe�����C�+��0�<vt8~��a���^hi�E�zvM��0L�p����*ty-�ZE*�Z����a��-D6q����箜N�x{�|��a0�-���D��wu��ؽ�S�ڷ��),q:Hv`c��Xi܆11{U�^(n��
/ 0=��ᦜ�k�M'O�L8W�R?}�T�M���|����Qڮ�"g�x���?�I¿<� ��s���pp�sϽ�0�QR�wD�믿��nݺ5���h�����p׍�k�-�U^�7kY3�{DN�g����O^���T��Y'��������"�Y�� �hr!	�+7�\���HY�8?��ui,�=����x�T�Ƅ�[E��v[��M
%
���,�&�j�c���\����Z�m��d��;!��u�[sN�������v��s=�o���r9�F����>����Ez�;f��I��m���3��Q
���|�H���,�&��̳��k륈*�X��QE�A���&˛��訁�5�o�x,�ֳǩ�#[Z����@��D��l)甴�+�yچݕw��&�=J�" �P��®m�{�N�مO�x����:
$Ta6�iE<ե���+KL����
�1��S'aJ{B��@����!��ߦVy�ҩ�F���ѐ�������oa��ڼ�w<��m�D��eYz���+�tF�ڔ��x�.02R��x�O�����&�G��Y����EǾx��o���J6��Ǐ'�y;���ԑ�0����dmMM6".�;��WQ
;BV��<>|鳟`�@��]B��޻cx�8�;ߝ���mU7��^�u�R����������D�.s=�9���Y�k����3?�i���=�P�׸S�����u=/��Y�H#fC�����g�n�Y_}��ч�J�s�>.�՞=}�����X�>��0	(K�ۀ CzR	��^	Zy�6�֡����8�d���]�az3�t�Wٛz�-�j��������E'q�w_�;��RN�V�c��2��u�.�s�N��e<�t��[W�
���n��C䣑,�׈R�������th$��)�s��w����5Ǣ����n�d�k�l@�[����u/�YN�c���4~3d�|�HP�5.sa�,ƹ8�>k]<	 ��q)��7O���NP`�]=ٙ��ФB�M;.Q_,1��;�b.|�9?A���E�u׉�ۗ�"or+_-�#"
����7�y���m5�E�y�R�	�s}�ō:Ǣ7���������)�ߌ������b�{u�yO���f[�G�G�"-�̄�*�R�]��?����-�PqLJ�E����b�sk�6�w�m�,��!G��hf@��E�x��He����;�vi�֕z��=G��5�ۯ�[�]��r�CzG���a{ CQ%ږ��Q��Lo�7���K����X�1�l3��%0v	$���[ J9t�p��֣L�ʑ���OT@a��nº��Z�56�w6�f��κ	n�v���@�V��!�P��[rd�:щ2F�'ᮢ������w߻��Z��G��v#H�3����G�G!��Ƌ�H��g��0Ϟ� �qc(�O|�I��_�X>9���?�yܲ}3����ȁ�a��㞓���4�x�����&�������{�� ~/�~�\�|��utػ�� �u\�E:D]&Up2i4���WV���R���\��7�.�����v@ͻ�Qy�'1�0��>gc!C�*o@�!�HJ�K���>�������d
L�������7m��22�,
}�*VE �U��M	(ح��*^��h�}MaV�qC�O<N��S�վ\�ߋ�+u�`|��ƙ���>�����;�9k������a������~�ϩ�ϝ;/^%�7B��o�K�����k�Nq�`bTX#Fzɯ
�&K:um셖W~X+}�y�?¸��`r�(�h=�uܖz�*6Z��rH4,��hY��)��')#[G�xU��O(����4�m�j�lU�d�w@/����xOw��b����u�8e#�F<����\~�Y��^��R�e�{���:_��r\?�f�7���@7�˾�~P���b�5���<��&�1E�%F�-Ѣy҇F��N~~�(t��A�����C�`o�23�_)��������-?�-�t:`�OdϗE6�A�BUڝ9�+��~o7���X�t����[�\�fh��.��j�����G<u�Ӆ[`Q����Y�e�S롗�\��uޢ���cu���R��R3�M��X�����*����ϧ����3�����n�ӛPN*_r�7�H'�/me��3wo�ܚQ���ث"���|<����]E*T�=ק������X�Ȉ�9k�y���G?�E��c�ޖ������5��o|�f-W��	?h���O<pװ�<�>j�=������H�����?HJ`#B�����	Ť�FB̀t4��[]�rz�z��p���BV�-_���	�TLw�&�?	�����j�f1n��矘Vi ��^�0!Wю	<�� �륺E`	��)��P�\���(����]����"`@�W`�KȚs^����>7��?�ï�G�,v�����l
������k�,4�[�(�+b#%l�W��j9ZX!N�x��jM�h��o��/�˽���z<�*����D>����Hw��um�u�}���������<J��~뷆�{��5���=�\�̿�G�1u�Y;eT9^�D7N>�[h�Q�牆Q��׈�l"Jt��=7���`+��HMzz�&%ʙ�����^ެ�짢�6���\��S>_sQ?��R������
sת)'c$"�h�^�~�sJ�Ǹ���_���Q�5e��i9������`oND��k=W��{.>��J���%�<��C:��l�Į���Y��O#���1��"w�BG�����K��e�,�n�L�h�Η����N9�A����hH��7y�7�z<�B����⡶ܕ�7���zۅ�A@?_)��L��(�����{��|�Ub���J�F[s�6�\�޽{�ε��9(�N�2�GE�G�ExՄ�IU�Q����O�a�!�^��׭ �Q"�c4���h�U[�҈}�r��hQ��]�|Kr���n��j��X���P(�Z�ʖ�©zo��?IL�f3���ն��ݸe����?�~��p��{���vv�P��Aj���u�	�k�b��رe��8m��:���Ƭ�׳J>Snup�[�D`vflطs˰o�f������O%�`��+���a��)��
�NB�I�����@t@�#�m�r0�bL_d� B=|�
�4�m\�ᚖ���5ap�5||��}ۇ9ش�	�?��/�0�{�]�wP���p����UfZ�Mo�l��1�!����o�*8�C�Ғ��ٸ=�n���es�0r��b��5o2
Y��t�o��o���
炈�n�t�rޖ͙G7'���`���o��o�*ٵ���?�����?�T�a~=��Q0:0���[��%T�;����[��U �*���v(c:���%�l��:t0-|Oѫ�ƕ����$�U��dHV�.���&{]㹸�E��{"�R�떉h�����1�k��g\h�)�M��7W���9+�E�O��<R�˿Tx�^_�)c�>��wߥ��,�Q��-]�ܑ�^@l�܂����¹T�K�Vi��{�E��ږ��MD�<�x���8r�k�q'>�c:��Bbw��)������n�(,חs3��Qd���@�6!��(�f�^���	�7?� 5��\�:���u�fH�FF7��*�\�n�[��d� l�Xs�������������C�>	���m�;�+�*���Ϝ�w�guғ�vh�T
���~���'A�ޤ�ZZ��Dy߲Fk�l�[xL�+�&���8����ǌ���� ��:V(��,���Av^��f��{�}��-�#J��-��*��E���ί�Xfvf?Cx{nx��w��(�x��C4��v� �
����1_�{�-+�w��&*s�#`��K���]��jt��� �e
C��m�Ƕ��nڻ~�Ệ};T���/P����7��4���)_�F���(X��߂���D1�W���q|�!bDJ�_&��2O�h�Gț������͖?��<�;��&"�v;�A�s�P�����l���l���VCv��102�����4
�̈��s_ۣ�tv6�{�n�s��\� @��5�mKW���p(%��8M�َk�4��w�}�N���[���{�{«�?
�Ν;#+zw8C�K���.�F�Y��?���i,}0��(^ߟ=��>
(�s�1�F�~��50T����A������ʐ���"/·�S��(c���Y��g��M��ɦu�T�>�3�7���,�ri^w*���_��x�m�� *bX��jV5Wt_�۔��ټ�;4����=(��d<�eqe�z]��G�s��_E���˟�RZ�c��M��P��j�@��k���+�j<��C����Z�����(�UWmu�nҮ�no
��z�j�`S�0����o�Q��?������=?߅A���[�Џ;*$Fa?F7t��)4քb	I��
�E��+]"�4���l�?�Nݻc�p�&%�+�l����T��p��p���6Qص}�p� yG6�['N��C#�'�v��ݥid�5�= �>K�Q;��Ү�iK���3�"n�f��m⡇ڻ���Y�	��Q,�9E���H
�����?����fw�!�p}8rx�p�й�����I�[��u<C��i��ѷ	S_B�V7�!���Z�	[5� �	�z߈
��K�9�V�o-O�s`����y�Y�֍�$>S(���w�������h�s�:Áh�ٍJ�gO=;����*�-n���]KNr{~8�o�h�V)����R���hN�q;Ƚ�o��<h#�P^�B5C[�M ����nb45�Ԓ�7H��A�T��9�Q���}�����]�T�ɏ�Z��5:�#���jѺ����U�7h���p��)�	|=��6�ƹ��5Q�ʖ.�R��?y������G��tע�9j�e�uv��0j�����Q��R�DalK@��t������������.>�{�	�d�e��l���c�(?J;K��Yq�s ^���2�Q���V�S��R§-1*ڢ-����P��{��Q���ɾ̚)o=�ʳ22Jn�����7�F>;5yss�`}֑4NZ$4��KK��~�:��FD����M5�e�o��T	P�:��:���Awd��Nnl�P[J�>(����f��bM�M�׶�*���2эW�j�u�}5��2J�t��c�V3 |>z]=?���2����qG��hnԋ��O������W���%D���
�`������,ex��������J���ײ�������˿���w~���� l2=��~{��o=�]���KU8��Q��Vm��Sl"Ѹ�2���u�g��R�+�2�e�!lJ$�$}Y�e�7��&2j]��O�y��̰�u�R�g^<6������ �]'�2���a���U�<l#��H�۳-�����7#`,����\C��S�fl���5���MYP�w�OOu���Mݲ�ĺ�nnӖ���
���;��T��47L��4|����7�7�^�N?:��ҋ��I`��q�,:���j�eв���MflU�����O~�>��)�C�.���#�:Rh�_>���s����Q��_��Gk/vƶ5�u��{4rE��NCjd(մA�����d4�N�@�����U������|���'w�a�
�P{7��LH9*�ei��h��}ͰY��O9��%� jE�a�8���=4$� S��S�yLgC޳\O<O��k}���>c?a�1*T���S�ҫ=��R��3|:֞K�����q�K�b��V$A���K��h��8$�d�ƃ����g���Ջ�,2^��@DO��i
��Ƚ��R��d���ߺ��z��0Y��qݻ/m���w��_���;��W)��_����C���L�R�n�[�]Q�z��F��׭ U���J_�i7\�!�������������z��������]P�U!�l��F=�n��ޛ�x�_�����֊h�f����7���~�f&o�?�c�y-�pѐ-�mt�?�����������~틠�g��{�G�Y��K��rnzۅl����zЅ���0�n�Ox�����"5TQ؊��n	�dZ[}V��۱j�Z���;Ǉ�����S�%�?��q������B/G�F�eI�U��%� ��s~��ru���DX�&�]�(��0Sy�#��m��=ÉS硚}���	�n�p��$��Mx�� eYi]���ؘ����ר�>2|ꓟv��7��޻��edx-���]x�@�Mn�h��ER"0��ّm��i<�bP�%|�s��\�
�����Djv��5|�����/��] �9�� �u�q�GgyT�}�;U�s{29��k�㬳.���`8�!�3\Iʱn5jԍ����L�ݣG�����T�e�B[�6���~�%�Ͼ՛cz�/[�4O�����p��<��0���v�}o�W4|������0o�1�u�U�ݵl��q��y܃g��Z�Y������:|	x��c���V�o��&T��S�T��Ζ�aٮ�ͫ0�t��7��=g՘e~,]c���2p�|��j��viʚ�&8���2��`+�:��o8�(\��/�<ɽQ����i;;��v�Yw��W�{*X�`�}1@[YH�K�z�,�K���[E�D6�aKl/�7�Ք��z�j��D��|���FI�T.#�&'�n2oW�����
<�+}�����66��h����G�ص!��e�<i�[ϑu��n���\{x������u�н�Qo9ۢy>�!����u�r4��?߿�?3������y,�;���>:< %�|��ָ��7!��I��Y��4�_��}cQ+�(�ϧ��A��A������g��9rǗL�aL37E�^gдQ��Jd�t��x[n{�h�Bj��#X�Ӷ��筀!�܎������/\{�rϗ�^@#��]���G}����3x��gO��6d=9��1�vQ��q�x* .]�Fkǭ4����>���G���0 �zr���_��_�{�[���l��ȯ�n}�|������5v���/V.#�P�x��	��^v/�)*�)��~�4��8�,\ ��ֽ���wx�����Fʤ7�x	e!�(z5�Rd"�-{��-����������`�_g�N�-0��ݲ�~LĲ���!�[�W��<�����YC�b2�77��R��&J$X�2���Ͼg�am:]7���={�D�-A'|��6JU�7��{s�/��O~�c<����U����Z�����h�L���{��dS�9��FJ�D�[�nOo�/�6��r*[\g(m���c�ZY���!�j!�!S�1�A �Mz!\��L4a� ����.���>֣t�`���q��8�[�}�S�(�µ�b�����W���0�;%�ڸ�fƎ%о��{>y���{��'�
�b��$B#Xͮj��=�W�N��p2��T�{D'}��g�y^)��}L�J0j�Q�u�C�lE�-n�*��s�Z(�K#V`�b�/I��O�$`\��K81���nxY����e���W�%�u}G(tۦ�����)i(�`X�G�3d���p��mH�q#�k�)��q-��J��(b�U�������!�
�U\�{��~��*Pםm�wME�4�+��Χ�{�l4"0���itO��u�~?�u�
y�g��� �����4j��};�6kmA_o$7ڕg��k1�/�?��	�mg�Y�0�-<�}j|K�Wc�r��k�f-��u衏�ٞ��Q-�^��R.����̡�b�\}B+k�}��gs'���_p�J~Ae�W�P��Ye4~�^J����C�!���}N�7���� l*���ܗ�����-�6�x�
����ϜZ�z�9x�Y��?��? Ran�B�Ρ��x������K/��f	O��h�������3燧�r��q�|v�ҳI�#Nuy��I;�N�7}��(=t�$����~�l����r� �T��������0�M&�z��^"Mq�:w��BC�Ϟk7H����W]ʲB1T���	o��.���7��K/z~~nx���
{۶�	���1�~5��~����)s٘��U�~�*ts�c�4��E�\�.�B_�1�s������J���eª��F�Ч�;ʯ[�GTN����P�>������˯�!��ڸ��&���	/���L�A�u�^5�S�1S"��+G��[�i�Ҕ��<v6I�t��������c�����Ki�깍�X��PІ���(t�m�l�����95�7p�(e��C0C�IbR�s�wf�C����vu�u&#�^�F��Zf�<��g�o९g�\.3f�Sx�IePwʫ��
�
<�����9~���ϟߨ��W)�:�5�����ە�h.�a}�?�P�h���g�
�!��P>k;��Yx�y�	�y"�JД ����Q�|�����Vs~�/��[YJ�H4zz�$��$f1̥�+�3��Ր���n����.��n۾u�qe���Lʦ�)�m�"�6�%��%��"�eU�G��_�R�.4�35�\�p3筷" ���3�
���}��/������o�XZێ}��׋�d�#�!
>���.<�i`�1�۟ky�8�xN�t��7��<��ؐǈx��L�2�L�����U�����+�Ϝ{�p�L�4�
${���\�vO�R�#=����÷����ЃSQd��W�-�ҵE�f��\�K 	�- )>���&A-"#�8��+ MF��\��@�� fn��	x���o�8;��{�~�Y�^ZAK�ת�|�y�-��x�`=e\���Py�Z�G�X"(F��[��]�"���{4*�\��[�p�H�ji�� �����0���zr����o{I"���/�"�z��1 F���{�ˈ9���fa�#���:���>j�/�e^r��ި��� S�f]C��a_u����7��ؓT�\�L�����:�'��� �Z�U΁�[G�r��|U Ďu�TY+�3U��s����cgiժw��hߖS�G҂��F?���-Nf�m`G�Kl���<N�b�A��9��t׺ڻ�tuH�0<�o��P��x6*bT�e��F@����i~��կ�Ɨ�O��S`}ڍ��w�9� Cy4¨H�6.cD�n�4RH4��'Bb�"�X�������kyF]������:g�'���M-� "W��kn�
�S��H��g�w䆫�N)뎦�������9�������tEdv)�B��
ܩE�r)~�gz�����[5� �'B�m��=7���ٗ�W���|��# �����h���$U�;���c��8�Y�Gp�q?�!j�F��"F�X��n����-� ��Ƚ%�g�K��X	���E���6kg����S�4%�ؑG^���N/�OaE�M�VC�K��ϡlqu�Z!��,
\����4�Y���5�w�|���뷇̈́z�Onx ��ÃG?��χ��.��we��{_��'���C����e^�c�Bs��q��<�Y�C��Q%f8���&Ü+�k��p���$��s�
��̪���5�m����Fhĺ����FV��S��UE&�󺥝���Z�Q�%�/Ɣ���\r���4���6"J{U���1b�=��=�M[*Iic�y�2�z�E�\���ź��H?��b>�A��^�ىiV�U�K�m8����#G���q���s�o�k��~�����);���� ���AJwV`�MZ����1p?��G�@gv#@8A_l������@E��-�@�#b�ޔ�:+ݬ�D۲t�����{8���$R���/%��������n8�u:+J�s�Ȝ���r�*��0 p2�eK_�A�ԛ�"��DO\���s���%�$g2u���Έ�ն8�~��ᕗ^.\<Gl��я�����9�{y��+�n!@f>eD,?�#��A��PC����x�:��>�;Fi�y�,��iQx�uZ+)�BGi���&,�x�=��Ӈ�o����[�a����5�[m�(�4�(��[��t/�pV	ʘ~��F" �e�5���g~�_�j��ЮA���m�K�ݕ7%p��z_��X��{/Jo'!M�va�i�B���h��W��f�d���
�*�� �s�P�5끱�R>R@!ˢ�VƉ�R��z���������1>ڕ��X�e�!AS���>�я �"׆!���/j#���u�� ��x���ُ>B,<�y��:Ы[��	ᎍBlbry8t׮᭷^O>w�P�ۇ�ss���9̢h�y���"�˒�,"X��?@�pWB��6�nϽ���U_{�V���r꺩B�u�R��88o奲��b�s�r5*`O���4� ���jc�w�][�s�<���Lx梢XkzA漛Kx^(��2iq*𫕒i����(�n
��"�[��*�[��]!�G��M[�q\]�=�$��6ڞHڠ�ٟ�Ǽ�N �T9�� _Ŝ8$����a��k1*/{$��w��.��[5�c,U4n��&��c���Ű9���b���H�l�Yˆ�3�w��1�sx���a����ṗ_.B�,�KQQ����h�u���������2����pP�e��[���#��]�"E,
r�����3��.^=���f�y�sMkh] �r	�}9�O�:�{�N4`�u`EMR��e���s	�s��ft�"N�k�6���d��w��sx�q����k��Q���X C�n���އy�%�o9�Ir+����" J�s�$���#��#��s6֮��>��? ț ��Qm�+�nߊ����mu�eE�T�������2�f'kg���s�)��ZM�T{�s=�f����f��hRX9���w�C/�G�lZ]l_���`�z��)���]��N�"̇Ww��S�}�P��m8�Ojbϱ)i\!��_i��uz$��m�w�Ǻ�j_� ��|Z���Sc�T��<�֌"�o�aT`¹*C,�临s�2T�;9~�A�y��(���T��76�g�n����<;<	����=4D�~d?�����˶m;#��1_����������7�7���ςt�}��hn��j��n�lټ�\9�0xЏ?~������6�˞@���`��W�ܕ2�J�Nzz']�ҧ�J,�r��kߑq��Z�QGO $�)�Є⽄���4ү<���j�-�g��|`��S�	��.n�ǐmt=KD����mD2����������2�cIQz4�\�%��'/\Q��T?O��O��ؕc�p���MŰm��TYx�}Ҵ�����/�@�6�`�Ɯ�4�*c1'��� �^P�*}���R|�׹�{w����~ޭ��HKk�RX������z�}��5xMFcV?��3�e�]!�}��9s������!R7FgX��bd�}����P����#=�Q�PK�V�T帷���I�"j�G���������0�)��m�bӤ�Rk������笖G�B�e1��+�רܸ|�"J�<ǆ����({@��V�H*�5���U�P,eX j��Y���,��")�i�?�#�����"7xq+�RX6:�����Snq?D��%��kb�Zl��N�uG(�3g�<�BO���+�����z�iS��6⡛�r+&�Y��*�X��+���9�icu!��fߕ�6��c���s���Lj#զ�{���;�4��{�B�!�<��z��Mx�?J3���B���`���Xʆ�@�^Z��� ��g7lb���>	��1Pۻ��n�]-����t�76�̆1:�m�x�}V�8%<����j��eNeP��7� ��5�F7�F��品)��Q݋��Nݓ�ס@�GP?���^Ν;3�w�����'N�&���]Ò�I�Ɵ}����[��O�n���$�~�zB����p��"����'��>|/��pE�;}�8��ΟG��$��j��'������������"�ERQZ��Ly��1�w*ʤ'cX���
zh�y^��}��s2��642.
�r������n��H�R�Q�#�L  ׬�_On}3�Ķm;�Ӕ�A�*P�9ī#^ߖWh���:sN���(`�����|��.i��uDy!�ס�r�
��`���a��O�� ���} �>ɹn���3�=֌Q�������W^ɱ��և�MYT�2��L�YI���=��B�Y��+�h�NX-Ӎ��ze���.v�,��9���,l-w������NA&$���mɟ�h*��>����6��������SI�ŕ�
['"�ܽS2$��Wբ2Ճ�ܠ7�R��:a�ײ4s~�,�n��>�T��l��c��2�������w�?���`"(�q��u��
Q�MD��Ll�>���?}���J"u��@���J�	4���A�,�X��LDjy��Z|�9� ;��&;R7��R�"���
�f,��_�˻��|U��M�W��G|���"��;Z�Z�Z��_�Th���Clk��&t�'\@���� "@ݿ�6��iJJ�VK�l9MYp�������[��ZN��H�.��������^}�J	��sӊp�w��Ʊ�o_%4��{�j|���sj8v�,�׭��]0�ɾ�&�j-��]z`�|�:���p��C!����r���gtUEZ!��t@�E!��ߚ�^5�F���Uom��ֆ��`UI2V�Q΄w��a�޻�m�ۆ?����e��D��$>t� ���{|����\,��#�5���mG�T�voR�2S9**s�zW��%���T�m���9"�����3���֕F��X��EB��[��x�έ�h/�r.}�υ�Ӛer�1gT���w�x�25N��c���i�#+[^���3ˏT 7m8�o�q�hog=�{�ܮ�q7�*���LM�[e�rDs�^\v���Q���C��*�E��8[ޫƶ�c�N�I��(�E�]o[e�O��=�r(t{֠;F}�o9�=��g?[�|�zT�6e�����!�M��j��e^�zu��!2���Ip�U��~�a���I�b��2I�<��"(|���x�W�ȉ�B����4�=},J�,�5���ƧX�V���$� ��S�Q�� �Z��i��0R!�q����
���-��#wz*����T���62�<�D5cD�1;IYޖ����w�� w�p���ͷ���b����ڹ;�����4.+��!geEpB�Ş���T2��NX�Ls�� �R����H9.r���k���<P�S�3ރ Ks��J@�EZ�s�W���\�!�p�v�U�����T��S��p�:�E)X��	���������?�R�ցy�]q��v/~.LX-�չ��ZW1'�Y�OO�ŞZ���.G=��Ʃ�o�p�I-ߚGIlH�j�Q�P�r�����OH��
���m�=KxT�Q$2�ݦ��p���]�B��j�8B�{HZ��RA/}\����\�%4���!�Ǫ��{+߷�ښѓ�ݷ�9Of�a��C�G��|�r������e��SAn_��֕݋x	�	��MO�p߹D'�˷��4O�>B������w�'�Ͻ'���V���5t�|T
ȉ25�D)oU��"ԩ5|e�c�f�_�����.�w�����w�Ee 9jR�_�.zzZ�=�6󻛶�2�۶��Hv�|�k7�����w���
k#T�՛ẁ�Q1w�������?�P���u �RV�[���M�Q�_�җ��=?����~Ơ�4�/�9����>|�p�ǽ����tf;x�`�D�خ�͛[�.�1<�q�FdMS��=�X**rRh}��B�:�A�Q�������	�)�8K>)�Ҡ�-�-�#�|�=*Q�'Ξ��Q� Ϊ¡yԆ֙v#oF�R�b/��G�?E��<)�E��b�~���ĳ s�DU�H�sF2�m�3��2zȻ��dcM{)���~���(w90h^�yv���C�'N�����~�I6��(H�(�m�Ml�_
�N����)���%ݓh�t�|���d6��	@��k�~Y�Ub�s���{�֠�����]X����M��4d��js����J���>���-g���u^�|���Ek{�cv
��q6���Z���%\`Z˱��܅�����GN�*�	���b���Q�w�y+��'��cTN�SNzIn��`�?/�{7��� �*�����ق�ۏ�|=J`7V��,K����+g�#�n��y��"��*��P�lS�b��5���ꡊM���/��z8׹�z�l�h�.+x��H�iSr�0=z���g?�	�k�W��5�x��g�W�=?� t�G��ko�z��p���{�`k����t�b����x�g�_z�<��tM�Rr4C�6y�n�jX�s���6�R��������E}Ҕz�K�oW��QЈM;��s�Ʃ�1k�v�X��2���:��N�J	�]�S.��u>���}���Í �(9�[O�\�PS �����Q�=e��K��<���<W�T���1 O�	B�c�NA �kV��P��+�����%j���y�Uu�4?A��iM��H�ֽ˦<��?��ᩧ��5\�ç>���պA�z!���hL�^^�u�΅����a����^KeI�,�3�l�����N���9�V��S��%4Gj̞ ���l.�����������s��"SOz���sou�խ�4~���';����3,ş�531��͉�S!�l{?�:�G����4JR'Kz�Bn%�������)Р���|2\�0g��L�X�
嬍Y:�>���wh��j�@�9
ގ�\�ԯ�������3_���Q���L�y�kJv��tp�K���7��%]����Q����2����1�k�rh=̷F@SԅO�jJ��(j�`?�r��s�uW�w��\q]W�C���̾���&�^��l��ּ�|�+Jx��a�u*�q�P��7<{�w��ل��|d����?�DاކDe^�V��%������/㼜<���l��cg����.�R�J�"�f����@�������.��rk��5���RM(s#@:��gl&�2?�2�ַ~2��HD��������>w�(E�ɻ����S�����a�7�z�?x�p`��E9\%���5�	#����s����mÏir�}a~p(tǡ�=z��p�<@'�����H�2�����DzJ�V����?uo}���+�[�~M��sX��G)FaS6��1�Z2�Ud#�'���[�����Uۇ	������a<���!��#��5��ZR��/���`ޗ�(u����hz���l�F�D��D9��Vqv,L�Q��7����}��P��ӷ��}�N�{=�֍��Y��Z7J���~4�ѽ��.���2�O/k���p���|yf3�݁~�z[N�oi��@b(��jD�d2dD2�m���G0'gUWA���V��-E�<Y���JmY9!�����U�1J1�E�}e�16*���f �����LJ���X�_|��U�֣�+��\UfDC�� M]W��?�U2�j�Ү��q�05YkVT�ڒ��r�D)��"2�1q̲8�kʥ�C
����%���1" �_~u�:s�{k���4���Rv���x{�΍����B1��{μ�����Bq5�ߔa?��@��m�c���7a�l�2`�r�.�)��'�7?eN� ��eyf�g����-Q[���e\ʡ{�i��Z�Bp�!@��\si���;Gy�g���������3}���w�����?����g�C�JJr3�M�lm�I)'�����o��mO�|�������αТ����FěWQGn� ^ۘ%l�l¯{D}�z�aU�	����|;f̬��lt��E>���ڸ�p��~�0A[��k7�M��ax 2Y|��q�����;H�ov�����(��D*���P�|�^��%�!������a�{�O�3��#��y�ҕ��#`�� ������M���C��t*]�z�5�N)�R�k���|�s�:C�d�B�ѕj���gZ�b�lhpp�S �'	�&="�&�=�z�!;�ځO��2(rrג
͐�zz����i5)3��l���Rr�%��='ajäajc�̑�z�5C��My�֋w������W� ��a��n��+��݇rè]�&-`w<��xe����R-"�>K�u}�G����&L�x~��Mi�B	I����Y�&�{ɩpP�7q.I9��Xq2����3i����8��FA��|��� ʕ����6\�Y�ab�=�r�4�̌M�4o���Zn�Βk����S��=���P��X���
4Jf ����Mos�+�{����>M����|hЅ�^
�nql��`��0�}�m�tם�l�,��$ę���'�vX]���o�B��c`�MZ��������/S�<�R����J�B�6r卺�ݰNg��G��g���͔������&A7á�[9�`�����л���aʛ�`p3&Z���T_{��J�Ɖ�w�6M/�®�:W'�螺���Z
���w�4c��P����_�����������=>|�?�\dr؎�����j	��畅��̮�����aw�:�����Q
��Q�S�Ү=����5OsT��6��hj�CeT�y��U,�\=�Z+FSd�ByM"<�Pq��e�wx��O�tt�D�r�z�1�x��i��w���"B�'?{a�v�2�y�>x�o���#�w����e��+����|�QhUOsN���<��ZO��}D�����T_Ö%�Ǩ�^स-YJ՛y�<b�A__�%��fx緓"���K-��#���	�p��В���Si�{^��4+��y�*k�G��ʡ���1��쑶=���(��U�A�Ⱦ���s��#�9Rk��!�,���wc�˓��F���B�G�=�vT��T������'(���xW��37�!;�C���b�B��?�1�/~k��_���p�VV�+��m�R��:�*W/��]阤ɍ��5�������FZ#@2�+�A�e8�H78��
Y��5ra���o���Qn��D�lq�8����F�d���H������4�����9m�i�|r�e~OM�&�1�4��9ڬ�f^���0�:=9}}���DP~exܝ���
e>��:!�C�yB�YL�lkU#�_�X.��̟�O��B�k�. ���7��A[�ϒ~=t7z�\����~U}v1m����ũ�f��"J=�t��P�
��W��r�����x/��&XFQ�U�ܬ!~Yb�P[��區��|s��?q�������+Ã�߃��cSA*�y���G��Ͼ���ir�z2vW��(�'�9�#_�|����kx�����}�P�lKK��tn��ix�]�����G�B�Ѧ�� ��Yb�MJ�e�s�?Ԗ͛�d�w�����A�� H��x�s���_��_����Q��>�7Ets�"���ӝ��Y�ǆ��憓��"�0v8�5���Lo;b��A���|fEՍ����u��o4\���w[Qh#z�q�أj}mEV��0#5n~�~�)+���D��>�:_?W�f�W1���s�����Q��ڃ�Ǩ��s5e\�R�JԆ{L�Q~w�܍�j������xu�=A��``��J>���*`���.8�{2J�Bc�K4�Y�N_��
�<�x��u��*����Q����\���$��k*��eO,�[��0��<�g)��~��P=	L��d��r���.�yE�:t'�����a��&92���&�����+
ԁ���/1?�5��SsD���O���C��Y��>�(�]>�k ����=`�1X0S$".��O�y��*+34x
�D����إ�2cB-�T֍��+�:5��6���y,*:�Oڕ��W�K�B/^�*�"Y����	��ԡ6y����jFC����\3&�<���,%t��6r���Wy�������ǝ�SǪ�e�{�J)���+d֭i�k���6�߽:/,��D5�p,�1�h�в�G} ����
ݟ �	�:t��a��Y��o�V��h4�%o���������α������^ĳ�D��B�(:�����w���|h�tZ�>�m����{,��ͨ��4�J���LِR0�~�k�~;y�4΀|�N��������ʅ��RΡ��"�,��kO�v�5�H�iD;l�=��sk��m�<u�*y�R������6K���z���Rxױ��ڐD�`1�T�� U�5�1��)���T�.LyFx��(�}��#����"�%V�@��:��.�hĪ<슆%E�wM��>�����hV)�5,@E�T�������wϹ{�l&���D���kc�#{�{�m
3�>�a5kꑀ(�6c)!m�be�+��5KT뽢�'���-O�I�����>�;~���ʔ�a]z{��M)\�5��	'��x�z���`��yd����j2F٤�d*3s\Q��COz=�����b��{����s5��<s}������*״]�i��9�U�)sl�<�/]Μ� ���p�'Z2V:�#+E6��+e'@�h���z��8��}��Np4�Q�Sj{���9��^��˝���x�n��iEq�t�*I���Vo�O˥��9e@n|>iɚ���R������*���??�������y'e)�.��F$k)�ch�f	��{k�i	l_QTA '�)y����%)�>���zt�����P
b��
\����b�,ky����Ob�9��ޠ��n�P�`�+;}�t��NQʶ�4�y��%�X3��07"�� �>j8F�>D��=F*`�UJ��=�]Uޣ�է�r轼�MY��T<	W�sm��n I��6֓yS�Ҩ�UFEnb���ю�.ӣٶ�-L��z:��h^B����*%��=�F���t�����Ի��^m�_OuYԾߌ��F#k�"Z.�>>�H`�%Kr�w�Do�K�(��<���h���HS��Q�az|�h��K0�k�w�olM��e�c�T���b�O��t�X�{�Ae��Ux�GBۮ$�K�޶�✶�(�`�ۢ����ާ��{����!�ƷzZ�_�&!�Am�"����?��9����
�������Mb�t����hY����5���3g����F5�VQ)SqQmkժ	�JG��3:�	��Gj)_ݏ䶎�bo�1R����V]E�z0m�۞���H�^k4K�p�f���@�V�kx�ļ��M�7=&��Zr�L�\�``߀��=\�z����.ڤH����Fjh�T�����o�B�r��y�ڟ��i��.&�֖z�i|���bv;s��Y�-$������.8������~yM�Dh�Φh�7�p��>���)!ַI���ؾ[a�zV��UY��e����QF�E�W�~�1�u�q��b���1��w?����~E.��5���m�ַ�v.K�9�?NC��I�S@U[6A�I.+�AE�f#�E�P��@@��(3 z���5��:>#-��������f<y�2�����;k{oFa5χk�h����H0�P��@��WB�z�M�I��egT�el\�u��=�Tv�J�ܐ{u�?&��T 7��+���y[3��B�z�.�&l�zZ�Vk�4��¡|�cN
cQM^<τh`��1��5���m*m�6�I;;c~ݨԜ��6;��S
��H3>�;����^݃	�Σ{��*m+��P1���]%\��|u��XZ��?�Ԅ��	����)�B����	�O�������
�I�*���zծ�%<r��_#�B����^7��:��m<*���)'t�Z�Жr}�9��w��-��.��B�1� ��K��\L�u�q",R-��^q�'�@e�"_*_���a�X��,�+�a����^���WC�d�bn�P;�1oB�{��9N�H)��a�^��%d
�G�;M=9Y]v�>*�	]Y?�IOl05��b�!(}o��톗���Nw�A)�p!��۸@���L�R���
�Eu���ѣ�=��#�v�%�-K���^8�'�Sea*����j�Py5��l�2˴=��%dz(�^[n��[vUx&�[���E4���j0DpU�U���m(Y��R��$���u�Ⱥ�ٮJ�U=p]S�ڇÐu�Eh☨���_^���\d����,M*u�^�C�bG%�)��^}���|�M&$@�R`��{;J����	��̦�k��Μ;�/�yj�}P�NTh�<��S.����",9�"�Uw]���ސȩ6h^o�n���d�&8Q:�!�Lad����g���K8��)�*"o��pl��W�Q�"z5����A�./�6�h�7�h�ʻ���O�Ys?m�eR�km��(�����ϭ�mK[\��Y?͐qB^��ܯ�$*L<t�Ή�78�!�Y<F8��K��/�YI@��f��$��2�{>����;��<���nh���K����{��v?f���ki�"s_��<�2��x���9�EO������ն1����iH���R�#�5n? ��k���C�޽��s*��+Dk�����'��K0⥏���m]ז4���� (lFf��Pk�)*CNe�m�v*O ����3�z�<�7���j^Rk,K�-��e{���4P&�Ȼzm�tq�J���o/B�;sȆ9�k�g���9p���x�<QRx�a��]#���q��Q����iC|.�c�ųW���&�u5y��̉{LB"C�v���!��3�\�ק!��s���D)�hJ�����I�%,:J�I~���j����. ���޾}�y�Q^���WA^�-�x�ݹzoL�
OB�X�.Feg�^)6y�K��քf)��~rj��Z�Uy���V.�_��J���%�ʫi���T(
��!���C�B��6[)�R>�g7_��X��������F�<��M*��?;�ִd�)��˦��'�@�{MH��3�۶��{�ߤ>���,��T�7K_�^��u��
P6��@�Z�@v�R�ʏR��Gگݼ#�Z�PRy���ѨK�Om�* �c���lZ����W�s��{��a³�'#�6��&�<����Jr��~T����/��.���`��gT�/���}h�;�QcR�q��￴n��w�W��<f�Wj��J�����<�0ev��u����̺?4�g��)ˮ4�Q27�qZf��M�]e�����s2��v)L@�k���5����X��8 A���2�;kZ�r�
����F���c.o<���_5�뚺������fhTX�;}���r�+}��w}/�9~Vw[��zP��A!7��N�UqKh!k��׾�ȷ��&MaҔ�2FE�܆���Ŷ85�-�z�=����� �LЪ![����p���-�YO��fY�LJa���(ps�!���K7�ٴL;9�?q@�>�E���W��G��dm�����)�6���H[����d+��睂��7U�e��xV ����FoH���ۉ~�=���j!�]�:�؛/���E�_?v�'�U{����UٔZ6�ĄMF0�vSx��v��\t���_^y���th���U�>
P��l�'U&����y(Z�10*�ݏ��S�j�\��%j��m�z��Qǭ�o��n����cc4gY�uab	� ��A�ڰb�^Hb؀�傈.�c�M���CW������ȩ�7�S����=6?��z2���F;x��
��Bz��+]�ڍ���{ }"�Z�l�B);���S�4�����c͛�^A��B�"{�oC2��0��ǉg�G��q���4��R��L'V9�7\���*V �o�{R��/�~5=���z�i�#���[e�Ե��e��(���
r-z�2m�U�YEq�P�T�i�'W�{-|ֺk��5�Z�)c����r޺�j_<���j�3�BʵY#{;��Ws�μ\@n���`��x�Kq�5��汃$;m�,c=Џ�g�r��d���-K,�n����Q�F��+�ןj���^>L�;��W�n��[6��KM���	ʫnB�R���%�������҂��#���&3e��m�yx�Y*�m��s6b4y�%�4�z�\zO��et�,��7�~���;ÿ��?����ȅ����x"5��?��&A�Oo�gh�D��,q�݊r��30�M@_;�ޛ�^~�,kCp�DL��m�k��	��d����q�J�D��g�Ƙo�R�5Cwc�4��_nz	��"�^1߹�My�M�_em�J���>��+t/���CG?����>��G�6%X�E�4kcv[݄V����&�`r�Γ�
AB}#V��݁
�*p�KU��4)�ڿ�߫�s�.�VC�K�ӂ�X9b��{[S�=4�OX�#&ESh֌w�VB��R�ȚR�p*!���ߍQ��w���}���n�������y8|�a8��9�;A;���*���i6�`8��oË�lF�t�Nf ���)��<*��Q�y�yTR\��cZ7����v������3N�kc/��-��!��X'�ە��Ä$׳��P��'J�NP�FAX�[��Խ�&p[�fdI���S��mf�a���J�u���rƨw��F�:F��wM�B�R��R�ˆ��AY�/�/ ����V�š�5��~����s��(�j#�c���ɨ�l7�_�^�ųF��a�ʜ�~�O��z��$��:�F���q��t��^K��t55V��bX*��+�>U��y|O�6bX��wc��^�㔜{���cu�ܿ�e�����e�6D���X�\�+�*gL�AnkX= &!��>�1�-T�CC��`��K�?;���2�ub��*�uQ��x%�aD�h�/j����N��6�n?{k���M��Y�SP������o��_C�&O/=�S��<���;  � vk�7�%͞��nn�A�r�4w�n�ȟF�4��8��<�8������X�ʍU����w"�M��U#ZC�K�#{�{ǨY!2�����Fd��7��=��n�S_�#���;����?��z��=y��}e�ڮ0k���pvE��	@��(��5r6��<�EQH�� =B	=����Z݊��̇@6v��k�W����B���c�s���n���	�g����,WJ2��#^���4ή��M�F�.7�@aQo����5���ۄ��<m���_�:]������#�
|賳�C�)��B��nH<�T��f'����Z�BF/21����.�T��K�l^�jv���~j�k�x�M��C��i�;��7�:>���2��+�ʣ��Oמf(��Nb����$��Dq�[gw*�+�޽��t���HJ��+�c=��$��,�I�
j�����%�]�\��E2{�QT
"8�'[�YE��z��.e��d^�:�*�*���bj�� 3Ӎ���b�FU�v���2/]%Iŋ� ����K�����\�,��U�dH��hZS�}-�*G�"
��\�H׀��^�TT0����m�w�0G��j��?4fF�p{Wv݃U���y��2��L�w�^��52�'��S���q�0�:X�1�Z!�c�_�QEW��3(���W�:I�@�E�1Y='H�Fi3���ӛK�E��r�9z��4<�{��ڍV��5���!u������[!�Qyʵ��z�z�vPGi
,��S3#(��.~%|E?�ʆ�|Fj��ŨK�
q����ˮI
�4�RX]{Ԭ���>�#�;&,߹�Ǯ�$z��8ձn������C��#�c{�С��|��?Y��e�p݁�e�/����!�B2�w2^��C}sv�9f��@W����
��|��n�_���B�a~k�ƨU_.�W�TB1��w{��V���}ЈX��KH��I<<�t6t/-��xS�3' ��*X/|��D���t��Job�-�w�᎕l9���ۆ{��3�w쨭��?K���;�Ev%!_�=��B��ă��J��W�:FJ	S�Gypx��#�������O~���"%s�-Mn�y�y_�M����e��	�"$��5VB�<5�����T�^�uK�� ���j-���-3����۵�r�Q��b�1�mA���o6��'�y�(�DE�U8z�*2<�fl�Ll��"_O6�B��ʹX��C�UZYG�U�M���:j�����8�����.��¶v��._c�R"�xg�u�鞴M�s��(Z�Ѭ˵����m����{�0��g������7�A+��XU�^\ka�sKeh��51x�qk����:#���i��Wb�pv:<G$=����(�/i�J��hv�)0[��Wg��W�k�|1D|��ܐ7@5�0��t���t�#��
�����Kjʰu�ߍ���;�W�]�b).�P%,�®����V��d��Z�σN�awK�TO:)�H��}g�ȈT9W����PTk d��+�g��9���9<�dSR��35���^ܼi����ް��Ũ�y�����4��,���?��]������] k��Rmֲ"�wt��EZJ@uϢ��`x�6k�F���9z^~-?/Ɇ�
���̡G�����zL�_u�����댣�Y���{�ĭ�B�>�Q��=Gk���l^�<U�P��k�`ޣ%����������vV�1�Zл�>D9��a���({�l
P�l�KW/�l� �6C���'e.\�ݐJ������|u�N��饾m��i��D?{;%A�;#��&:rYs���В���Oȶ����]%΋ ���'|��޲hh)��j�:k�c��f��<Z�)�!��8�8���m�r��u�%�o!�4�����%�j�����4ae.Ѷ��6[I�av�UpH��F2��F+^�%��j���Y���TI�_�*�)��������fR�C�e��HE����"�5���zԥ)��e����#���IW���ݦ%�M�W��IG�U	36��>���Q����y�NI[{G��:)�yt�|������*�A��=`��P܆g���r�]�b���DO�*:׸��b�2ec�=ZC-�8�3w_�̽R�G�ɫ�W�[`Π� r�ȅt�t��G��[���J�VK�O�uj�+m�cV�X^s��
`Oe�.�A���k/@Jed�8�!��ލ�T��J�D&�y[���]�r�����U��u�[9��l�M3p���yҶ�R,q��;�C�bi�����~�.^��Qf���P�׼������]�zJ�X���t5TX����c|0�6�ɏ��G�A��"A��^������V=� .��߫�B����2WY�
��l岎�CI�b��x��ݴ
�>1��-�������{���.j��?{:�}{�K��
g��=á��Jٚ�]��#n���e8�4y�rB����	��^�
�=V�%�2�
*(~����7��|���a~� ��=�W�Ͽ���/}���{����E"Ԕㅌ�Ӗ���8��lл0-�� '7�"ׄ
�Tȱ�v�p��U��2���Ƶ���`����q�2�eIR��4�D'���
 #��z�7�'Ә�oh���oܓ�Y+Y]�	���nƳ3R�s<����[_��D�f@*#��j���dnу���L@i:��x�Q�^97F���������(k��1P����K>�E�������jF���\��Wv�}׼lE�*ZT{�Ǩ1�)�W#Zm�z�<�� �|W�V���u���YJ�Sk���5$ś�W�?�,W�=��<�1�9n�x�*� �r/u��u����]q�j|��Oh�y5�2%��Ek�����Iv|�$��ک4���u���b�����@ȑ�Izs̧�ep���-31#��! �͏���R��V�uQH~�Qr��ַ�H��-�)��{K.��@��Z�R���㱂Ar�肱�M���������m��y����Q
�����y�Ϗ�w��/����K���Z�K�W$eTi[��.����~/�h4�֟w�V�>B Ѽ�x�V�SI�.jw:Ey�׌c@?nZ6Gg٪�e�0Z3.�N�W�ݐ=��kҋn�<=��x�
�ΘWQ���a{J7d?��к�w�=>�������'A�1K��$��=�n�V��u�Nj��ފ��8,=w�MenQ�ý�����HR]��WYm -23La\L��,��%��MH$��3�����O|lx�{�	B0�m�����P�ax�/�� !�t@l3F)ڵ�j�x;z��n�2$��x\�^�� ���߳"!���(�b�Wͻ�y�m+�}g�����US��\@���:���J�֋^�V��@	xv��2�*)�Ne�3�l>����
N!hl���7^YS~/ec�q�P0�èxg��MMiQ Q���Nn&҂����^�K�YuM�窀����[�)+���j�J�;k��o�.���+S��ז{r����=�l����VYiy�Ω�[ՔݸU�������Elb��66��B�IM1����E)��a���SbxM�fK���A[""S1^�Hw�a���7��0��(�Ҁ�h[�iL���#v���W��rx*'�@X\{תUMO�g�ZQ��X5�W��
JZ�ܴ��ٷnc�D�N@ش� 7M��ē��֔EmϘr}jb���)��=Z�g��ޫ���j���Kn�@����r�	����p�X���8�k�ڿˡ����ۯ{��G~��o���'��ϔU�� G7q�Ȳ�w�':����S��,����Pt��.��<��9�JW��ʼJ}v�Z��ݒ�����楤�(���m�\rX�>��CV���<q���(��u�Lϧ�6*1IHS�\�~�1YO�x�^�����7}��|Fp�ŋ�$U�	~9�+�Q���:&��B2U/x#a�l@@
)_� ��鱨#VKj�j��-�tFJ	8o���M��]���E������	�y�y��O~�Ӕ�m^}�ᩧ�f0��&0�rO��q��-���T膱+�Hge��7���q*T�9�x�h4���_R0�KB������s��R�׬�@�[�,�v9�z�Ƭ�o��wc�tLq�e�nb4�jVeC֓�!<v�7�w֫�+���c��ެ��I�t\n�n֓��+��<���n|�=�=��yo��e77i�+�3^S�����GԸ:FO
]B����W�\�cm/f���n��%#
��A����B��Q4|R V�s��)���U�P�0��
bI��j�M�����0Ÿ��@�9
�F?R[�����9*2_�������%Rs2�z�o�O�u2
<`���Z�;E�8�m�\��kF�
8+��ll�o�p����G�40*�P��Nm�y:kc�h��e�)�kQ���k��9�~t$A�Ǽ�fER�g./��������ܦf�u���n�%~�?�(��Ɠ���o��O~����εw�
�mM��O�K!���n���&\v����=,>������r���ѫyLSAjn�z7�S�h� y��D�aK0G�E���jy�,��N��j�7=��5�^w��%�J!�ICZ��$�p���s͎9}�\@*ָ��>O�tۢj�Oר��f<�^�8U��e�w�<��)�cJ����ޞ�VaƉ����Q��W�x��p��iBㄉ)?9:i8��+
�+��u0�{�9�Co��Y 
�e�����KW��g�l��:k�>Fu`���=�ha�H���$ż�B�:�fg�����&-��Y0b��3>�ɉ�]θ�<�z�`��I�2��LI$j�D0����;�@�}>��5g��)8}����S�8������K ���L�b�U� �8�\]Wr�^7�3*�������`��)k]�6��O�p�S�Ѱ��2�F#i�8v�b�����V�W�T��徎����;�jc��*��h�����^���ⶣ�y�l�^��,O��*%F�>3��ܯ�o�3ctdl�0�deT�'��r�P��!�=�$+C�s���|?i(17��ƍi���:p"L	K�U]m��Ϥ[7�X�ф�yp �)j[>n���^l�`�#�m���^�p���]7&�]�ʯ@K���*�3�\��9͚�TH����&�Z��I�*��xk���7���ٗe�u�wj�5O=w��#A� 	��Hɑ,ڎ�ر�(�Z�W����%oN^����!��Ȗ5��(J�8�	�����y�y���|>{�SU���$f�]`��{������w��8�~�?S�a��7Pָ�MGLL�v�'{�;8Ws���_8�.��.=v��O<��^�I�r�iC+Nc������gs��{UH]�In�X>��Ra�`���eБq�ߏ*���ռ���11�AxP��ī��JoR��5D�H���n��Nh	���	�<�!�:UH��t��aN5	AG�t?1N,��_uPlf����֙�����|t= ��M{��(��o}zz�����(t����x�ާ9�������`�" ���qOӄ�O��b��&d5r���	�,	oI�e�5��͓�C!7������dx�E�t��s�}9:�eD��
��e-]�2��z-r���t �a�<K�B=���~T&��ғ��zD�v�pI��=nz9b ���ǈ'�/#&�Z�'l�����
�\y��K!��3R���Cm�;�>��6I�Mf�x��Di�h��8K������ @�%!�#�.�>P�]N��^��=�w�2���	�vjl׹��$����iNg|w���~"SIATi���9�N����?YϞ�^�=�)o��3M����|�^ON���&n������om�9�y�J\E)��h�x9������{��l�׾�$�ͣI�/���
��Ԅ���=�1B��h�#fp�!�f<��D���(��c�mD<2�������*�#	{D����� EZ��=D'H�"*�L)h\YZ��Kܞcq�b�rL�mD����8ׂ	YȵiL����ަ5����w�R9�FI� hRcZʎN{ �ďr�I!�ւ���=w|��B*t�������w��ݿK�����z��<�N�hݛ�R�_g�wT�S]G�7�^���oGO�E:^���*��b��ӷ̹��[�Cc:A�G���BID�7`��M��m����� -�0P2^vH�SQ��^��K-��c�x^
B�#߾�n�GMٽ�����[�6[�k��ff�bn����m�0�ܻ)n}�fl�a�B����/ޖ�o~�s.��i��4߼�$�5<�ȹ������g�����m����7���w�ſi�,Fx�����[X^��:}�/##�51�NR�*���R&?�gM��5������_��*�4>�/��W1,|�Q��Q+N|m<��*<��Fl���]�G�ߵ8��C/x~&L�قYld�#�����̅�"Sچ�����4��^��|vP%�k4K��z�B���I�"��������w��tC�f��b�>�X�_�܈�5�=��)��}��#L����k�e��+a�1��s�~�s�]ĵEt ���;�	����{��Q�g�|6Q���y��O@�%,���\v����D���W|�Y\�on��sf��YE�A�摪�#��ܼw�=�1Ҵ%�-k#E�ͣ�H��d���M����!���:rī%`��`��p���O|�FK��
=B	���@�}@ӢlqluG�~z��s��*W�Ja�V �o��i�\�F,�tn���F�%r����ҍ���m�p����p��zpW�D�
��4k�p��l�\;���R����_�̧?��_|���k͘j
F�q+�:�"�ruq�� �E��S~?���Xy�.����R��Qk�;g'�қ,)��@P�����p����E�r��k9����w�d���8Ɣ�P�{X��O|2����nld%sv��h0i#	B� ?���;�34�ѪwF�!x�D�s�3��ͽU����ݏb��m!�ז�>=�wwP�F�<c4Pio#�`�����������e��fh�SF^�F��������y�=J�h�y���S�>�<���{��a�S6G=��[K�����f��x�/�I�Hң34m+�"������3:�Jo��P8P1:҆QYg��e|�Y�����mg;�"I���m�S�a0{kgiZ����2�c=�.�N}�R�ʳr̤�0E��������A3�ۆ�U��"�h��$�\��k�	��Ur��Y�$4������iC���Q{�3&�ah�y0,�*m�w��\�^z-�P�i�vFa�{��J���!�H[D�?�;���z?�9k�� ��<K��|�:c����6��:�9�Uʫ<��ʇ��MQ����Ƕ��Pj�?��盿���As���w~�f���!��|�f���g�ɕ���7����4	.D����U�q�{�E�u���>װ�g��OC����͘q*��j�l,�I�ݧG{C鵻�$�EU{~8�����q�<�����"�(�Ѿ�9.�=ƿ������T�t��r�������C����6�Cw�9ʚ0�GF���L�c����Q�������޹�Η)�z6-eQZ� �X(��ܝ�3��b�M�  :O�g����zj���G�~4��{�ߏ��'?6*�I��3o������Z/�56�^[��Q!9X#�z���� �������z�,r4j �������ߧ޲�<��#��_jVP��^~�ы���w�!Źs����6|�@��K|�M�'���b�k}����-��Q��?�'�L�4���Av������wx�4A*��ƕ���7�n�^�_��fk��/|�����o7�;�,o��L���~���?�v<[7�ʧ�e��yq�z*�܍��}��ƂҊjy��9�p���X��7��w)nOj\i�v�IU;�$���G�l�
+j�go���ni��K�>�]�a�D>X>�$�/\OˈI*9�~��n�$3�u�S��D5�H<�	�����>
ì�Y~��i׻ޤü�óm��#�z���o1��Wǌ�k�N���E�'1-�B�p�Qw$Y�%��}ֱY���f3݊W^G����|w�+hSU�W�!��f�6��ڴ�!�k	c��"#}���C9��V�ȝ�Q�L��n�|oǶ�e�V�s��G�n�.R-2��GJ*�0i܊Ib��8��탧�@�L��*cֹg�!¬�Ñx�c��b�H�tI�4ܝ��\1��p14㕩^��Zq�� �M�E:#y)��E7�s�^�����ǲ����]�/GbfDF*��d$G������B��|�"�N��k������7�L�\~�М�����<��u�5Q
�`�����j��͛W�����������,��\��W���*�����b�g_K�4�8��1:��z�H1.�nPDw�N�t�Bl��u�������M�ކ/����γ���S��Q"��Vtk�dC�ױ}Ӓ>,�jC�Zˎ���6�G}N����n)���ԙ�a+�G.>�<F}�Y���k�gt��SgC@=X�n��v��H֭��lDH/�1!�z�a��/\8�����͝[6��4�y��aA>>JN������w�S_v5���B��޿����1emO7���'�'��c�P�2B�
+��a�C�J�P0o#W� ����9�
�}��-��!L���x.
#�:�|�B3��:'~e�6Nw�0�{�s�#qy��x�o�8�����1#<1U��P���u����q��p^c�-���vJ�I�==,יU �B�㤰F>S~0jԡ����#��W$!��Tg�Do����фH�ۥϞ���7�RD��i<��u!`�U�������du[B7�z���;�u{;r��B�������E��Ѽy�=L�������q�vv˞���x���"?g�(�ߧ�g"��xQ�WK���g۬�m,��ք^���n�V]Z_l���+�{�7�i�Y���"�z����Vי�
rr�`�
�XnYFe4"$���yn$ͽ��*�`���q���xSWØ{�^	m	�4�����n��`��H%���(�רlG�O&"��Qޚ�6��=}Z���%Ⱥ�H/D�Q���#a$�����5<Ԝ\ȱ�+�c�H��I'�8����с^o���J�\�����ԩ[���g��G����>�~��]غ�LB@�J��=�\}��&鄥Ū,�)�±��b�U�'�CO��ֈ���?�u���+G��]K����#%�?#X(�<#�IC}w�kO�5�2�^KE豣�*����襴�?�GX�=��[���%�p>sU*�ȡ�8y�Ts�q�
�S�<�,�>ǆ�5F����杫7���o�e��ɨg6��W7ќ<s�cΠ�7�w߹�b_aR�B�����:�uȆG��$��������.9�7�4��/7����?�̟:ռ}��8���y֎��
;1�, �h\k�M��4� �О�����'k��4��)L��,+�^�k(t��my;J=��(��V�����l*�\j��x��3���ꈃ�u�����K/k���!	I-�:(��7���i����0�l�bL�G#��X��kǝ�P�~�5l2,�sJ#4�D&�(��ni
.K�_7l:��}�����l\��慳�B�b�HI�V�����_�ͱ��[�/�.�q7׼��G��`m�oɆC^��k�kP˥M�gɱ3�`�adb�Z&{�J�������o�ܻC_vHj�]��
ē7JC�gs�~c����z3C�e�����(�h�yWW�ھyg����f����� L(�rd�^��lf���}��"<����>�� =�>	��6%�q%C>d�F�'øK�Q�j�x���0�N�e������B�{�T����Jz��T���%�HDo�g��C�9N	��T��|�4��[4�Ʊ��Z������x�S���G�x
B9�G
�&G�y�Ԃ��w�1��/؟�	��ӵ�׺�kחZq�%z���ɯ���Ʌ�}����s���x~�ŭ7� �����*i��¢C�
E�Ǉ��\b~���BG�4B���������V�l�}XcnyH�F;�P!�h����rRkz�ȟ�?�k��g�u�_�淛7��l��2���̏����^�����Rs�)n��a��_~�����C(���:P���ϝk��o�6-gO7������?�I��dS{� ��{-<�1�(�Uo�� X�#4y�� B-V�THj2��>��%�>�T�)��d<�x̆+�#ސJc�TũS'�ڲ�W;����r���9C�wQO�^|�;C�[?�)�%_j�@�lݿ�A�x9��}u7"��]�B�1v�#��g�G�x�<G�s ���  v��s'¨[�q#�6�"�>��J4R	��P�vޱ���;6�!���-�3�����9�8�֜��~��Ј�[hD9b�m��kg�DH��Bm��S.]W�a~\�=�����`�5I�������ޛ?{����:d�:�ha� T:�z@Z�އ 	F!�LS��co8�O`��i�Djc7Z�F8-�/U`|.T#���s�w�hʴ��ua�Cb���о�=�H��k�p&�so�h�`��V�����b�raa��S��{�0z�ʹ��0N:^�21�g�fHB�xA)sM��]��ht��6�Q�^�������}�1�K�:�B��1(�u�J�a"�`���pB��.^y�����"�{��_�6�?��k�~�������]�l���>3��!�T��3�jC��wܒ�R<�B<��2����w��5<z+����l޽����vm.P��EڒI����G/<��>ͰZ�b�}v{c ��� �dhSoh��h����~��<8�Q��>�C�PzI��l�"'ڇ��&�8���8��Ge��<x@o������揿�fMB�^o`��)���j�Y�q/f�!�c��U������	šQ�-���O����5�2B�Cd&��d���5jӱ�	��mHv#��� w�ݯ�"7ji�ރ�D�f�;s���KHC)]�C��]O(T�Y�U�&�T��4���83�5(Reg����&N�a)U��a�!r\Sg��|W+�r�&q(�P��j�[$�E
�(�� �m�%�S>�K�K��YcLPo������f�u'�}vx>�[�N��ʅ}�-<�;����5
x�sv|�h\����B�����(0���@C KO��:�{Z���B��O�e�G�]���:��U���t$Q*J4S*?�Cq�U�;��hg�$��OC�&���Wa�߈5�VF�Qe���u��#�;�Ht��}Q���a�o�N��:��G�&Fnlȣ1���my���*� ^{�`��j�^��9�{G%�1u���s�F�H�3�uGe��&�7׉�i � 7��	+����^:�O�� ��'�ӈA8)V"P���:���S��P�g)������qF�P1z8�B��gѓ�)�B:#X���q��,t��/���	�_��^�r�%��]���2��x�D.=@Wwn�g�nT��RmI'0:X0��U�#.�x-?ߪ����ɼ���uJ�!uX���IH䷺\q�)z�FO��5_����^�\�jdW+-��|���l��?j�ܹ�ܼAv����L���<����m`1����M��k��\�4dv�]r�!��O�FA��n�o����|������uE%��A4 sz����;�|x�\�n3G�vgt���;ͭ{�x�vY�>ˣ�޻�^m���ퟆ���(�K�����;��_��P���9�����g���g����}ʯ�7�^G��	G�����2[+�՛��k/2���^�b�(�g���@�4�O���)��}��(� ��屍 d�?O�^G�)rMź���tJ,�8nx��HA��L��F2U�"	U>���m�=�����u����l�t@�7�t�{�����G�g?�k��T���aj�gK���	q��:���ll�JD+r��_�(���d7���gG�Ď�����dx��|��c�I~��6��� ���f�y��m�7�0IY|>���L��U�*i���H;6}'[܃]��h���p�I9aX����2*��D/u�ϝ�5�o���9���1��������s	4�~���W�������Ҡ�%63��|Ny�F*L1J2�y�vfA�T�4�k��2)�2��4]w��Ix2�E0��
V���K��*���&�D��{��{<�0���uי���b���N��i[5L�f�>�T�L`0j ������¹��'�z�&R�1�2�p�=;�L_��c%ω�C���Ɍ�#���,��m���˱P�M=x��7��k��������y
@i4ei�󈨻�)�?�uif�]*��Rb�l����pQx@��b�J+[+��t�o:噬���$�a�'f��^&(����{��6?iX]�#kWCXi���l ����L`�z*_ϣr��娤�̑�ם����A��y����8�ę(g��
Jr��,k�C�������^�.������懯�I�o�}� s�J��L��g�p͌��XgN7���f�HǹՕ��������!B��v��=[kd��\�cey�y��+�_���n�CڻuoeI�����C��B|�f��1��1�>��Q�-�7��<�(����͋W����9r�Y~�W���s�$��m*+{�'	�7e�ut�J�,�:H�2�e�s-�S��NC�F$z?]4I��)T�ڏ�e����1:֫1��"τG�jTH�:s��fm����KЮ��LH��e���V�?���^��#z�����5w�>��k���������0i��w~��f��^ZZ�}e�ڻ�ܠaJ��w���j�S?��#AB��ԑ%f�*M�s�qϸ�:R��]��5��g��?{��5����f���WY���	l~�8��'��x�\L{��p�z�5B�o�%N��_�00�������D�a���p�^�לY1�֘JْJ;����gg�rQ�΄)�|p���������Kqh�z_��4�n��e�ӧ�6��?����=������i8�ϟ�K���v�OK���x�x�^Í�Q�K\[�jr��I�����M��ɺ_�T��{8)D
&g��i�T3C���g�O�;s�Tsc�k�����	h�2��n��2��([;v_�B��T._���/��7>����<xx6C�.��=�p�1�<��Oi�f�N.�͎�SX��:e�לy��m�;B�~�ͭu��2��q��F�cR��P��zZ�Z�6����^�~�T�%S\�z:vO2g�ʜ��dBieu-z�v��h�pax
US)��?w�酱�5��y��K<ћҫX��jum��x�=���Rs�@(����F��!��qz��d��$��� [83�d3M�{����I�+�<N�׏��>z3ؿ�Ԑڅ.zr���̟C��Pbޥǟhnߺ�ܿw�&�o��+��Լ��_n����Z�n���%/��ֱ���E�Y�te|�ĮP��1��i=̃��2�>�f댍�I]�#�RqxHԷ/���A@����ٍR�w�y��6Q��a���(]#��w�}�XV�|�\����d�HG*�n�)���i	��>3��9P��	p(����jDo��9��<�B��
��e�U��Jɘl�0�r����r���Ϝ{Kv4�3��<q�D*#PAZ��W�i	��R�<�%�,E�{�V���~q��ѣnB��;���;�M�"okԣ�/ǈ0|��7ud����Wx�m�,��R)g(7Yb��ez�ɺv���+��c�l��KD�%ԙ>ED&�[C�w��r:��yD:�VUY!G8a�a��Q�x���ᣑ:��VXx��v�k<Rg�y�1.���d���>�>���+ݐ�U"\�H��&Mj\�aH�~���z���ݨ�Q�q�;��p��L�<��M̳/�U ����BD�B�[��
��������K#�M� �/s��9"Xܛ2��F�~�Ȯ�P.R\���S����C�7����� ��[�Bu=��\�����<���Sa�u��a�4mشP;�̕���m^8_3\G�Q0F��uu:F�cG�;�}j 
l�˭G����~�f�����)�]�6���V��I��b�Jx�9ElOp�\�3O?��C����u��z����*ђ��@�4'��W�D-�<�;`P�*����+���[�����?|=�h��]{�5S!$�Cs=lę�y�n'���#�t��50�18��ﾌR��&]������`���A����Y�;��
V��o��5�׿�����|���@����y���w߿׼sa2D�{��5����(�9���fԟlk6�<+�(r�>���!O���G��4�j���k1��0r|j���Ț^hz�9���O�A���b����8^�]��٪�<���p�^�2]�T
��7z�%"��hg4 	R�%� 	-��Q��Z�t�g�Q0���}�{��#ͅ˟h�=�l���?͜���'Ϲ�46�5Ԇ�e�o�[�pm���� �E�kX�~��ݸ�u��p7�\Lb�84���C^3Jś_Y������@�ͧ�����z ��2Jѱ�;%Fl4pɰ��%���a`���G�Bt-����:�Z���.�֥	BF$cr]>փ�����fWF�,i�Gh\��>��@�U�ǕJ*�x�i�E�O���;ʓ�Bf�|��}�s}v�z��4Gߦ��|�aı��дL��9����tc�� 7�v�<,�nu��<FZGtd,������h`-p�K��V	��qQ�%)�S]���e��F��0����ĵ�^��V�3$�R:E��)I�C��SA<��d���~C6�>L�}�e�ܧ|l<to��ŋ��~��~��_�Z<�8�lx6�;��Ps�-��"��B$�L��.��,H���>��[!����IO�:!�5$r�V
.[wZ�)�� ��W~�|�s��1=^3Y�d����M�Q�x����{X����_~�2F����;������fS�v�^�ܴ��fJˉT*���*pC��~��#��ؼ�d�oSC��z�ܬN\�%to���ר5�<nn�c�Ż��^Bl4'榸�G��r���*�lj� K�����=��3͕w�mΝ=�s�^����{�o��5�8H�e.?J�ރ�F�ʞC��%����+b����WX�5����_d^�B�7y�C	�$��ģO0��"���Tx�
l�y���De���yd���l�3����g���n���L�c
�%BZ��7u�A%q�4Ó�2��������mv���-y*�+:�+:�2\�M��z�������Dֿ��Ƹ&0P�R�{�TP�<����xt�
�4@�gT!��S�������R��׽�Cś*��a�λ�4���ꗰ|p��s�M�!��?e��+ �x,���WǛ	���Vct�t�h�t��e����}�?Ԗ���i~���"��r.2]l�ċ�l�2�3ܧ�Cy�z(�}�ʠ�@n#��������2U�Ai@���5B	e����G7�Svz�"i9;E��v`�X>i�M#F��&?}�1�V��ȁ��.\� �'$@��oY�*�SPF-��*�`�aǽ<|�u�����PNd����Y��싈���x�� ۩nxx࿟�{��t�:�m��q�'����WSo��7=�����d\�*�С��J6��V���v�ux	*��g��usG����J�dj����z1Q��.�6�/�oWu�BE���[��zv8�#BV��	)�}S(�	6�ֿ�H�q� a��^��g�m~�!�0�/.�n�U��LY"�72���dS�QdG0-e�7���3��M���V��«�ԃKg�s�ᙛ�X���U(]-x=G����Z��f��Vs���4׮��\��Ǧ"�֯�V<Ke6׷��$��=�pq%�1�}�3��O?Ƈe-'����[5���]�C����pvi�s5�N|,�'�m��6L9�2�����N�����X<i��?	>=��L���qbclj�9wz~��X��g=V���;B�5�^�8u��J�{�;����''�)��D=p�lF�3֖�\r��M8��7n���й旞{��9��߰r�.`D3Z/�[k��[���u�K�X���K��εJ4��?�l?�.%�Z72�Fv{�v������a^����&�f�8��!�{��y�q��zޡ{!�vI����;e�ʾ��7�Pm�U^~�[7��=sv[Ø�F<1�s�˸\�q��MິL�j�K��(Jk ��1�$�QV9e��DK0z���{�ܠ���<I7�F�v��Up:��c��9��JA�t��_{���0m��tEK��g�g�<��3���&����SZ�a�M�0"�٣unF`���1~�������Cw޹F����}Hwɓ�bX���  �I�1 v�$�=�G�!J}-��8ǡ5�>����X)tD��/����޹����=>;�q,�֒K?pi�����R�.sS�rm=����Q���!�k919���:F�	��Ó�i��9rz�i)j��nQ! �[
��)7!���G7��v��<TԽ���;F/�GR�,�M�a?�$��J���tu{��w����:����}ɦ"��� ��\���"tsS�}��5��&�-1eM�������r�+^�fQF���ԓ�4/>����1�2���W_��N^>�O�[O��l�;�V����|��Q�x��K�����ʗ_ʦ74�09��z���W�`hc�)]>2��6B/�A��yB pQ��B��SA�:D?�2�%� ���)��I����`=L�6�?~�R��(��òw`�^^�
��O�z��G��g�'5���x7mM���T�l�ȋ��_��F�����x��k�B������O=E��ts��"��&7	%�`RC{�-��]��0V��(u�9���1��v��*�Nٶ��S�b۫��?��[�|8�ۧ���(��?gX��y�qE*��g�7��"�B�]��gv��$��?4<~��ɳ��bDmӼrx*��T��5��=n��T2�Y�7pa�u`~~��Xo*F+7\�A���ޛ�$���`�1�'�6kr)B~�b�=)���12�b������H�$J��1>9D��0������$G���z\���i�|�:\�&[=�,䤄R۷���u�~�a�G(��u#��ǝ����`��q㔌ҋ�	k6��=��Ĝc�u�:^��իW��~���X�_�9�y܆)%Z��	fy*��n[/$���e쯻��⏥�v��nY!"�Y�VTt:>Cr*�l�ϼp�k���gb�e�z�a�g�~��C�|��]�ܧK�|,�Y�鲟͓����UX����-���S |�l��~ȆԚ=�dB��6�2��R׋��V(�$
z͹�N��{W k��;W��5���G����wjDq-*!�q�(|�<���&����Õfx�Q�\�]��3ǟ���bJ�|yy����#?��o�Ҽ~��T�j��_iN/�i�]��b��UrJ�lQú�@5W�Ad6ro<?���l���<d�g�>�H\3
�V@)��w:%r�H�P�fs��у�p�')���eY]�յ�ם^ZF�|�3fb"�zy=��������R������!��^����w����/�����K`u�����J_>��
��O]���//�u��ur��r��YD�O��`���&�>��,�>�A��x�u�@(i��ID=���Ͽyd�S��;�����ȏ>���M(Ep���"�5w���5��!.�h��k�����ll�ޱ��s�-��Jn��GK���ƥX�pA�8at�e�.�=r�`;Ȅ���r9�{��T��d(���!�q�^v�-��<q�L3-�ޒ� ����!Ah;��C�є��K��e�|�K�n���u���r��ȑ�,/Dއ�U��<�I���{"���0�|��gX�}~_#�O�܍��"�v��^%�؃O�\��#5�5;���8�7u���W��/�����g6��';�\&q�&n���G!OR��`�=�r�a�Oi�ƶK���T��26Y����w��<�DZ�q���fX��
�ŮG�z&q]�����s�����i�q�����瞍\���uk��{�)N��ajx��o[�v���t	��>����GH7�Ru�VO6s���P ĿTT�d%�HV��`����L�a�u�@�����/��4�hhX�Iәw�C��z��m����(���?l6Q��u�p��vg��à%g��t�ù�����fh�^�D��;w���u�I28�Լ��¹-��")�1lM�����|L�B��Y2h�,C�v����;����ľ�A$rB�`>!N��<������4�7�8Ƣ���ǰ�9n�F���$I�kc�)��Mmvv��=u�9�~�d�"�L�����2Z��>C�^*B�>��\ �#���|�`D�Z'��_a��T�"�z���kD:iU:3����OC B�]��#��`�yu��܅�;�h�������M~��G�]���l��������z�t�uQ8��ѿu��)�X&�%��իH��,��n� �����|(Cd�GJ�Tp �_tW�?��w�fɛQ�7����������$��p�����8��zO ���'��GY�VHl�������4���}+64��c"���Q(�_͡��]p	>͚S�dv A9?�|{�K@�;5r*�Y�����G�6鸧w�	���.5��§��g.`���,S\c���&��0�#�M�1ׁ�J��1#'m���?�������[o���7���������G_�vwz�~��vdX�Ji7R�M�OJ���(�|w*��ׅ���R�'9UEg������nkSUzZ��o���N��>m�Q7��,����G?mN�3�܋�b����h��v��Azb�tĩ ����c7�?A�°w��1Bɩ��v�2���|t���q���k�L�<u:Y�[���#�^��<��q�Q=K7�����|^k���^�*��k[�ܳ!���y6�F�����벱���G8|}e�z7l�E~��[;\����c��$�-�J^�Q�`G���x�He�]�8�)��#�w����\���JE�W7����!�%�s��Ǔ��j�4���d��g������o�x���O~�q�@�EHv��=��pNC�>'��(,���n��m����\�Ao���7���g�ˏ_�S���o."�ei���9~r�m�!�G~��m�v|�*�a�ƙۻL����M0M���Ge]�r�Ր�Ǿn�����so�������+���h�'��{0�v��%F�/��G�w��Q������G޽�{=<�xV��������N4��$�m�0�YEA��0�c�˨Lx��%.<y�Z���4J1A�������tOtf�c�8~o�tK]�T�7Fk�W��M�������.uhl���`s��4jb*�r�ՙ�8OCsxġ497b��Z1�4�nkVz7�u�c��vpxtbj�ejl�-�d��ټN���g�w6����4����^��j������0��b�l��Ϭ�_�_����Cy����k��O�x�3����c�A��r�k(�옵C�h�j:7Y(:7d�@���h��ôb�l�����6�B��:1&�K��[�Ӑ��KS���(��gRK]'{]�<��6�֛��A7�w�4�.]���s�Vay��nR?��՛��Ս����ۥZ  HUIDAT�]KچCs E��ƹm$C���6�a�g��i�)���'QGJ�v���åuڪ���;����v�G�a�b0�������^]�)�3j�ǨR%X2���[G:Ӝ=�u�����8�@#�.u}��J�c8�k�)o�(s�Y�gas�*	���n
�s���G��e�*N�N�Q����K�)�i*��	@��eʆ�	�0~����`��S��������,�O��g���\|�R�s�!sb�1^a����
&��5�W\��g8��zΊ�x=S��kع�F�N�7kͳ7=��f�Ju�F2��=h���5�L�"���Ŭ�e�w�4s��{܊���`��rnR�/j�s�v2��*ǣB3��ҋ�m(,l*��R���7�$�U�g���{}��������	G�L�w{��Н�{��U����z�aZFz'Y�9�������vWf*/'��?FYbx�F�|W�F�"�qzvz�Ү{��d����F��N�M��E�����he�;91��n�H�͕OQ�Q��k� ����=��<�ϣg���5�ǭ��'k̓+D�Q���������%/��t�SO?�l�
��I���^�~��$�v�}�`r���w��${f��2gf���~����B�+��o���W~�W��������(�q��a\E
D?&��G������q#�s��ݒubr��0d�anM��XLU�Z_��[OU��e%t
9��ءl���"��µ�a�|���Wv����{��w�����c4�җ�D���[��х.�Ʈ;��H��IbO�X�2Iݘ�a8�G�R��Y���2�C�/>�x��~�y���j��g��^�&�,�y���u���lR'J� %�XC��1��k�������v�2�l��2�9��BIwc�Y��w��H�FmXh���c�q6a��:vi�3���/��1I���Q���|tTNvW�Y:ųرL(�xX�U>�K�)Y��+N��v��`R�����8?�vn�k�k�u�`��>����Qϫ�Z���{���U�P�a9�Ŧ�Vb�_Fc�ퟎ1��������Jz�b��t��:�W��lךs�(7%2��8,a����T�rLI���ڟ5�}S6��s����-¤��#Y�1"n�1b	v��4��mj���q|��c����o�1�����|6y��{Z�m�����������ͣ�L�V�`aF����n�%�BN��B�9��� ��8=���ud��q6�r��>.q��=��x�s��S��)��ӡ{��2��J�,Isg���)����V~��"�#;�g�-y:���%7'K	^7��mSNe�ۻ���Pf��ȥ+��,-^M��5�,=�ه��P����q��%���dD�8n�N�7o�n>�y����2�떽i�sO\���n��I��5�FPE	ɱ�:�
�'u�ɧ�����o�ӥ����/���כ����6t!��UٹI�D���Ʌ��f��Hc��ް��4&!p�N���.��b��<q��Y���e��d����܃R.�PZ�jT���%C�2�������9m����4�Ce�h?�*����ߣ����L���"��%l�0J��B ���G�"7o�Bq,E�n{�u��)��d��4��ܿ���� �G�J2��KO�Y>�\�v�9�7��M�g�w��3of_k矽�w���X!Ң��� ��p��L#xْf��ϜXEvor���k�lO쟊����)>$����>�`�}l����¢]G���Q�J_3�s ���!?ϧ(1Ϟchu�ڔ���Tv�`�~�l�=�V#�����U� c�ǀ�qs������~2	�zi��-+��w��j��=*$"�ӯ�����Mw ���K�A\D8��C�� �~��t��ˡ��k�\�:]��Xt#���ꆸ���t#�_��:ls;F1) x�ܷ}�!�]�+>�9�_�|8:�U��NH5�s��r�=����:��l�%�ށsX(y�~.���EW%�$hp�H㮍C��{pww����� �!H���ڸ$�;�7�������թ�=���s�V�����Y����E]׎�@b�׊�]���xog5J���ߔ.��!��x��������<=�&�Ȕ���˅�u�MҘt�I���Į��_���n���n�\��)~�p�~:��2o_��w��s�<��"a�iv<E��kO*:^NoE�w��⾸g�F�`ҭ�
����U�a;I9aճ�G Kl�}M�S�5��ou�g�= �I4b�e�Mv��%���#�<�ȭ�
Q㺞}hQ�ԩT�0��f�Zn�x=��5�T��� v}ZǍ=~a'�<;�F �ɂ��7���� �*�`���Roj�NJW�Iz�W�x+�V:t�S��Nlj����⪝ ͚�m���ڙ��B�hL�.�儊PK܋���G�9{v~4�&{�3�ݸ4�:W��*�+�o��8ӋR����q6{�L��J���)Ͷ1B6��!���I��e[u�g�v�p	�J0�`��0E�JF�B梠��n�O�ȷ�o��"q����*�H����m�/*]֔����8$�u�j�=-��Ƈ��w��`���ˏ��q]b��I}yΩK�pJ[���<�/�$��_��E$;�aKN�-aKN��&��Drrrh�=�P���Nĺ�U$O�G+��Poq(PCŭ����Ϥ\6)#>n�K�0��1b%e/BW��U�4B�#��k"��e���+�.^�E���T����ާة?�6MZ�������㢶�I��3�m��'�;=N_���8?+����%���t�jcK���A�-��
IDC�]K��(7b�?�����~-��M�r8Hز�E�?�^O�ǹ�H��:w���y��S�Kн�5w_��W��H<E�g�=�x|����S����t�v[��şQ*/_K��D��(�~~�u0�����u�
�LFȰ"i��l��p����k�p��<�Eq"��;4�
nI�=,�(�qm��|$�L��!㽒� ��E���=��~t 9C*F�{�nOcCs%��L��\��|��h��2�(��J��g�J��mE��ց��h@g��;b�Jy <����-W���6�y5��A_殾�/�'-/n��������/��?-�a>,��H��X�����Z�5�	��c�w�fhkw�R_O��2�6�$���mʲ)�]�>���6�����]'���\����/�D=����Q�LD�&�����8��mG9މ{ަ�/��B~���|�f�
���uSc��w�k�@�q�N���&����e����Э��(�����71C<�� ������o����Asu����s�ߐ�-C�[�c�LG3R޶(��y�����H�~C=E|�}.q�w'v���6�n�-5a�QS�m�����������ƀ�K�GLB�<�˔��"�zף���w�����E��w��c�D/�Aa
����~9��6��?9K�G&�$�H��2I,��4��ծ%�c��{�R"�g�� �5�lfy�V)��59�Y9�w��A��1��1s���Y4Bu����F�\�-��FBt@��bz�֦�p����aZqy� �?�\�R�ꯌvwٶr*Lv�s��Ǌ(�ħ�4=W�8�j���K�$B�flٖ)t����0�*���L!5��W�w.� �i���V�X΀�{�\&%!�},�K�}���MX�B�駅R������>��.��K�Uw/�x���f������7�d���ͤ���l���ø�p��:ŔX��@���/�d��������;<�i�}���:m,��~a�.�H�����ox�������woA�����<�1ғ��Vγ=���>�L\�x!^�Ͷ�<�4�e-�2(│�����?v�a;+����Xt����Jç	]�H�l�&��q�͛����@Z����[;X��KS���������Y��@�D�'���!v�M������#7H�������<��\�����{�J|�������6L͡�������-���E�KjC�g�A��V0E�oc�ݍS��>�Dx��{� =*l���kd1���A����D�>�u�+>�͗�ud?��=�[$��d`�4�U��Cy|�%���$?��Rr�8uXDޣ����k�"O�a�"��`d{|UX��4�����T)��vCO��{�Qf�Z\t�WJ���q�*I|�򟍸h	���_�~�����%\����})�Ϟ(�bqsB^���	����J��s�R����M3����ޕ�׋r�����V�L��zʄ��Ϧ�ĸ_��"a��<��o@�v��ߵgu;�L2k�c��n^>�(����S���N�"�}6�?�������f�ݚ�?��H�PSf՗�k���Z�W_(���W���>�i$�M/dA=�����	;���O784�H0��t���8�"q���#�Z�ʐ�1�F�E�^�R��)�����:�Nh1����ۚ��}&�֚
��0��ڋ��R\E��ܞ�h��y;/yZ��X�N��L蜤=����.�8�FJe��d~�}��&H����7ZGϏ��/��uX������v�&f���Qwn)�^0��w������	5�5�4ٱ������vV����^M��1rظ!gQ2ć�A��h�d��'��d��r@��W�����V7�i��c�(�,������橷��j�x�<�a��_t�E	���>�&�82���ܚ��R.+̳��8Vɾ��?IH�^_X���Ą��]��;��V�%4�4'��٥�S����d���
��I	Y���(2t�� �Y���A:sp8[��?N�zs2��/�E?l�Q��srS���?@JϢH���S���pC�U�36�e�����I��%��+j�XJ>�)C�5!Y����}SQ��nA��s��T��L=��`�3����1^��A��)���-}��"Y
����b����Z�nz�+k�DB:#v	ݓ����r)��P�����0��.Hc�Yu���S>4�W��5�$$�;i�J�Y���ß�&1'��B�Z6M��T��?Q�Z	��yE��0Mk��4l��=�V�ߎZ�з�cu�-�3�HbC3����ihB���d&���	�(��w�g����,�?�O> �v�E1(�#q������R��J�?!-X�Ǻ�o �l7߶U��=�H��]�ϛީ���2yP3@p����:z���Yч"�@̬Pz����|I9P��bvFԢL���c�H]�)M�Uq���_��y`��.�i�#]^X�[�*��V��eh�BEn��[!���SY5~�j\	�v���.l�,Mk��>_F�ګ��8�<���8� R<e���bC5@�t��ň����|xa�CdS'��-��5���q�Z�x�=��u�w�#F#�w�fp��ߢ0��i�z���f��]Z~�s{p�e��pou����F"8��CT[�5�����'=��WJ�9�*��h�l�~��BD��G/����-ŝ��D��=jX_iD)��;SW�bt%��2�l�.�_�"S���c4�uJ������إ��v�Ć2�lW���1.L>L�:�l̪P�%����@�/�US/A�1�%0D���	Ks�^����AI/#��U.r��v�=�N�����>�Q	��k��4L��-�w9q���9QfŇcg[no�Έ������U&�rm�lə���9y ؇j4��(�oY���Q�y��kŌp�+���B{�����C��q �� .�K�"����6*I�Z����[�ka�W�^��W��7E_��r����?�m���|y���8�>����no��O�%?#�l�u����6!?�k���!��[�e���438��Y(+]Q�9ñ~C=�௜�#.��p�o�/Y`�3��4z����,�o��nBT���4֙���?��B�Oa	�2T�pL���Q�F��~x���凜�+���&�'@��-�I�D®I�B�I�D���Iq���X��@zy6�G�W2L�~x�V$8'�v�?�쐪XB�#|��︧��KB�OI5�0(96P�ϼ0�c�3{��rj��<Ve���!S�RW���;|�&{�, ������@Sr�)��[(2o��&��w��_BdzH���k�j*2^	
n����?�A���	�������7{_�O(����k��J�@]g�����I|�� 4�u6����'�D��G~u�.�L`���3=�>>����r[pH���5�&�X3�ծ�=��A=p?yza����g��ח\��b�kw�}"ל�<ɞ��aMK���o0N��ϣ�.M��������#�.D�i��r��	���{�\�������゘ݯlx&��	���D����Ͳ�s3��T���EF��	W<�e���#5����c��[|��+߹[���#%Rm'y� ��I�ci�s����b|ܽո�5N1�*v��i��p4�������ƌp`�wyʹ+��ʒ���'4��۩���m*�+S�C�$��b�B�k�}��3Ơ���S��ϙ����N\)Jq���.�^�`$��Lwx^�_tŪ,����TJ�&˖�G��G��C������v����#����դ�-��kQ�ךy�A�$��N���N>�\���gwQ�&��k�8@W+�ػl�'�X��	��Kb;^oL��͹8eo�ocg:��c�ϑI��
d>�8hRDH;���$��{�o��9�<��Ta��p�)����������1�k�k��U�	!0�H�3 �3L�&��#�F�3o|���'���W����,.0bK���ҡ�OO\}#��F޷���,҇���F�Q���j����9�����eM���=�{;w�+b�;F�ht��&��
D�<�'N�e��j^Vk��ؿ�lw���q[*���.L8�[��]/t�-}��Sl`C�U�Sz̡7���<�;��O>nJmc��	���
ϳ	�&�T��2f�JH^=��w��:bj��V�����[ɌC�����Lk ��~�.1.�r�h�G#�Cg�	12|/�@�� )ة�]U��'s���>���y%V0mrm`އ��	�	��M7�6��u ��R�r������}�⯍�1�<�	 b�f��Ŕ�����P�Q�-vr��iذ
�d5�nɏvb��^2���Q���''Zہ;-���OO7t����@=�q��t(W�;�j�����	�� a�phDHEjl��"��_�G���;�!�ҊnzAh���@
�<iH"����Mn���s綌�B�?�R�э�$��=)�r�/�㙮��;¸x�e�[]c�D"��4����Pթ�}J�'�qYN,���$fߣJмD$�r�%JӶi���zH%�ē�$�e�к(JW�ݩ��(?�Z[�P��R���y�$�f��3��a[�?��_ŵ�)[����ET�����_���\�C���
H_Ie��ֿa�Ji�����D6��I�mQ�m���rgM�=�)���	/6?ӄS8$ES��U�V�D�Ub���V&n�p1.�wxaP�+��,s�$��o^k��hBf/��"����M���!�5��O�l��	�j-���C�bҾȪ�s#���S�~��j��I��_8��uXPζpDYG��!�RFvKO���B�S��P�)�=Ձ��(Jиm'���iC9z��W�!V�vR^h91�zC�A��Vvj�V��/�7�!5������?��Y`Ʊ�3�\@�u霠(n��	�%�05?mǒm�w���|HF凭��i�m��Hu����2���{m�i!m�R����Ũ/ %a/@�G����A�T@��c����/��:��5ޗ��v�5���䝯�\^k��CWG\-�u6����7Q:B$E�x��,s�6��Gו�J�9zwX$$�A�ɥ��>��W]p��)��Q�)i%Qض��GG@paA��u�q�P�'��%`�9ٯTń���%�P��!�ݠ�(�~h7�
��SY8�,��}.��Y�e\-��{���M!8yb.��uƈ�p�z=@�Y��f,�R�&d@�A�E������v ~������)�u��+t���R��.9���+�$�M|j���-���`��a������k%t��;��Z*�8��5B)|Uh��ӕ�xM��?�(��aM$u6�����*�C��6�'�V�E�a�<�`�R�E�X�D���?!����R�[��b㎤ܔ�I��]3<�y������8�(�����大��c߂��il'M>��S�����5H�t�%��Cg���P��#����e.�\mJƏe��]&�gF�$4��Q���O�(�`����*h5ص �gt�Yr��X��XvnEk�rz�yW�\�P�/�G^��#���1�Y����N��;�OG2hUǬ��i�Ձ+��E�۟��]�`�R}��9�sgL�//�>.'��*ċG�1S�T�<5���F-�C^'��oF֧u�1ǥ��"L,���u�|H5sNI��� ]���P�<8=��<��ŗV�,3>���~�_
���{�!�g�)�ݬ�БIRLI��U�pĆ���@�鵯���Za��X'NǥUJ����O�]�r��Ai�2>��s�WJ*O��=v��0�oF����\�F!~�E�-�5I��*��ֿ�nK;vn�{�G�����[����*c�̢��|�ΰ�)R�[9 ��)z��|�k�a�Uy��.g{�;l�`>�T��vM����4z߿�g�/���7&%���r�_��U����M��c_p�E�Ǵ�I&���G�Im�WmϹ�b*&�	�P��Wʤ�'8u��
2@K?���]׃Uޢ�2+��q���2�k�!=a,��F���ut��OIvH>(����}�Nd���~&���I�Ęs�e��4�u��m�Y
mZ�}(n���)ީ�	�A���0ԯ�H0ZNUj��P[�V��ǣmd�:&ݡgC@�l��(�?�UT��[/���2GH��3/6���&�����;O�p��
�y���/2�싚CZ3s�u�M�?�d%�t�8��O��Mw�m�%��t|�,R?��FIA�8��_9�����dJ���a�v[#x��Ώ�u�*���U�9���I	x!	�f�ʩ�z�h�'��.���Hwr��� iD�<=����?��J9�i�����t]U��S�� UK�K��T件R8TE2O~�'�3
r��I���>$�V'��^;1!C�EY�Ƶj��c�ڽo��%��S�RhF�*e��t�Ŋ�����A�W��`�A���!���5���:+��h�~�!����ۛ~�Q���� �c)�`���3Č�S���_Ҍ�
���µҖE��e3(����^�6A��s��7�-�~z�B�W8^MLѻ�R*5y�07'#���s�*�9d��Aa���E�����U�xs��&�3�`�WE�����B<����]� �=��SE*.��K%��?��0GV���XmS�♪��%���
w瞉�AT������� �<�V�}VN��bDm��l�F۬8�����S5֛��7��T*qC����+��n�5
_X�^��f�&"=ҩ!P���gG����jl����M��c��a^�j���}s�sf-���l��̽��w� I�7rM���^m�/���x��#!�t���:�ˌ�Zǚw�xy�7��K�UnI����~��� 0�0�|/N��\e�vE�θ�-�:�)L�K���z4�=�5J�d��n�FxN��T�x!E��H��7ܟk��	���K�߰G�d�D
�;҇���⟥�aV�!��>�PJ@�����]=_Fy�vC�eD�.�5�,��DKq��GG�m��aQ�MR;#bfY��s"̳��=�b||�<�{'A�g�;*Kr+;ZR&>9lZ�
�Z�b�%:d�-=������c`"�,�{@9�:���1{��_�{P\{D2��2����ۂh+6PvI
�$YB�8��:��T�/�p�/�l2��A#��������.���-��c��^�E�}{���m]'k45�!fS2�О(���9���t��M�	&�ӊ� X:��%��<w�Z��*�JYJIL��rg ���Coŋ鲔��o
f����Dkld���Ҫyo�~JW��1[Y�[x?MêOl�oG���T�%��f�JUTP;��L >`�~����&R:�X ��~p����ǕeT&B��g�ѯ�ҫ	Ĳ�B��bB�b�xlNE9��pEͽ���eW��B�$�a\&X��휂��t~�^��uGBأ���'�M����_·�;���D�G�g�\i�\,��,h���*�1۵\LqW�ٷbn�z��3ԋ1�t�o��Jg�Pn���pŀ�A_J��1�.�q�}�$z�]k����ɧ�Z��!�`�$�1&͚�O�Q@���ƫ��I�+7��cvߤ�g��S�
�/�ye=�$��7wa�$!�UU)�?��[��j�_z��b=��\2�<�����MϺ�ӥM,�dO�x���x~�ʞa�N���=���L�ƝY��TU�#>Z��ä�\���;l����3������_�U������uZ���Zy@��w˅ǿ=�M+!\��O}FV?���[��k<����Ja:�p�����0�� ~Wt�{v#������l��&X���,�x�<�7��B89�Dm_�Y�$���k��'Ĳ��<�'6H������Ǡ���{��z;s�´�ρ~*΄]���O�isc��?�׺��A��A���	�e���ۓ-Ҷ�}}�Ž_��=��j(�AK-ܹO��?�=Yٿj!'��n7�>'E��6�e�!B%�V�B>[�:���������J���20cX+�>���hpXE��k('��!f���a6�m?��U�U�M�ww��W����C�G@�k�Rhɘ��T��-�ac-`e�-f$���-�4��)���FM�/V�!�g��"M���1��K���6f��L��ƾ���BWڛuA0��5��mqjy�;у�>��7�������TWryգؗ�|oA'�d�9�["ԟڱ�sс���)���1�B:�%D0	�㠈���� �tL�̒n�P>7'@O�<s|����чo��~t0P���-`
#�'ۭ乲)8?��^�<����������_�y��o.3u7=%��7��أ:`��X������L�d��lS�;j,K�ʴ+bZI$��>�3�p������]�����9;۫�ù$�`z�k���O?<[c͐S�1���<MQ�}gH�Np��m�/��CV-�ח��?U6��,����Zx�縿��F�uk1� �\>�u$l*e���pC�=�=�2|tv�e��7zn�;�L:�g�2��S޻�``��V�WNY��$ޘ���V����j��(���6d%�ك��:I`kx�EL�ڸ/ȈF�������X�gF�KU�1��SE�t��z��b�bg39T^9����&&����G"� =�xc-d�2qrz�ӳ�[GG�}~��ȭPU��7�T�䅒q����bJ��8�?�in�C�W�p����u�,�/"���g0D�
�2�9�D�b�~R6�#L- |7�����c�Ym�l8h���x�tm�*QL_�M�u�M�)["����VIwğ����N슓�b����&��'�)p�ld���Nd�J�^������#�Y��<��7���
6�+G_0g��t�I4	g�홁F�'#�2�2T:Л�k���G��v#!Zd�+Χ�_Ґ �oc[�GМ'��g��_���z$��E��L�F��`��i�.�!�c��%����g�O0���k��f<�b�\��X�ڗϸ�)�I��BE���Ō�(%��й���7-�Qv�]��M7;��Bަ���{�"�$-��&�}���˫+y����$<�:%_��
�zξt�:��<��,5~Y�����+3>��1�J$T�6 ���m¨�>�J&x��y@Ȥq�haQڎR}��я�;��{�g�������"�i7B����`O���z��mp��TKl#��vO9)�ʿQ�w2�#ya"wC����D�
TI
pQ>x���-XV�=��!��x��R��j/�H,�U=�2B�e��v]n���K9�yrLƠ0�9�E`q�Pǿ����AZn&KX;��?��˦3�?��\�5R[�OeMe���øH4��/�=@1ܚ X�,�y�]�~�5�T����2!qG�xx	v$���ڒ_z2���^ϰ�=���v�Xۓ�����R�Z�e#�*͊���*�����w�>��(DpBB@y���g�3�Y��^�t�X0���)7W��v;�%���e��h�BIr=�����KH�$��_�݉.��ˈ�������O-{R~��y��5Et�푗lG�K���o?��-ɀDd�Łl�]� ��	�l���X7��5����jZ*�N�GϤ�9�/O7ς��P\ݿ: .[�����Bq	D�d�`x����u�������p	v��"�?g[�͇�3YHh&���ښ��P�:,8����*��$���OD�g�Y�|������r�NBU���޿����(�rC��{���S)�ܝ��l�����C��Ś��i��zk*�<C/�&��$�z�r�Th��E��W>��V^�r�;z+�޷h��`� �%L�ZL���|�ߡI�B++�Y���Վ�,BwJ���x`���XI��c��0a6};#�Ժ�)��Xt��'��9��c =S�{1׷8��m�@)����X�i��c� /���)*�n��ZM{�Wd�iI{\6¡�n�����@�=3G2S�A��_O?�ș�O�s�f��".�K�]�Kٴ�R����)<�~�VK��.�U�h?ݾ��j"��%���â��YV.��j �%��d�����Z2��'f-�7�� ;�/��RRd۽�+`_�d�"��O_��A۵�]��|��e:̂�f�sᴚ�
���&8LϠu��+��ו�����[��`"�����U�p��-v����Т]����۫�0��ţ�K��\$��L8x�o?xeY靟I���H�-y��1�7���ˏy0����X�,�[cC#��O������*Y�^�V�L��I[�J�d���i�vEl	�)k>3���f]K_7���Ȳ&d�1��� ����=��\؋\���|���$�y���K����4Ǣ�x�B�:�G�z�A��A���H�������>�Wf���*d&����}�z�杯���q|2���d�-IWQ�vU������W�b��J�,`S�*Yf�d��M7�h#�y�6�/��J[e։i�9</�1*9��*)ED��H(���P�UBa��VTUT��{��n8���ԘIQk��&���VC�O��;���߲� ���RNFI��FLm���0����jw�{����*���5X������(��^�i6�d-v)	���Ӧ���e���2�r��$)|�����5�_�q �4�hZJ��u��.f�&}��"O��m�
�� k�`u���T����F�"YcJ;�&_v�I/u?CTs�Y2Ӹ�㾬�q/˅p�`��Z@eD���Z��.���/a
w�*�n"�d�}���"Ms�9�kk��L��2'r�M殕���#�ᇶ�t�?F�g���)eU���*!��3,��cL����X	KY��!Іs�*������C����֔��Ѽ¶��5�s�%��T�"ՙdZ�oq(C�c�y��X,�壙7h��<x�WJx��R��MyY�+^��Y,��H!�����S1u\(�4*o�t�f�Z�	K�[ˌn����L�Y���Ng?����"����5"M�x��%9�8�N�����I���gZj�f6R�tE��f΅~e�y���	L!qЕA�r,��㫘�2�Ҷ(H!G�y�����E�VzlQL�i��?=�g�66���HJ9X-��d�+���Q&,����|��&H�����(&3�5��df�ݷI�%Ϭ��bA{�ï�^�)\�S�=��3����ѪI�hH�e����凿�*`Y#��'�:�\�R�u��N%=Ѿ.��W�0�L	T���D��P%m(��N�C�(0����s)=b�7$*)��g�c+�^�v
��Bh6�����$�?����X�s�p��ꪓ�r�cś�k�tշ�������gi�A��/ro&6Ȣ�����j��;�[�����`mx��1[�b��D�B�����-��&V�S�G�{��
9$�#J���?.5��w\8֮H�^.��m�%�)�,+c>���W�kf�f�m�3��4�R9y=(�y1%����m�y��k:-R���2�]Q���l[�*�*�r�T�Ϻ(�����ܠ>GP�K`���O�|
w9��E�ў��*�E�M�����US��fT���o�0�rm	l��jzR^F3���c�����_I��B�]���5G�4�Rpq��|�.y-�#�h!��ṳ7���Lf�k�p�ρ;�+b�������������8D���ڕ2{��e��ۓ�x���:�mֿ�"!�� ��1����mc�,��;|�Rd}N�)+��C	>$	3�t�|��MD�̶�]��Ă��"�`;Sf;R�u��%��<��cm|a����x�	aݮ'a���9&�SJyf�ڪ��ʯ��q ��4�k��}ה��x5;���r�U�}��1�h�Lx|���H+Jt���h��w6��AH������s�|4}w`�h����|v�q,��hY�q�P{2�HYe&w��~9U�0�L64 �Y��/@�؄���S�"���H��j����"ԉ?��vIw�Oj�!��9��,�M֣�\�\ץ3�m�kb���)R4��Nd�z�Y�Wju����5)��C��m�8{Cw�5�xSl�r
_3�KP��D���qH���XƆًu�q�¥fQǕ$�����������t���g,���^���/O��}�`u=$nb?&�V��<���WnG*�vW�mMCav^6H�*�ƒ��%��C��k���=�\�@��Bs�eQ����V��9x�#Yٟ��m��9�DHPv_m��߱N��51�'�,��CP���$�>��C����Ur���ݎ]���Ӷ��K��[�:q�:}UA!�Θ��h,����'7��4se�I/d��x.!��[��#�SR���l�rGR6�:���_��⼒nt�3-�-��z�'(2���5�O�獏��h_]�^!��*�1�������:�����;�sn#��/$v7���2�Q��h͛��}�du�����WY��w�p���	j�nB����-�ȵ���?謨��G��bn��i�-U��o���إ�iK�Gj�{	�4TD�1X�w6`2T��1'tO��Vx�ȘZ����1ĺ�L?�1,���
��鳷WN?��t������R�+,IYZ6�� %ˡ�ǾPj�v�:�Ǚ.sd���~W��pޤ��g��I��g���J�u,�!a�qB��I����l%�8G��{�����.��k*��$n4�7'�V\�M��B�P���2P�
�=�S��֧@*띘�޻���-��$��.O��ץ<�;��VUS�	����3��"�Pg������5�^r`���F��y�����>牣��4:��]�Y�Y���S�\롪��I��"U��F!攴6�9,��T�����0�����{J}NO!�'c7O��f�Ի\Q^��Ԉ%K���{��6�?�~f�wR8U��xv��1�s1��H*�[6T�H��B�Ew�A��㐳�������i`�>��3f��%�ȁ�;L�wM>����������l�k�����2��"�Z�𿑑TW��PK   AaXU4Y�- *- /   images/9c0c4208-33ce-4eb7-a42e-8f166060eedf.png���se��=|c��ļ���m۶mMl��ę��ę��'ϼ_�ϟ�����:����ku�>�J
RH���   I���
  ��o=�B�{�ef����]� @��K�G&  ����EԼr/{`r)�����Wf��2�s!؆��)2�՟�֯s����w7�H��AБS�h@eOY�z����VW��3?ܘ��^��?m!{^�>���?�DT�d��d��Kb(��Y��q�7H8w0rx�%��O�1zxX���ac��!���"���`"|ڲ����FW�N��}�"%%��I�q���٨�����7�"�{�v�\jki��y���r�B�ۅ�����1�?�y��|2���@���W��okbB�4���lbϥ3���$q�M_��j
x;-�5dƙcވ�`�߮�ǼM�%�+A�.6 Z������W�E��_�/cB׿��u�]�&�}A�Hc&MR������EYf�̫N���r׀���.��l(���\���_���A!swk��=fffp���� &����6�?�#X���Ǵ���?D�]2T)�7zL���Fp���=���dUE�V�%vK##��U=�)���t�f���U�M�U}O�ҋ����g'�!��eb���HǍ����8)�By�~+��vd�^��ټ��
m(̕���_]s�I�K-X�>�yy0�>#��e2�-N� 7� ��nZ�	�V����%���wL�[�Qc` ��7�� gМ+�0�
�A2zQ�k�-�Q��������y��vvuՃH\��� �Z�;���$r��I�"��F�� �9�9���	���\�@	���TU� "!����FØp&L[��{�-�����p�k�ޑ�D2�,;�(�^!Py@��x_0�f�D�lF�!D �*����UǜF�ljB�q�rR'F�,�����'��|?�V�^CI>
݌��wz�ǚ�AM��WB_�s�F��A�{F}b�������^�H;�Z�!�C��F�D�A��-_|;�
h���	J�9HәP��Kwq�=�|S^
T���ڽ\P�n�qT��#AFcZC�����Ƀr�Q`|~�9?��ɬ4V�P]Er4�QY@%`D��cp]p�����;cFu�b�a?z�zBK*8 P���i��޾n��"�m���lo0��m�k��;7]z`�vd�����ϯd���-&V$̉��*�����Hi:4r��O ;@�	H��՞"�ځG���M�ݖ�^�v2� �Uns_���� ����B�= ��ω98

>�*n��tWy�
kAH	��ދ�R2�w���Ǯ� �j�AG5a�eJ��~�y��.ժc~�����-�V�|F6�v�x���A�߿��5���Θ����%}�f�Ѡ� ��LǊ�"��rb���8}t�Y���K��ܸq\��q3@ll�
|R�Q\k�k^�(l�<r
����z$G�%6䨒�\?D�PHf�΅���iC�i�B�w�ڜ4��߯��f�Ģ�x��#��UP&|��$�D
�l����1�h����[S
��g\}�OZ4�)&8^;�E�A7|�� ������t���z�f��Aϛb67�__i���Đ='��CĄ#� �0q���4�#����Â�{�&�o��4�¶�wN�
Ԣ��uͽHx�)��J�����pv ��_I�bWU\z*l���E���ǯ��';A+D�;�o ^,�H�8��`��~�O�p���Ɨsƍ����쓭+�ۡ�# J^lս����gx�zv7�C�X����h��&���3���c�0�\���o�"S�P��'4(����k�M��A.�C�2r|�d��v
�x���<��vy?+�`�Wo?�C�@#�,��ԍ?���f�dQ���"�-������ѰE�i�����r�N��swf�v1?V�a�o��E���/�Y����();6oƒ�ą����G����Y6_p(��{ "��;�z�Ad�D��+���.��8�n��8�n����Lrߐ &'�c%E���y�����Kr,&��rizK�3�ZH�1�]`�(q�k||9�S{ L�0t�
�L�B�D��b�a������W=����$�Xw�~�8w�t���zWC��.�.��y_b>;�j��Ǌ��;�+*��L_pf��3f(��N���-,��Z�~n��w�!��BW�ų�;��᡽ރՇ@(��'� �TepW�������Q�ym x�X�<m�X�RH�=M~�7�H�� z�m6O�X�;*�3��W�p>�_����x/��= ��)
���"e#�47ze�kĖ��zR�Ń)����C��~�o�x��ͼ��q�KO��z�8�z�/~�(2;��(�7����)�2u�%c��Q���F1���"_r�.P9 >��*m���:�����Ll�lD�1�o>�Ńh��"��'�`	2�RE�ߝsX8�r���"����2�&ޛH]Ș�����O��w�X��CuΩ{gz����ZH��M�&_�z��V�8��ޛ2�_��.�3�}O��N8�fh��HC�[��D�6g� �rE��^�|aX2�"<	��c�6Y��la��[��Ga�
�,�`�������T����Kl��e�Vƨ�B=����u�-H�C��O���
,����%����_�{tM�s�C6��H3�ꯏK1C�4� ���ɇ-&��;]�����V`�r|c�t�2�=���4��X|,d����P����M,�߾�$&��	Ȗ���9�O�W���i͏��,��f}�O�H�QdB��^�G��Uoӽ5�ި�3�	P�bM��И�$sC��"ī��gM�c��Cl�-"�v+Ω�]<��}m/1f���IC�8H�]S_��S����G���}�xc��J�ȭlOG}|�sJ�T���dLe���AH�= ��Ɨ�z��J���^��gls��t�-U;�Q�x�Y�'\�&��b-�l-pb6Vsc��o�������~�0� �$�W��?9�e�zfm�h:*w{k+�G�o�"$ΏѭE��_8��H�~�G�e�{�5�98��� ����[�m���"<K-8�����cB�W5���8��������y��醐8��O:$����r�i.����Pȓ7vȕ�NP�gY�.�t�p$I������yX;�|>����l�0[
BI��.~ˍ$���"��Ϗ?���ă�^�ό�݀'_��`���B/i�r���ߘz�u͌��c���!�Vu��h���)a�AC!��=�����e�ur�[;$�{�y�O桢�����٫�H�r{}\��p������u���}���4_}H��uTϼև�Y���x}���N[�pZbF&Q`[)�>��z(I���f�$����G��(h�Ȏ�##.6����gE�B%��!�
t�B+n7�!���Bo��Ċ
#���}{ �
��M<rq�So
��{�k���ޱp��D��c(��Qd�ӏ;Q'f)��dk�A�,�B�X��T{�~>#��̝���K��C�������o���Ùh^���{��e�������'R��q
/��4�8��O��Kbw�8�_�sv�`��!����2w����'(�_qa����Z�Nlp�L�ܿ���|�B��_m�Ñ�͔���
S@p����F����j�%�t3%�9C����O���6�T�K�b4�C���H���u��ALkB=g�?�������d�*��rS�)Л^�6T�(@��Ap�T������Y�B̔�pڍ=4Q���@�i7��v�a%H���g\^a����Á,���'ǃR��B���ss�߂���|�v��x~H�\�+�����w]R�f��=:lr���(�́D��+�zs�7��h�BWv�K����8zx��D�E�A��[��z��/�#�爤���mmm.>�}����	}</��9�f�N�����R*S�\�� dx�n�2t-���ґ�W&��e*~�U/N���5A�)������w��`ZxkM|B�N���B���ˋ3��؈��=lS�Ʀ��A\����=��^i�(�����<ղ��)�6���-����5=0��D����O���u���D��c�ȋ�,��[pɄ�|��lb���C-�+���뷟�H��6b���������r~���6��g�:�T�mu|N�"a�o��FFwc!V�a��zjV��]a �M��s9�ջ�^��~w�A�%`�a ��}卑�}�'k�귝������c�����I	�3X���R�������jEᛗ�k�VP^�K'���c��3�HV��=	[УoS �H"Fѣ�Qt�o�������B�}Sx��+��g��%��5��N�K���I���o�1~l���g��X~n�^w�[$o�Evb�Bc��& �,����:��}���P*��ӇcB�C���4C-OnY�1�wg�&��� ��p�=����n�y�l����[��o],:
N܂?|������lmM����a�
���ķ�^�m����1����Iꧼ�n�4�?���J��.>[��>��� {^`FV�FAW�B�"���	q�x�lh�`�:��O �,,"�wIkv�I��w���*�"R��s:��Z�&-���8�hW%��� x@��H��$�fYʴ���_
2}՚�l�����X�L�E�=�����M8�E/%W��2�|�s��&;���%7�3�LQ5G<vĐ1C�c��'���'�,�
����ȩ��_�a[�j-��Zt�H,�%Q�e�0$u:,VƔ�����*�&�����8���;�;/~�6���k���ݏ���0�ذ���ɕL���ӣ�`7U����!�P�ѩ�\��bZS&�����`g�;�X�5(3�a����CߖƢ-����1���T�ӹV��C<�(��'�
\-l���m�NΪw��I-;�v+K�	'^z��Q&F������g[XU/)}�mglo�Wa���>dw*���I���	^�4�1��3\����L��@c��!5��� b�|�>�D���)�n�n�Ƹ�WҨ���<]3Nf)Z�%x���j��'
v�={�j��y�\�r�|�,�o�BK����-āf�]uެb�qq�	C��6B��T�������I*�85x:5ܴ@H���:,cqSS��&�p�Û2;���Td�I�x@�6&}�i5/���9#����=cb���s�z�4����Ļibc3p':���O0Ƣ"�wd�C��@�sk�JF���[I^�\��^�>"��.Eqz��/�jQ�O�!֤E���"����0ho��6'Qrh�p�?�n�L�<�W^�;�q"��N�x���_��5:�bA��A����K�y��Uae�5�#��e���z�O0ዑ�b�N��՚L��<��iґ3�R�d��k��9�>�r��P�?�h��LƗ��[�+)��_�۱N�:�Y�d׬ܐ*�E�Ҡi��ӓ�?3R�Ad�S�
)1~�	Q��R�<��n�
/;s<<"2Rj����Os�j��7��2?�p��^�w�DB|��#*ɒ�J�/1�����|0~�Y���^�����vmRd���2��_iECu"�ę���;����]f�\��B���g?�IM���L��no�8�V�/7ԯ�~X`:-U]�/�,�	Bχ)YO�y�MD���o�\=ކ����=�D�{���e����Ԡk�,>ǀeָ=+=����ռ�c���O/ٰ)��"���O�����%��N����3$G:9�C��Bn��&���	��}��W=���ؒn���O܄�?8=��b�����l�ȉ�
����i�2)�w��K�qzP�o��c���z��˕c$5��	IQ=h-�5����O �7ZM|;8���ȅ��q��J���E���蟝�@K�`_`kw|�N�;�,E�����֮Q�/���i%%Jp���]&Sǖ?�^�U�S@��8F-�k��"K�M���z���a��[���B^z��j�&�Ӥ�p�U/��hkE��ڻ7�Z��IU�Z�P�J����emdu�7�=Ό��;�Ȏ�07\�`�~xv<}�3+Z�-�Q5aHn=�r�R=ޭSc�n���r�'pe1�;C=��b[]o�-��ߏm�p[�j[�4�ص��ԩ��JSU�F�_��)%�Z�R.>Z�&wf��Ο�2y-1�Q|�􂬬�2e������"���ѧ�l�+�'=��I�C2/�:j��Wl{�B�oxY��$��h�M۪�D9l^�z4+JtF��%�N��o�e�J��5��M�W�rK��c
|n.�93�2�saoY5|�;�a�;����k:~����|��C��'��:y��Qį���1As��gj1aڞ3�v0��h�x~��_���4�z��M*�ؚ=9h��.�*�������Q���b߿*���r�=���e�/��O1���牰gLAo��呙`�>B�׼���u��C#.z!�n��jJB�Ō���:�5��̤��~$�*��u֨�*�^l	/�K�)OSm��{AϡX��j�7�X_]T��8�ά��6ىf1j�D���h"m��M<O��n�Ð�Z����N��]6F�A���̂��YYN^���]R�M�8\��=;�N��E�ԧD&�:D�B��X]��b�+��/����1HK�MEIn�3
��tG�1��˄�H�Uf�VZwE��a*�KQA�#iU.v�fm�l{�#���J�i�?��M(s�u�ؽ��8�[v���`G�&2OF�}�V=س�H��t+r��`���p�>r�SmMV�;�ͱ�Ϝ0�8���U+�3A��4eIn�x�ϫd����W'��'�$&n���o5�-_��i���$��2�*&CH��!d�b��J{��8V�ō���nV���H}y5EA�Wh�Ȕ&��uA�mZ�G~Ű�<Ge��wF�?�Tx�����F�����-=�B\ݠKq"�Sb��]�:�y�$7���e�4�2��"��uU"�iJW�!m���(�!G��?Q?�ěD��9]��H�5�]S��#�i�������(�"C2�X�2�r)~�H��<_���N��<���c֯���t�<���3���$��e�`uz�٩�@��&����Ǔ��	8,e9��e� ���x��
�u��
G'�t�Ɠ���k��+u2��2e�v���ȏR4&q�9�꽙�� �]Z�x�cF���Ƚ�)��9Q���E�ö	�߆x��K�7�!O��;a�-����p˽ijnN)N��<BM�l�l�tWxKiK���\<�D�������7����g��w"$��\ub��&A��C{�C~r�ƹ��(�
�m�NF�7���Ż��j�f��_�G�T4��J�R������|K��-/lˊ�3^��t�w�e�'�1����Ju|���W=��պ�.�t|f��ɻ-�����O"����=�
����)KWČ#�,g��O�ڪ�rҍ�o�7�O~�ڐţ���I��+�)wr����^]�� p�6s�Կah�"%2r�%����'h݉/֦�gC�kX���wt1�����L���#��Ea�.5�=�/�děStGJ��L�)��DxJ ���܃�Pދ$�T9��+w���Gb��~v�N/�Q������w�'.�s����)�E��g ��H�ɝM��>�
��I���1g򱫏:��u��;�g�˥4l�o�xV ��ez5V|��J�W�d+����*n�A'�h�����]�3h����� ��ȧs�X:������&}�	k�Vi�i�o�9ik#��n�	x�G}��,iK_�${c�"�Jϒ[��խ"���
�������3��=�.T�
m���~��7��'�d��9���;a!J(�zՠ)��A`��}%��\��Y��\Ĉ��8��?G��x$V+���?y2˕+x!�;�E�W_ ��֜!%%Q� 	l�y�Q�q�W�/�.t!�YTU߽��;#a��[�
��'�t8�"�%��A��Ch��O����Uɗ��U�~�_��3"^,C��x0��Nxm��#M5N��J����L��-��y�׼2��Q�j�����db�:~�'�^�J_��(��۶��!�D�$Ymu�&@0�L�<�ӳ�^2�u����y�\P�r1�;�x�%������F���i��{��v.�a8S����Ͽ{PPH�8���gl�X��z[^�vq3���l�T�!�Ye����,�C7���g�M��9�F$P�Ώc	�,�Sረ�Xz�9�`�=�N����M�v�H�N�0+4Q2H���!Z%܃l�%�F1�:�D�+F,�N�,$m���G}��C��'��~`|FGN#sR�#�)�9d�����\�V?�(d�_@�M;r$ؘndE>��W:�V~��)Q�+� �L���O�m����L�Lơ��0IJ$\�F��&Ğ�.��=�	���i�ӱ������W�Ю�@K㑋7�rznz�{�d�^X�	~�KZ���3Rh<�}2�յ�v{�۸�Y���w��s�N�Z���@�p����7�o�K��C����kk�W����Ҵ%_\�~Ӏ�_�9��C��?}���;�)��+�.Eп����*���G�k$4�p0��3���{#P$��x��i�;-5L���ǒ+�A�z"�l��o�����:X�k�M��U!W��V;ٸ�V�R#D�$u�:w#<����������}�O%!e�J���)M�k�555��/Cu(�8����\Ē�S���g�ҩ1�����5>C�����v�����#�����q�_\�p��h?�f��S Q�݅���b�n�]D�%���
i(���5Ch�E��-
���ȶ��W3Z��-]��^�V��2�6�ڶ:����8_:�qV�����u��~:��6@��뵐�����0��9��em^/�'%f�ƥ;�qN���NԦ0sӥ瞡��"H�o�O�E����A� �L��BV�=T�g�;��G�q(�^������rѣ!��wh�4:�������à1�Hbƞ�ZZ����{�_ׇH�� �$�~5@��)
���j�\�D�׫晳��o)6S�V�T�r�co����;N�KKk������"$�M�.��aE�@�q�`RR�H	�i߃L�xAf�S��p@�p�DϨ��ϯ1��:
���G�4����w���UG�M��:�|�9C�r�t�ë�Fƻ�"�탢�OH�m�8gqO1�kGR�����b�nh����Z��N3t����疒#�����a���Q�� �4�LĠ&����_����j���'t��l�����:��L1��wК��Ѱ�YXtXwu��(I�L����I�k����`��%��1�_�HH�Ғ� �E�fu#X�A��>3��3��UN�B�K�/���%L|�C�L�ߋ�-r����z6<��� ݗ	='�������K&��%�R�(�$i��Q�p��!!���^	�y���V�T�-[fL3[�-��'���a���d�֯�G�[fy�ߪaH�-�Q�/�G�p�ܨ�b�$	�8�z����?G�v>���3U �I�o��9ܚz�']��w�Wxd9�.h�b��4:���g�\��X���7���W�f�m%.��Z���Y
Y[̪ ����N�뙵���t"p��A_�s��`ݍҷ�O*�l"h����ˬ�`9SO���6�.X�>��i!��4(�Y�,���&��^
�ϝ܇o�<�1��ܜ|���z��9p\a�r���rvƕL�Bq5�U2�~2i���Fؐ9�Cg�=Hꇘ�=�4(O.CDa]:����-	�qa��#�N���0G�q���:�*�y`lQ�?��Z�d��_��#4�2���8��8	(����S�h��3F���ˢ�R��a$~0'�P��0����{�JS���g�i�+��j��N�^c�A}5(7��/�#��Rc���VP�d��
�������-P0���x6�N��'��|��QI�ũiq�f��8�j����s���v��$C�L��i���h4��e��s�§�<5�n[}2�'1��2���'i��c�*�k��f�w�1����VEn)�X͓]��xR��}G��q3�c��v��O�et�xpj�1�y��
nous�w23�%�`�c��!=6�hɮ�B�}�b��I_+��?��f�1�%-��M#�?����"c�����"������h��L��R��y}!5�j/�p�F"��gs���ҡ� �١O��c��q�Wfy~�,���_JB�`�c�ԏ-[�̘|� o-6r�DZEA�Dtґ�!���C�㸢
�&3Z� ������������89xIi�Sl_vi�uN�|������Qņ>o�̈́$Ɵ��e��̇WUON�����M ��	n�u���}�g�id��ۆ� A<\IP��!�-gϭ�4�m+/n�L�T�f>~���p�f%��@��V�;���B���9��LT��~�aV�ߋ�T��g�9��FF�`1z��2��\A�:���`��W����e1�q�\�R_n1RGny��;��i�eEE��9]����0�+F�~Ӝ�kM�|~L�vP�ohG�M���<k����F�Gk���'\��4���'i�ZAZ��6[Ŏ�]{s�7T���.2���������箽������%V���}� �j����O����qÿ��a`�0mǥ�c�� A� ����I@���� �m���Aa.ѳ���y����o�����Ĉ����^����@V�h����B��b�okDe��>G�ER��E���J� o�-���V0O�V��R��x�[l7��u7@�����
> ~�-��p�DI����.�N���v��N[�ߗ]1��q �{Uф��\-$-߮p��e~]�w�GѶ[�N�e�pv��"���b$�e������)vĨ��8��O���˲�y����2k�����Ra9�UYǖ���㕶��5�v稤M��Unr=����jm	����;�����"kX�Rz�y��O�S.xಝМ#��P���Բ\�.B ɕ���K��~�YIF n�w�@q�ckP~O�������N��1.չbs#|4:De�4,�����Cɯ��v�C�q��9�e6���K�p�0J�n-JR��`~�=��I��eIM,k<F��d6jT��,`y�л��nP��R�^���H�Ⱥ��E�����1�^J�s��G*�vANizN�0�� �K�� �X G7�1��:4:�> qtA<�A�_�Pt�rU��Kj5�E/�������3�\�lq5�M�����-,���o�w5�ɹ�������,P� hp������lS���޽������u&����Y� Z>-^5�kj����71Y�X���z�^�*����AQ&�h��-���;���V���J��Q!�؋�/ҥ=����(#�	�d��.̯�e�kE��nR�[�@���*p�l�{�Ki�"���_����P�Y��p����Np�g�v+�+Ks�0H�H���V5:ƿ�'A�YH`�6TU���IުQd��� ��H<��.Q���w{֞+�q=�߽E%����t���o���'0�2���S��G�)!��X|[��3�X��X2���Y.a��E��?HA}Z��j*a=��9z͒EUFBST�$H������j���/�(�Jՠ+i�a�B��≊���T�ƥ�1L/
v(e�{߯K�cq�\g�������6�@��A��֙@O��E K����/����c��������p}6^V��*+���W��[�R�IbEe]Y^:S�T��=,�7�O�d8���bԺ��i��1��S�k9���W�Ą8da'̴l�����϶�\y~����u�ԟM!ᾎ��ǡ�-X�8��f�2��<�~�P�L�S�	R�M����y��!��ģn�&Ǵ��_�3w�<h0��p"ʗ$������9�_���UW�z��ԟBtx^�`�����[/�0k��o��fU�����
���� ��48��mB�Hٕ�`��Y���T�h������Va�M��NTV~~?�g�h/�Ά�d�@F`���zP�wV{q6.�C�����j�<�j���\�PWa���/�WV%iS�&%agwR\K	U�p��ÿ!�L�"')�@"l�N^�V�z�6m�#���	d����5��J�FF�.F<�u:��[VƆ�Y��`�z�ɠ3�e3��|�0Un�L���^PC��*�t<fv���2
9B�k�gr8@����&k
��I_B`�F����l��������䁟�K., �ӟN��_^[#zG��$�)�Y�����"ۈ�K�v�����T�t�s�Ŗ��a�;i�c�}������_*{pa�ʊ�GX�w�JT��WI$�o�>���t�h����B=�J����ೆ`�ڽ\�Y��4���&8[�ɇp��=��L�z�J��1}��ْf��T���<���]�7@i�Uv���x�� ���,��%s#Y�mв����>���	p�w�0���mq�}>�&c	����x�h�]m$�7 .7�0L�.�G�����~��ރC�盂�}~甚�s���}������F#�<]z�o#��H�Z�v��m���~jA��ł��V���6h�\?�u�>�+P�S_���ے��`�����#~(]��WR���F��M9�Jz~E�S�u��hC1h삑��(��s*�WI���{[�	�� �(	DVz;aW��`�I�7�J�3��=�DM���\���4��ҧu�Ӫu�8�#��f�2�n���Y�5���O����[\O2��&U1��`��\��]�DŴ]�l��(g��쎁���0"ڿW��>,��6�P����)}��M�śM]&b���
mXAB��<�A�������^�Os��\"n]��CP����gV���2^�����;������߃�3�U���YC�)����qH�ͦ��0�i 4"6ի�����!���h�ilP�!�U��l�/@�t]"���)��S�=�)A��&X�/Ax#-�JtuA�����S3��C�W�p�m7X܇UPÙ�R��k.\0�@�����p��V2�$Moە�q�OI�湜K�`^6(e��BU �&m:.�Tf���r'�9��C�}Y��|�NI�?�l�j����X��	v�0�Q@m�aOn��F�8=Ɔ��VKL��ǕNK.3n�����Ԭ|8���`�Y%�d놁�y2�̇ʃ3�ߨ94b���������^\�h�-�&1�LN=�����|���'d���~�����E�{?�ν}�{*��j���cA@�. ��cR�������I�
�]���M���5cҖ0m���5�I��[XDt2@%,K���"[VM�{g�����wH�6vs%ŏ�:���8���9<�x���l�D0�Yԫ���V��&��G� �C��ޗ8�,�[�HE�E��p�>x�x���0�]?��EU���1=�Wo��eQ'ML�m�s�b�>]�Ű��c�z�)o�ր���j�'OA�A��8�� ����j�'PjR�^�+n��g�$��2���-�#�����?Q�"2YV��� #卾 �s��%�x�!��}���Q�.cdO;o�����4����e��N��3��m[
�F_�y`�$���DO��� ��}痌�}��; i]��G#c�܋psE�k=�A���,�E5e&ȲV�Nx�!�1Z��?�$.�iߑ|�V6FdɌv=v;�Ʈl���wo_�����q�iN��G�g��|�i�G#��nGD��}�$~���!�14�n��3���OG�O����SՂ7�T����>����/nF����:}ɦ���E�%�2�$�ѧ'��~�!�����K��X~C��'d�%L��wgʔ���c�䕜FH��g<�_:�������p�y�]��`��rv�>>�
����8�~s3?v���fB7w��f���*�%�{Ȣ���D����1�>r�+I/D(�v����c�W��b�ٮ�9�P���-����*���\�כ�H=��b�IgDf;��v�'��>H�{;��y�^�3���&��E��/-V�R���ї�C��E&ϔ��Y*�i�$��F�Ƿ�Ӎ2Ma'��3�<���9��b*���=`�ٌ��)�L�\��_{�Z\���xD�ڐyݼ�|�gK,�>	��W�nƕn�j����"o)��l��6
���hj��P�U���U�#� 9XDb�gJlޙ�C�An����,����W��"I����p���۸ gf�b�	�&���@�;Rg4-ز5-��xQ�%�����T8>��Փ�u�4h77��1f���~ęD���
��9�f����[R� 	�uj��?T�i콽�ԍM�{'��k��9���D�j̻�FTV^9|92�U�z%&@x���!�c���y�Y�Ɇ� DJc�ČI$���ʞ�4�����dY&4���%Y�PZP��w��:�k��綥�#�{��y�xF�.%�Ṕz����p���v����:�j�A7�k��9~:�-����qdȲ~�E�/ʼR������ߧ�;=ϛ�(|��9��ac�`���\��R�(}eI��e#�~��%�p��#�4�4lkn :^\��}9�n)p�Ҩ�A��Ե��V?�he�M!B����_��ʃ�mR]����[Eb�(Y)۩����ͺ�b/�i}�)�/Apq��_�a�\VT5���<�
_�ٵ	7��c1��<���l�k	7��>=6|�8�/_�f���vA��RLp� <��B�1��<W#т��B'��Q5���m^����Ӧ�����f�v_�nHn�yKgj牥7�A�YiQ�����CY��e߻ڃ��+�!c�z&��>"(��Y��B)�����gs~����B�,��hj�b5*YY�geg���	cW}��v���*�R�u�A%�����d
�u�X��?D��Q�T�n���w�BJ\Z����v�0\Br���R'S�������(j�
�ίy
����XH)@F���Q�So|⢧���؁�p?�v�5u�@�I_ϛ�F��ҐVD[������(+�}���E�+yS��& ��dP/����8����� �B�ïp��1�r"�EE�+���%Ų_�BOnϋ�fј�\��M���hu{Y�*^��WAj�@ݔ�N%ǽ�M��H��X��=Z��P�x�y�'�O��1-�*�1�M�(}(_3��_�h������X���i$5s}���ez'�ҝ�;9��V|ȼD<��}���0�_�����2�BpMl�b�Av)�s���k{�����j�1� Ւ��	���{?tK��7D����^fnfv&t�X%�'�V
�Hq�牆_޶�_e{M�dtٵ��J�l��L�/\�V������� ěMHR�n���Ou�y����r��PQ�6c�g��\2�t�õ
���L�(���S�t���(ȶ�iN���������1����xK�sIh�g�i�ζ�j'��.+;o~(ZlE�ny��s��J4��k�?J�
1 ���ͭ�(�Uz2~՚�������N�{�'J���_��}���վ�4�φp�y��R��X��a��8�*Ƥ��@t��m�4�_���/$��?wY��;0��p��)�8^�k��D��[&�o�u@���` ;�G�w������>����Uy&�e�&����k1����M�}6�^8�f�{%y�5��-K�x�H���D_�x<���z�!������z7�ab�����V���Q��O�Od*�R�{c����cs������y#�<���x3��-�����𹻻/��Xܐ���@������XVƹǟ_V���n1�o�9�h6�u�%ߞ�/I���٭�]L�=�ɯVg%����z7���{��IF@}/�����=����H�� �d�x?����8�r��`���(�m]nQ�#�gg�fn�4�q�����|IPQf˩D��Yj̢
)�����޹�[ �(�Ҟ�]�^�P�Ҷr �s^l�c��o��rPZ�n�c1��c��j�mgJ]�pd��O�qӊ��z^U�
C��{��8Ͷ��|V��ަ�z����f\4�� @��w�Ea<��n����!��^���O��V	�GN���� &N�J�㢝ø�9-)2*~|���z�&z�ϗ�7�^�l��O���.jc���G��u0tZ�p)��U��u�i��u��kiH���˙-A�ul�z�"��05��4 **zn
�65��4�S��$��b0��*;�C|�`p��(�]m��-`S(�jA*�u<7N�b�ś�YRL`��	#s�����a�W����`�<:眳ar�t�� ����������7���u=}����3�M�����)� ��H�CN���⇉G �x�%� VR����������7o������z�o���E0U��I���<���~@��%a�������d&J^��s$��z��htd�y�Z�p�0f��T��u��h��>Z��_���~��(���(h�/~}���З�|5-Z���q�34f&˘)��un�V�i0��v�0�K7/���w�<G��&7��qM&����A�dJS�H��I�A���lA�|��^~�#;.J/^sJ^�E�W�������ja�R�$~ϵ##c��6��]�G[h�ƒd��P���D�*���9�� �H�P=�*��u��&���<�X�T�e(�����EfϷ殇�s�s�3).Il��#6��#v��((kG{7�Æ̶�������δP6;sV�_8��>�w���І;�R�k���z7�ٻ�͎$����ڸP�����sT���P/���g^H 'm\'�:��0Y��K��~\�b˓��s�+�n3�}{�ʵ�Ǘ�41>%`��%����u���<u�w��Ç x�0a����������9mt�ͷ�$��ww�y��N�m�g��jff0E�<�3���u�
���=4���j���7�ꕫ�c�B����/����O ���K�=�v�yy۶m�2��s{hNwm{��R,;�jSG��G%$�����������o��N;fA�֮]G��Ȗ���N;�Lz��H�����=�0� �V:�y��MXLf���8��O~v��.�9{�����Бô�?��E/��?|��$ʀ��n��~}�mx�'���{��~zы_F����8������B�:�1��Dp9�i�Q-ʋ�ep)�*���*�~n��Dz|�/�+��W�����5�H֓)`À�ų�B!�X�r�S6s�u@��qB�����޶`�I5�2Z*�^i�BFn��i_�FC������'��&��'�Fiؒ��u�3B#Z�����	�9h]��R����D¿�n��v�����=K��̀��.䥡���h��d�V�
�&(9����~pC��޻��N��~����F�W��E���]G�a�B ;:Zi݆�42Ƒ�}��_�K.y�8���l���2E�i�ưl�*:����5��������
��t�׾
 ;L/��|��k�ä�Ŀ��(uw�jۀ����C�C��w��6m:�6l�@����z����&�V�Tn�+v��xƙ��ɠ�_���(O��DA���w!��p2��O%C�m���`��Oe���L�|�k��x��g?����n�[�*U��	=���lN=��I�M��X	��"�����UkVb݆eC����T�G��S�VQ"s;��KZ��=����i�8��QO T7
Bn4�-�p}ݽ�h��t҉'��D�3���6z��t��(����5��:{`����B����մs�.��t�s�K+W��s�=�~z�/(��'9���\;�=�eifʿ��e�����4�w�[�Џo��h>��5�V�kК��0GW� �9�|�*�ǩnj�~�+>N��'ܼq��Zh@�%kW�N��ō�hn�!�s���=�{�͘u�J�H�����9�9s\s�1��sroKs�T+ۑ�Y�ߺ�)��:���;+jla,�ޛ��L�F���� 9c��ؼ�s90X�z=L��E����n����G���q.FKC��J�%uj�Ƥ���ښ(��Q�^�J�G6���|f+�P����N�b����S��$c#�4�93«n�>�'��0�)-A�Di���c�Vz߿^F=�LIl���6B{�R�a��ߧ}����EG҃n�M��1�m�Fܶc']�ַK��\�6	�<�����x�C��0�O>��#����\#�j���!?��Nɰ�����>
0�F����)ۚ�����4���_p=�y3�;�f/Wa��l�����vW� ɂEK��{����j�]L&WQWJ4�+ѩ��+��m߾����k�'?�!��~#���>�w�`vX簛#�ڏ[L������/���=���������2�Vuk�����i��AZ��W��D�F� �q���C�a<?s�b�;�Ff���F(8��g��LvI�A{f����۷c�az�.�=O� zd�.���v�e���i�P�YU��~�Jz�Ǩw�B: 0m6�Ԓ�S�\�\&�MUآ����s^��dz��b�e�ꄓh����/��(���J���w��_�%p�/[p��_�*=�=�L���ν�et��G�`U�L�� �[�*���T��r3f��5H$��։X?ޫ{S�Y��nm�����t}�|�����"|kU���ؘY�ɺ��v��
i�P�M�U�8�/S�Ι��pg	l���az��
�\J��6��o�N�R�ʇTT(�P*As�L��n���b�@v�Wkb��IJ%H��|�W��֖vz�e����)��:*�VsS~�Z��RM�6�N�Dyi���f�o�R�÷l�N�%J��u�E7��kP�0M���au[���;~+�ŏ~~3~�G���Nھ� ��)N��R�$'-���!���(XĜ:=�m7L<�>��_��!�[pH��}��{@��t�h�?��n��׿��'��G���[��=�����Ĥ�@Lf `1���j�x��ߡ��ݳP̧IPG$C��u���b�´t�rJ'�t� �
(�k��ڲ�!Z�bm{r�Y�;0  �-��� 9�a���*fY�u5�����|���R{O'Ȱ��pJ��+)<^��������G� ���)����X�!��\)�!��H1QH"��,�o`b����W��褓N���mO<IņJ���pH����z���ݾG��W}�;t��������-�K�GZ
���-�0�ι��������}�h�q)��G�m~�n�间c�c��=�.��:tx�x�Q���D===�Ѓc����ṋ��P�e1�M
+|�c�Ob'vap-��	�ET^"��޿�X,/b#�e���hב+lGj�����)��a�?E�
t�9Tز��R�COyvҬ��U1���Ǹ�{���.��\��ď�~���u�������$�d{��PԄvS���.e�l�s�5�;V�%,�"�eNg3��5����FD)���dQ�Y������U��'��8}����)�1���� �z��F����j�+�u����qF�k�#��M
P�:�hVb2��Hږ��#�����L󗭒�kNVZ�f9��	z\$�8�����k}���т� �L:�O?��u��u����C��{�V�����-��S�8���a�� ��C���w�O=����/�z�sk ��4?�rG5��4@d|l�&K�:;�[il<O��}4gN̟I��������9�y���O�sA�-�W����w��A�%�iŵ��d���ID�t�F-0�*y6��� ��f����qP�XU�2��j��?D���� ܷ�E���cq�[�PJ�e;�a�r���+i5��S�O)�6�W�n��J�Q8��p�F���ә)��M�́(�{�90�a��5W���u#���ki�^~1uχ���J���SȺ��C�����pc, K���w�Sl��944AO=���Ĕ�Mo�G�?pX�W�_��/�t��:hL�A�YW_�c�`�f��P��9��C�x�Rh�Q%�K��ҟ�DLfnR��g��֠^'?E2i��{�M#G�Q$M�B�uǬ��L�3y�V%���&|* %
&a�j@7l
�*�� ��P�b��N��4��*0�"�Vq�E�FÇ���T�5  t�ܨ�����LE�-�j~�^|�I�'`��Y�F���V9dfIODq��?�rn
we+1PeS��}T��
@�(��yS�祂��!싰��Qr*.͇��r#�H��=�dzh��m*�8+�HO�)����5�$j6�Ck6�FC������T/N���{m<q=}�_�O~�s�����wI��Ӈ?z%w�����,�$4�g?�u�KI�."��֨����l~��`Ma���q�a�"�����4T8H�֒�t�s4�Zec�0a�>^�L�4��e˩d�n������b-[�`�b�t�s�0�
T�J�D�Z Z���MR� D`����	���埠%����:��[�T��.J��ǆܦ�\�k�h�jR���0^@���a �h� �)D�$�_c�`����5M@2�-��%^���3��fU�/� &����_�}�hxʠO|�&>tٗ���	좛r0�d�BP�tF �Ω0-���k9ړ���gP�U�#��k�������?P4��Nk7�B�P&s&)�m��U r��܋
��c͵�$�q��[�^*(�z�M���L|ۆ�����Q��X�ܐ�?l��w�W���&�6܌�t�1����7f?�c׹��Oq���v?tŗ��&�,�:���.�X�����;_��J����6�a6娷�&7�Q��o�T2_e!�L����Y�����s� ��6ܿ�ᳪ5����S��7�d�������,˭:V�l<h��"n�Ja�-E�� ,���V�j�kjJ�[��L4��T{��CmmM���u���qJsض9BU� \�1����V^�vm}�Z�h]���Rс�Gh9�q����v��z��锓O��B�&�b8��#+\������糯���0�/�5�&�d
fh�����Z�&�`"�Z�Dc0�"�,ýYxm�b8���"�X��K�������՛Π���o�LO�G�8���m�0��P.��8�m��l�>����_��x�z��[h��e���]���ޖg�T��%ҥ·�o��I��}�`���0]�����Ǖ�`afQ���ߓ��3��'�������ZZ��w��~xõ�/���-\�L��acO�z+POb���Gi��g  �T4G x�R���E7�>=�P�
�ǉ��-�k������Z[�#��=�S��c��a��G��
����9�2��&)�Q�M��T'>�/�s�Ĵ�U�+yfB�_$=y���r�N˗�N�D�i���F�5,��Z���g.llB|M�=/B�MvH^��m�L�zdT����(���gK�)ӿd�����0��]���/�ΰ���*�h�d��L*r��DZ|u#/(N;ny�M�5���$)����,ٱk�����h!hv�Ď�>��<�||&��Dm�}�\��I�]Dz��g��Jw����P%�}��C�S��C:�Ib0AH�٤篢IF�dU������t�M?�����T�����;�H�rc�40ڐ�[\Mjp"�A$�����3m|�E]��p��;�) �+0Nwͥ(6�#`0L�[��&NmjJ�j0K9+�dԤ������}���Z�aQ'�a+��6� ����I�TBX��J���/�Gnz�>��+�Y���M���>��+i̉u˖���u��-�t����;��,���oz�;۲-��BBBh!T邀�]�+"��

z媈^�����B�		�'�l�Ζٙ�޿�9��f7��������-3��~�9�s��s�9x��g���G�3=�F�t̠�ǂ�}�R]��L��=I��Õ&��?Ak�P�9d��t�إ:3�H"��M0��y|�ߖ|�$0�u�0'ΧM�J�2��`u��W�g�3ӕ���J]�P�g{��u��I8u��9=����ur4aB�~��y3�z�>�<vnم����W��av��"�ȇ�ݦ��1�s"#K��P���c��ދOj��~��{*�Q6V�6V}(L'�KR[)���H��Ps�j��-��Tޟ����YטD�e��.e6���ym��O�/�`~F#%0��dn"�d�}�6��!�B>���).UX�ի*��A))1���N�`7K^E�"fB�؞|
�L�p�kE�6&�B$]?;��ͻB��[����	Ǆ:ۅ$�Ɇ����%K'�����!��-�@�$��[�ןy��s9f�6�D���|��x#�|�Mqȫ�MaE3>q��F�$���c�\}N����"��J�qL�U/J��9;F��>7��
h����bbl�|~��5�)�JiP�1�=KIp��Qi�y
��s��ik�9���mj�39�@��+h�˵)
c�u4�y�M�qƑ��⅏�Gk�t
�2�+�#����v"�܅DɌT��Ʈ��4���2y4��03�R��ⲕB()�e*?��j�t&�c�:�0�b�Ohsk�B~�t�Ԟ��S3C�N���~�''�uy	������-��R���x~: x��J�I�2ic:�^d���4w��t�����9�|��h��:p�v;�!Zkr&ܟĭ>B�ܮ/��Hv��/��:=���U'_R��|��h��UHU����q[2�ȵ�[n����
=�2s�r)�"��jH	��/�"/6M/�u��I%�XD(l�\c�T��`�ڼ��.��Ӯ.��+dD):�mt'~�>6H+?�[,� ("i�h��[�p�C��NCc��L������pi�I�p�JNC%(Yc�c�b�ʄFl5%�@�ݩU=�2݃�N#&�v�ǆ��Jnb�NL�]f�UM��vAuKV����~�uh�6m����̦����s�Ꮟ<�"�0�Oa�J�s,���P��-Mfm��H�Rp2�3S&�pPؐƄd��^�0��3ɉ2���\Q�a�M��<V���<xY-s��A �zr��G!�*�3�S7F!CCG;f��N1��:�?�ś1�׋]�v��Ё�ujfv*5��q|�k��B�DǂUBkQ ���s�T�BP5)I��n��~H�]S=F���qq�v���іvIx����N-���Q�E�G=j8}i�Lb�؋��L����U��7E{��DL-�0:��6ڃ�8vE�[�y�,��@�a�h�30M���L�M�Ă�%r@��a�V���T�T��R�KJ�D@��M�	B1��k{�0M&V1%"���L�������'s/u�2Qhu��}F;���
�/v`Z���/�j�΋�D ���C��^|�m|��<&�,�O�0�(�"9M�J���K�P��L��p�8��O˵0|�b11
�Ĕ����a�s�H�X3Z�4�d���C��dpVXK.ث!*Ԅ1�\����S�6Cr,=S*����$��1��v�=n��tM�4ݏ\���Ac{+9� �t��
�	玴��S����V�׼�������A�6��3>I������b86J�kY<���X��L�B��M(�F�L�ae�W
MB������P��!zf*I�\�k]r.2&��*s�J�"�۷�_*p��r�I
k"
� w0��vj�����ڌ �<�����M�ln�������G舎�~��+�o��B�(J:�891�.�����X��O�T�がq𤯠Q(#4q�Ƅ��M=[��B:զ voég�-�����p�(��B�(���XiBs�폦FV`�	8���s��At�ڼ�-a�g�ٷ��]]p�AO�AG�o�5N�I��K��@R-;5?�S�_)��?a�>�D ��"�B=w�h�Ү�~՛���_� UÄ5�S?#ԡ����~���W忔��'ũ!$%�%���hQ��m�����c(U�Ө�f,@��%��zG���#��)�q��&���I�l�$~��c8�J&�����)��DY5@q�MX�L���Ue�L������eU2�2��+��lR��TUq~�Y\6�}�.��b��rV)ι.�7�ƥ�(ɉ�xN��� �7���,0�M΢���~��98$�6����hu9$��i�����Aɗ���P�1����|~&S@Sg;��B}ٚgs��K�Y"��Z�.&�&ǗH�����TVwX��VrdVQ��Fq2�`��T�Pj,�'���f��tp�$T�vwWc=CB���LQ��+A#��p��	S��1�!��p�3�1鴔�5y^#�r,��<Wf�o�H`�������2r���8�ْ���Ȕk�=N�r.�F�i�~s񧧞�G	�ɍ ��H� �m܀@���6��	-3f�Mבf�//�3S�\B�;f-@oO�p�r�� !�0!�P��8����t�:�)���Y�����Xi�p�����$�&T�ԙ&c�O���Q�9�q N%Y�~��t����������{#�d����Hjzof���P*��I]�!�%G�"5���]�7�x�?
�GǼ��|�@�V��9�,�qY��Z��(S&5LHfV�S������8ν�H%�L��ZH�6`QC} �7�Y�� rR��MFɄ���5NJ�˺b�2Hu4n��U��N6U�Jy-��L��걄�0�G���I��Bn��(��ćG(d�#O�����ʔ�3�l�N���\<�(�&�$bI�ȉ��@����mv*>o�tQ��fRi���!��,�����g�<�C��M��YDi�[i#;9�M��3L"��p��Jrtʖ���C����A�>��K4k;wv�sf!>�{R ��c,�~H*"��������,�ɓȜ''��܌�g�*RW����<���qx��iU�"�s���kb��FKW����Fd�-�sb�e����j
�5�J�&Fn�������`�n�ڵ���cCh�脙7�%	����yQh�۳S&�c�1�Ϙ���/(�+��=?�G6��b�=ݹ�sy,*����j�t~Is�A�T3��M�����k��݃�(��`�/�&L=����Di���9���hժZ=63.��G��i�)��g�<�H|�����뮥��S3��]-��H������o<���+q'�O�VJ#����9eXPjjJ�"\M&-���i�����e�H�U��3�1�������MPVd=��X^S�D�&��w���O��I��� 36*P:�p�P�
W�b|�b~�����<��2�I�~�̙���I`�ӎ��E�Y�����)��Nh�#ʱ��:gR�� ��s+�12x�ƈ�f��F���*�w�v��0E��[�>�=1�;mh޿�:�
�\#������#��X��	�b_q��!=������P�}8&��ѦFL��ȸ6C#b^NF3��M��5q�n�O�xƉ	������BnB��-&rE��)*��I�WX���'���dI��y�$	%�\��S��DN6spG�ny�r��6v$`�c�B�;�!����%F&��kI�	��J���g�N�cc��z4��S�!M�2Eȍ�����E�5���h��!)ʂ�e�mBQ7�u�Ul=��yM�wiY^9����)Z�#���$f���T�"L�����P״ɛ��Z�`�'��/,j�W��<>}���9g	��f�%p|X+e�R3)W�b�;�q�S����pi�i��M�_���*�t�w��6p��X�;L1��P�Ք�`A�K�(�e�QP,��T��.�<eK�U���fR�"��ǣ�|/n'K$��Xx��Q�k6�ab�2t���w�5n�6�����a��Ƈ�s��c����_J���� Ͼ�ݧ���+��>
o�\i��S�g~�N�l�mV�ch�F�d"!����0��(J���� �ڂ�� A�2��$�Dsk�t�����xcׄ�1i��}^/9HZ{/����$�rƓ�bh�(b'�ܰ�	��l������g�c)r�N:��F���a�U([)�9����Z�E���][�.	�X���ωT�TS��4���l)�14�!�K"�ɇ�� 6����Γ���.�5O��L? 9�b��J��w�n �Gk�v��D���-Ía��C���y,6,tm�]`)� !�t�1D�9��#���ȵ2RfT�!�g���JP�/��[f �	:��ڷ��ӗ>u������������o������u6�ˠ�DG�(�^��EZ����t����k������Ż���V�s!"��Y�jII]Ԙ��"��,FU-$q���C+no�j?�1})�QSܑ�Ym��L�T���>��:9�TrT*��&5�Ǜ��@�I�m����l���A,�ɱa
k2�F����i��e��d��jt�Z��U2|_K���ĪY��c�~�0-l��n����E��q;���x���H�)Z �|��m]�li�(mT��a�&R��Oî�iT���F�|� m�Z;gPxU�X6�hW��">0�T*#J�������Y�4+�+�a��Q�!�pCD`��԰�L�=+6 ����	�B15E�B�P$(��ա
!���̠&�$��R)Br~���{0�	bR(M�W��q�f�4aY����۰�a�*s���]+�<H.���T��6%��(+[��n!0��pw��Mn�M�@j��zv#DNb�~�1N�e43.��C9������!�u
��A��,;1�V�M��=�+�T�"�!Pb
J&��*�$�9�6�pgo{��3��e��4������'�o�:�(�Q�A�O�_���}����N�1�v*��*67	�F��(]pV����'��C�UY��N��(M5�Q��.]:�j�XLt��&7n���x�9�
�
y��^�rMi�XjF��p@H�$���
���ۡ�����ׄ�-nE�+,�n�j]��ɝ����N=�ɷmy+�-�����|��A���n��w�Om�9��6�"�t���'T�>�B��]oc͚5��ӧ
o����af�2��jF���p�N��yk^]�/n�����V:����3���NH���Ilo�$��b>��:y���co$Ɔȁ䤧�%6y����Y'����vE��
�ŬH�r��=��(90�L��)�A(�C�2mL{�,�?���voǴ��B�HvK�0-sRLF616.����~�	���wbt���f�\}���sȓWmT��|7|��:X� ��yq�r5
-�t��Yr/^�����=C�Uc���1itN�0�s�߸Q2˙� w������4�}�wo��V&dC��C;��y���K��PM�|�6-���8v��R�̈Sߋ�{9M��\�i
��o�v��e��ԤaQ������<���w���٤)١�<�ɸq�%�/��W��<ͨ���
S d�U-�7�~L�wL�L�rB�K�<\(����1�&���β�yUB�$CK��UJf#��%�����G�6X�A�{����K�������	�shS�f��c� �>SX��s��������?��50[��<�@F��{fbd��y�I�Ӎ�n�<�7��O1����Bd����ː`&9!���k:��vȯP����5�lh�A�_H�B���?���xv�;h�5�`Er ��Ze0�;�?�J����3E! ��E	���ErtI2�9�a
�tx��,'=#fy�Q���8��L
g	
����e�FdM&��\�pd�;�k
�Y���=B!9�r��hЍ|:���N��>��0�$�{��chdB�C��G~^zH4
�����a"gg�`n@�N��׍m�%A��ʔ���5�"�c�\�ΏE�\7�@��������7EXG��{�jOR��u)dk&��I�uB(>'�0�^�B�`s����	�@6	*��]��{�a��H��W�x�|����=�־��^|/П	\,�[s# $Cȋ��*#d�L���h݀T�J����h�kyo��JI�l����d�ұ�I�1�����L��&��qZ�;��tjb6�<)#(�vt��'Mp\Z�� �Le��,V���l�%����+�pME9�u=��XF#�Q�a���D�f��b��-3���H(v͕�B�l�mw܅9K���L�P��\��,�z�Y�z�a�ٝ���d�h.��.��D�D��K�W�␔����v�F+!��V���_����+�![�7�p�H*�&��sq�a;:�%6Ok���K��i-��iÊ�_�so��|��'gk�7�������A:6 #����vNG��	�~CsAo�X?�a�����^/��\
��浯��Ł+���?���B8�	�?nlo��Tl\8PX��,ܪʡ1��	��uK3�����n�\���B���:��)�o#6Si�?�fBv���~�%�lan0`z�.K���!9�6rd�_3ۛp�w��}���;P�%)D�H�!+�Y)����z|㋗�'�'�x7��\.B�Q�i�D�I&(����"i��&�2�͋�e������v����Z��sf	���� ���Q���ĳ/�{?�)E_>��*����+᦮�;�L�1��T�����_�H���I�S��۽#Ld><��Wty4s��̈́����u�k� #�������҅mBQ�px�	~$��ַ7blhXtS��tښU')�P��;l^d(�f�X
ɑ߃��8
Y������I��tq&�el���R �y���a{���ش�M��j:\�J_���l��[�����b�|@�g.=�t|��Ϣ��-��Ww"OP�<���%�JL�g��8Ȩ��_s�6_|�>
Sܡ�̮$2U,[�D-�݉Dٌ����P66)���#'�SN?-Ӛi%
�Z��o`��Y]��t�������l�02�I�\�7sԐӌ���Dm.�+�!��i2��I��sr��"�mHr�t�H���5��\�ot
��3q��~���وS���j�CN<�t&I�J�l ђw�R����O��L��ٟ�8N=�X,�7m-B=`6O��-=��VZ� j������쭚"U�jM�����=�����Fv�����S9�6̟щW�����H��/��ip:q��袽��,�)�9\�����c`�pth�([���h�`� �	��8�ƫ�^�A���k�����B5�{�{+�}� ;�&|��U�q���oGE:��"��"�<���[�.�d�d�����9�����]&��k��ʻ~ޤ���zw9Ov�L޴�Υj� ���6��w�[u�J'1�З��V<��:<��C8��Cqާ�D��4��.1�Є�>�$�~�'rfJ��m�d+V�⚴Vs���߉�;��8FK������ؙ�� ��0}$TN���s'��Մy���)���#���Ń�|�z����8Dʜ�����v`�{.������b}�z쩵��-?�4:�+&�P"r��9P,d(�QZIY%	jgI��8r�"d(!28.�nذ�B�����y8�:� {�!�x�@|����S+��9&��I��5k��)w�l��f�T����I�ać��R�J���.!�JS��
��ta$6J�7�@��$�� tT)%���Mr.~;�3���N�b���r(S���4w��r��݃����C*1�3?z,�����y�)2I.p[/�U�b���$~������QAh��B�<fP��2s��t��Z���~��SU�*!��Ql�{�G
X��-8��JN�uy�1�n,փ�o�?��[��C�.��<�+���E;�(����&T,L�d>���|hCȍ�ޭ�jo�M7\�ְ�H��<��1A�������/mG܉o\�Y�}�eXp�j:Ä��2���Q"&.C�"h�R>����*�
u�{OM!��S���U��Y����Z6��j�M�jE��`c�)�"�lT�?d�E�,f5;:�?��t<��<���q�!�p�)'����q�M���\���xw���x�Q����cP0�isA����"��#�ú���ʻr2V�AûKHB�b#gT���0+�9¼����B��(�~�����֗.�>���n����������#�~����m�t2]��o��2N��J��m	�eBU�y��L������6�|���Qb;w ��r���cǊ�a������;�e�T�0)�:���`p,�m����ck�ʺ-��`L� Rcc����/2�:���L��C�5��M���#M�o&��FH��P�3�]������奥=^���% 3�����}9v32��z��";*fh����H���b���7���ς���f�|�$�-UE�T5+��r�F��,��{�b��w`֊UX�������Q�AMr��P���9vd0�f����A�W���N=�pU��}�oOJ[|��F$x�~�&��5��ɗ^�A@�Ï�3}X�dv����Ԇ$�R.�76w���1ļ�n��c���"C��C�9����:��b�������p����-�jt�pb����ŗ>w���W���9m�F�i������:M̘&����W��{�K��o�GcZ��s|O��j��^>A3�`8`i�4�+YY�´#U�.�k�B!��9>�k��<*�:�Eu�� I4]�Pln?��2f�c����ׇk�{'~LP�����G�Bc��C_�EK�a�;[��Ï����B`�͚G�I�v�㙗v�8�M��`�LC��TP�լbRc *W*+�+�&9��"MN�L�i�q�}�����;�~��҂�[�7�}
;���PL���M��˿� �C�M-�&��lRM}�%"��=NN�T��%��#'��Z�U���H�0��_�e�f���{|��w�gdcyș5N����"�f��M.=r�+?e��LN�"������H'���f3(�hk:ܒX����6��#�Q�dQL'�Yy
��T-/%���,�Y�O1�\ 5��6n�in�N2�ˎ����ч���L*tJ뵢����-��'�<�C%�t�Iq�χhszSip�b A&˔������F���jt{��(x[Z[Zġp���ECS�$c]5Ɠ�E2ƀ?��߃'�����OP�����������!8 ��*=*\VO��9h�Ю!
���|�lx�b�
����?�&B��{R��Y���~
�.��Z#3�}��p�5ߕq7T�RP0HJ��^������m���H��ߔ��T5I�kH�e_��@Y����' �~M�4>��"���c�2<V��棘C��Ɨ�};���Q\z�gp���y���b�!����ãO�oa�ׇ�����/F��F�����&��B��<Y�ZU��2'h�B����u��R�Ȅ�3�'�p����k���#|��si�a�A�d�X���|��������/�%C���/�o�Fl,!I����B�iUr����N�:�=�D�##�B�l��,6o�N2���n��-ݰP��	Z�� �a��E^S�d��'&�p����:2E~*��|�<��LȥX.`xpT�Z�M��9
�:�"�f���5�"UIb�3���xք����ym�Ę�(���9ஙl��x7K�Qha鏚@i3�	���W�m;���O���C�l�7�p5�''�KAC&��r���+IuN0	9��:' ��!���'RhE�_�Lɟ	Mf&{*�ó��($L�´f;�%
�q
�XY��t	M�����Y����Y�)��P��`}���q�p�I�A��C�moo��?M�s>tO�;vP�K��	��l��M�M�]�>r7��/�����m�LfL���P���ً�Dק��T�|m���F��\��L֪���냧/0��T��}���O�,7����S�5}kdh�����%@��mVb�Ч/�M!���i��s��~�*�p�*��؋������G(nmF�� ���yяS�>y=U#^�i��Ր!]��⒦�j� 9����Th3R�%Ș�y{vl�UW}�)a�ց�8.��
lܲMm���3k$��o�M-�����&C��&�U6�6&A\[��o⦛o�u�\���ze����p�bA+�/���MX���x	��ذ��oǼ�v�d���hj%�i	:��� @�H5�S�"�ބ�	���Ķ�)��d�Ź�2O���2���VFG�s��ϥ)�N���@�R�r`(B-ގ&��|��V�	V��v=�F
�:�:,�ݸ�;7K�f��MW{�>{tl�������Y3��!i�c7?y�r9k|��B�,[�w��9���y9t�@���Ia�:�Mǎ!�!v�3���a��tY��eJi�dp���wb�~�U<��+��t��^BPq�Yx^M/q���CHΉ��tX��͆cy�����G)���:Z�(@8tm���Q&�5���H�%Q�^��E�n�{�m�y%����<��z���ȡ�Mz]������52����W����#V�p��D��N�û�w�;x��'��ߟ��N<g�~Z�[���|	�:�<�4}����?ЋP�\��U��8���p���6���07,�%�]a��<�_����/�,dȹ��)z��hg�Xa����V�(Ā�@�6}������J�J���Bj���z��b�;��l��#L'�5�A�?�VrD�>��zs-͛� 9�
�N:�,_6GN1��+���C�˓���v�ΟߏW�o#GA?G�ʜV�[�����HsΈB�i'D@:��>;�0d¨���f�TT��9w���A ��
%
;�0��sv>BXųML�@!S���1B���E��
��u=�����α�]F.`����aFrYi\{����\�H�Cr���FEsM�tE�����:0 �g<I=�β.<�	�}6^����K!Xk���d1u�||����3Ru��v;�u��;��X���W�<LѨ�����DOZ�P�&�(��3#�=��(o�`���S�(擴ߒذa#zz7��_$mE��Ze	�<Fi�<Y�Q��fLVeޟD��n��3�:e��3P'�9�R�8>��{��ߙL���B��%B��%,1��6�*,�]�S��d��8�;��QkĚ����^}�=�[|ﺫ�p�b�<��� ���g�˿.T�,]!c�Ь)�[�����͋uhZ���d� :���x��X}���1�k�3�cEW�6�y��^��b\e��V��HWd�na4&v�	ND��\Y[�5�)&gr#g��4�A!�U�a�Ɲ�a�1��w�-]��&��Gy,N?�tB�����}*��^D���D�x��E�yБ�
'ظ���<ś��:���2D��d*䫄�̲���%%̀����42d�rV<��͕�ǧV���+��a��tSȖ�Iɔ�ӋW�];6�˾�K��B����S�az]6�7�41s�r�
�����_�z�?�-�mMغ�_'��v1o��>l�sd��g�|)�u>�\���p���?G�ۯ���&G��!�p�J\r�9h%�KQ86�L����뚍4�O��5�o�=���NV�$�ƉZ.B�b�`��$/��鴏�W�C�,����g�v�Ƹ�9�|��t�f�#�?N�Oz��Q�`�t�^�7�ὥ�)�#?�̧5�ӵO���<\�yWRV��WXP�'�3yh�}��L��tH���&ub׶�ЊIz�\���a���������դc��{μtvNG�hV�)%��PR0�33�y	��+f1�J�Ã�����.Ćƅ'��'�B~&Ih7G'���Z,&%b�9pX0h������-�k�%SՈy�:�L9ׄ�MJ�ܗ�Z��"}A�ɐ��L �߇Br��I�����ш�G��/��@��|�4�ɼ#�Ќ'�OPH@��9��L�̟�%s�x�:��B�̄p�t��%CV�q.M�)d-CQ�_�&���Ln�{(fkH's��3 �!:��C
� s�%�ú¬�K�#~�-�1g1��;нy��'���V��{�,_N���^u�<�1��< �Ww�ү\'��'
�q�<̒��,��Ӭ���U��k�nB���&�y��ݯ_z|��ab���܋����O�(ۦ5����d�|$���?�5¾X�Y��|������������<(�o�#��4����)�b�iC�LL��ƒ���8:�e�r'o��p��%�։ް�("�;�ywEߟ�'H�?SB�F�lM�M��ć�P*U�G|�C��1x��J���*��t�	?'�'݌�6�Vʡ�L"9֏��8��l��_��_
3[�6�)1�=|�6�����Ş�A�ۧ#Q�@C�N�j���tMP�U�o�����YN��f"���ݿ�c��O�6���gX�B����/�6H2.J�A| �_x{ƒ�.\A��]ȃ�����ԦV/���&�6
�����Y����E7`٢Ehm����鴷�PbES��������vb����l��V��R���O�����ٝ"�ϖ�G����fF����\�vB9<s��ѯ�<04��;��<=�4��Ѻ1�|�KV�|U�dY7�i�ˏ�L�ț�J��L�%R��`֜��\:��k/�����$Ξ��.Y���fw��x�8�Esg�^�qv�'r9�4lU60|�⚌5ɉΚ��?�'�^6ǭ:��� 8�	�+���XJٱ2O����}�y�Yz�T�J��l�
�8�i���AϏ�'O�Z�2yB�Di�խ�A��v��γA���.�F=^ᥥ�Pa�G�gT��k��(R2}��e����� EP9�z�d�a��m�\hM��f
'\:><�"5j�S(&ikg^yE��<�:��Y�C�0�E��{
x��a��!�"�܅�Dsă�N?�����l��e�ٛ�B��q�}�oxm��x��'	�σ/%è��R�_yu�l�6�����Y2&f���4&��P���-˲����C�F�[�D߂�LmCF/�%Fl�xM6,]�C�M���[e����Q�$�	�KQ��K��I&�\b�1����3]�y�~���)ӯm�ǓϾL��׽��~� [�h+8�pp#c�gT�3
L�M(�c{F� g�]�����ҽ��4 սg�ql�
�b����"���L>�s�t��a��y��O�D���?�#;I1,�RR�M������(|u�0��LR�tQX�4�^�_z�ݨu8�v`�B��x���8�ēq�G���ې�ub*�h'9�]�⩰��E�;�1��4����WSȁ�����K.�W�
\r�	�=Ο1�?#���(�{i-���F�Xt��K1��I6oU���<���49����T��
#�B�Q~I�T����g�kffi�I�� :����d�?U�|V�b0�Cu���pfTm��ӽR�!zݝ��<����/�sQ���G!��jUK����!�L*����������E��C#hm��%���,������^{���z���T/!s�XMx��xa�v�����;��Q,]~���E�1����I���`pfHH���"�V�L�<
+��H�І�)�;��9����.����u�l}s3fΚKb.��yTF'���g/>Ͽ��}�fr~~
=��e��<%3;�	[ۅ0����t�y|.x�ꉦ�<�T@Ϟ=��9�}��������Fc�%���c�RNօ�"q|��?���ɪC��{'<�̜� 6nx��
^|KN�w���^Y/��ZC��#1�jlmá�W@����s>��� �~BY�Cp��f�92P��mg�Y�!�*&�R ����zv���s�8�@T�~��;mشm#��^��7��/��#�[�����ft���C�>3��B�f�.1KU���Ȱ3#sG>�A��7�b�J<��sx��w0N_7FE�Ak�NO ���;�E�#M�.EV��ϖ�Gv��m�lZE����n7����މ���}Z�
9����(�v&�(��zV����d	�h�&��L'j�dm2yjpO&T�x�����K�dU�Q4�>�<��zd!�r&�.�$Ŭm_��@�$,qS�OA�w]( ��C��Il�P�N�v]��>�,�7��V3W'Ei.���峈��K�n�����}/4��~֊=�(�GF�g�:DCA$Ǔ�O�߶�a�P�7]uQ*��t�I�G�*��,y�,�n|�s:#�ލ�`��&(Iu:uȘ~s�p�a�+1,?p%}-�Hc �F��3a�U���ۢ+a�I�q��PH�U�3��
r��� �!���ƫO��+/���_��x�MX��P:�=�|"��d��xb=�;`�niES�t$�e
;4)5sI��U&��*��`1�ǆSO;Q�Ou�|�~��`q�T2+�%�H¥��+/`Ӗ��y�q�ʹ8�����ߟG����v�N\��(���� 1m���'��J�^y�]o��ΰ_���8��hn�2�Ne� g��#;Wa����-J{�#D�6J���#��MW�'�/�Q���	�f��|Y�Ϗ���8����\I!��'-���z���L�Dg������y$w���n�;=}�TN���Lj��5�űh*�s�b��GB�=/�O2�%QD(����)a$w�3k\��M��������I�25$d��&y��h�j������8�붦��v�/�9�^�X7���z"v��Zc�B-_������'�E�<��m�/�~B�.?.���عe+�^u>}�eX�|�̉0�Y�;�� `�<K�������38���\K����P?�1,�ن_�u#zj��k�F�s"u�hx���U9+���4���]��]hq��Wc��F14��٩���׮:g��Q\y��x{݋���u��}��|ՂH�2^�e�δ��� ��0e���*���\v%��$ʣ�0\o�qک'�J�e�N
�(�܃���� �-Z�֖(v�ނի�7�u5������_�D���**g�z#�-�+8[L%������ǉ���0܍]�a�/�b1��ib�Q(��܉;�w;�#`Ŋ���3/���#[̊k9)�d�N 3	4�8�E��!����;��9�.����M���ܿaU]��_r=�*}�Ȩ����MBs�r�160����MNφ�RA(,�,L�HH�A�slp�7_we������m>��[��D��4��*��Ҥ��}�)Y��iu�ô�eE ���k�	a�R�h&'�m��Z��>�1��0�'F�p��Ga���KL�褵��q���B��@ּ�?�[v�ȜH�h&#�kF�b>�t#�25���{��S<�FE��NH=��C]L~ΤJ+����s(	���I������>�`���l������jAr��*V�K�RElٶ;v���Fz�F14��M� $�"ܫ}�;���aw���|�K�]�ZLt���%V-��*��,���V��R,Ww�BVN���N��OaɌF�����x�g0k�<t�w�I��� n��ګ��[��⒡�L��L�NvKP:J�j]�یzLk6Rb\zM�r����>,����
G�:F�rr��̦��pp���B��w`[o����0�q��Ƿ}��	�v ~����\�A�M���������v�*��V��7�sL�c἖�8�d*���<Ϊ��==����B΍e3X��,z�E2���;1}�Y�,��>��9[\xm���G�`��Ǌ��k^}k7n��M���h�ac�������+>�[{0����[v�s�K�?��0�o�b��9N�DD�&�f|tǯ^*%YV�X�-���g,��
�?������x*�˾�e<y�%�p��E�keTJ9r�>io��	�,��X�
>��0է��dq��b�E��:U��p�KSI�r�^h�۬!�Ήb-s[q�ϲ�:� ^�W���FƘ+�nN�B�V ���\/L����-�>�P��Ϫ�k����;�r�¾ݴ��ܛ��n�Y0�ZED��7�'�|�����/HY��3ΐV����44xR9s+ť�ZK�7�B��Ε��M�e#Z�4�5#�U���0�e2"��O�Ǳh�|+�����oq��~
Gȏ��:������횆�_y9�w�����X�h"a�l >!͜y���	��|�p�%��qu�d*2`���;��Ÿ�Gw�9d��SހL���tt�PD�@{s#��_6�?��6��n��y5;Z�ˁ w�Ѕ3�*t��a��I��������_{���1���]G��V�l�օ�m�HmC�����]l���g`1���zl���qp�wb|.��ٜ��g'($*��Lx�a1n>\�_�۷�!Bh
�ּ���C8���p�׾�(�%���w4���8pU�M�z���1��%�\i�X,��u�qÆo6�Ȱu!�f�~�/���h�Ohĉ�tAܹ*��퇾mo`��n,�7��A;:;�0����6���g�ud��B:�T�P�_.ĸ|_l�C���$�vr@�4���n/7�U�)�d.�M�w3�r�R�cB����nc/R����{���E7jQ�-���vo|ƾ�ɤM����������ظ2��J�.B( �� �-���O|\�$'��ݪ��d�?M��2Cf����!a�|���l��iN����R*�Eu�IR����9�t�P
8�Ս����B<�����Aˬ`pǯƛ[z񣛯GG 8h�R\y�شaN:�t��b���A�1Ϯ�f~P�U-�������N6:�}�*�m;�J��/@ȡ8S9O�Ec�J���(>n��К�Z:��>��n؃��_�A�g�?A��0�������5,EV���$�
��X��sc՜9s��"��\�,�9t�b��.��Hy��:�����ӝ.d�[}~8�P�d�f���D�,�?�@ �do��!tׂ��5�3��3���-V��'W��Ea����-@��׃{O�,�����(�-aX�.�B�Jʤ�B!B�n�C=c��en�hcP�úw�y��s�����(�^Ap�b��j~�|�q(�GD�/e !)�K�W��Z��&�a��+"�����g���=����@׼K�TVp(�>�<r���@��bR��O�وrI����DM���_mR�G��|�!�y��(T�2S��f���0�jt��l�����?���Z5��]Y_udP�w�%6�������@��R(�iY�L82��<��j>_T�j��#X��;	Q��"o�5����3!�d�N"��8�clx`�Ѥ����Ua�ct��X�G��5�Q��*���� ˋ�n�|$ЊE+���[��/~w�pڣw�Iؽg�<l�4u��"GarEb�d�#�)�T�%u��˒y7�wm�On�^E�9F����8~����t��)@4�5�K/<fuȼȑ��w����h}ʴ.��S���Z��jP%�bA&k���bx4)')˸�DP���{�_�9K������uh�3�� >v���p�#>��f<���B��]سk�8��ibh B0^�$�1
CM�����\��#y���1x]N�N�3�A�����A�
�M���|����z�@����e�42��:�L�*O�g��pY�����n�
��Y� R+��p�5�t�e�~�:�M���L:Mk�=BM�ꑾ�L��j�2�L[�{h�%ȑs^�C�T2�[ހM+�c�矏�s�Mi��vD�B�l�{�a�����'TW�D�:K�P�Jr�� R��4�(�x�k�ԩ�ď���R�*��I������Y�����hi���.���r ��͓��m86���TS=�Kolė��u�D�v�"=y��i<85�řv!Fҍ[���A8�Y�Gzq�����.�Pz�pVǭ%�D7��k��Q�H�;(��&�Y�E�"��iX�DZ�t���o��#X��N����#�ҋO��~w��5��,	/F<�K�b�0�I����d<WCeD.�̺�6���s�2�F��.]&�?_�CO<�/|��Xp��7�)��ߝ@>9�77|?���8�
t8h� dp�0/���<D%���2�%�i*p睄���g��呶Nlݺ��߄���09�o^~	�|��㭗��E鮚Ea��t<>�o*�] ��7DגBC�b��g�6{6�6n��ЇT"���=h��sΎa��|or������'�s�P=�͚'��
G�fe�z��Gp�X�BFB>>4�O�О݄j�H'��e�Fa��%�f�b��h�bL�Ӳ�"x���hw7��D��nWKѳ*���7>��/��F��h���>!~�*e��&�D�T���-�}R��N�Ϟ�Z.K�j3R�-\�?���38���$�j_K��𙗷�g��^Y��3��ckG:o���M_4A�"�m��22�Nt�2�4�C"%?�M
���Z_�'e�gT�˱�d�YB�>L&�3z�1|r��������G:e���>�-�� U}�	R�ː!�	�e��y��
�/^�27*�r��{���.Hn�ޏ	�[���r��I�f�G�YY&bu����T������D��;B�%x&��i�Xnb��m8���d��-=�B+����f�}h�o>ּ�w��~|�sg�rj��91QXbr�c�]!g�O�N�m1J*S���:�вUt�LC��^�����o��߅��}5/^c�p��1gz6��[���|�J���v2[���7��߹]�"C�Ru$�t|��aX�Ax(Lq�lH�����/�_*Y�h���:x1�����K��\����Ϯ2�b����V��]��=���Ne�9�s+܁;����u$>��H�DC��qХ�^2:`\.�^���n�mn���]��Ƈ����������et�#0��Ƈ��h4�����ULS[!���Q"$�a�D2?=K����"Ȇ�h�Fx��=��x��6�z�5,^|�t2�)�ӫ)�����ڄO}�d��;�m��qx��$�A�J�s'9��?��a��"��8<���:�{1��_��+8��U�сť{և��=�<~��������[��i�	1V5��E�.���k���rh
���a���["�}�Uj��?��h*���n��OF^D���%�?}�Á���NNUG�f�)6&�{�~���]]ؼ}�
ft�,&_>�psT=�+��S����(W��0�����q�0�r�6���(%����[tV�S��y������Z�ɩX�x�ѧ��؄Շ�¶��jV4�}2m�afs�p׏L���>.j�＝�p�O��>�E�Ɍ��	`�TU} �9�Su�Q���O$���O	c�?@�08���!
)��'g�3��8���4�"6��֋�{3#�u����Y��L��Fa����������Zǌ=E���gQz
<�m�����?�9�i�:�� ��xp�������˻ə���Wʠ��^�ɰB!�A)�t��z�`,�B�SUaj�'5Q�0�!Î��F��1m���/'Tͦ��J����J($jjG�� ��ЄˇrE͚45Oø��Bi2�9^+!?�>'�� z�� Q�e��3q��_�=�{O<�7)�M�5|���S���d��<���H�jh��>i���2��1��I�yRN�s%�M�^Fk4��|��Ds��	��%'Fbx����<��6t#����ۦ��Gc}���<����Z�� ��Q��ఙ����{/��{s���e�L�'������3�ۢ��\U�X���G3hf�e��C��/��o����D��̺\�.�T�>B�f`î~����$i��(_Q�5}og��Qf(al�u湵�����xuc7��܍d�C��S(�V����|E<�kL�J��+(|��l2��G�� ����߽w��wH�tD���Q���������\�_���2�����}�bֲ#gRc"�8Gy�B}}x�(O#⧐ad�.��"-\0���44��E�I�Nan�ܟ�����P�y���=Y8Q��ŉF;9w���{Lē�v�RC�P�2�}:f�� �w'�{q��_��"ͷL.G�VQ4�-����v��[~�m{Fnm1�2W.(�;��<J��CϲqfF1��ƞ�~q&��,]��K��zd��W��b��Ǝ�a�E�LF��*~r�va����$���Vjȱ �X\�%>{Z�����q�M7�ƫ�*���e�p�y�rA}���6����ƺ��������B!�TU�qDL{QUM�&��K>'��O~'�TB*�J��������~���ax=-"w�9�	qz�����!T] _ 4!���,	����H������������nU�wW���}�ǧ��Ư��B�>)[S�ѩ��GQIZ���*X����2|�]t�f��>ɱ��)�U��b��M����h�����g�Xw�;b	hVZڦa,�S�ƃЌTV��ө<����LFX��R�<��붠���dd�L	a݉�];��܄r!��X?�d2�L�$�p�wo�M��U'b$o��x5G��$�d*�f@JAK�0N%�̈́�R���f��͙щ��>�}菄Ff�m�E`�[��c�m߆s.=O��e5�A��X���$���x�X�D���//�͂<��P:#=3���u�z�e��9d���#�ÎId�{O<�:��y8򤓱��_�%�O�,�(g��������F����v��_�5_�Xȏ�g�|�Fa�ȏ��kx&���M����y;��G_<'r.��� �2Ar����t�6�N� 90�l&�ǆ<
w[�=
���qL�Fq֙���!"�nɬ ����̀���Fș\��_c��A�N���3����D�����lj}ɹ�i
φ��!�	�)�d�kyˏ{,N;�
7(,Rb	�L:�l~/�����}��XzV��P����P#���w5�^g��r�T���3Y"�Ц�b�������a^�3B�!�Tk&3�J�]�����"7��&5	{tT$�K�ǍT)4M�U�>�^�d�d*�3�+�L{��v�LF�H�D/�Rv�ǈ{��h�0X�����9y���ac�
bC}������~��@��a�6<��{	����/����KN�T���X�{���nx[�P�9�.�Mm�uWa�8��g�z1����U���e�s��{��ǿ#ۥ������/��s��s��Mgx�Ў|���m�p�m��
E� [���;kN0��=ެ���a>qɚ�m�ƍ��A� �=w�����93��x�8��2�������I&�tH�$�"ET�U��*��EVvuw�uuŮ+��R,�&Hoҋ��{2���s{;��>���;�忻�\c�d��s��}o}���3��:ڥ��Fh���i�%b�eq$V-�(��
9R&���[�
�Y���io�˗����?��:��y��{d\f��υܬo�T�6� 9�H\��H��q�W�Z�x��__�TSlp����va�U2����/j���Q�`�.��m%���7�v5M��O~䓢�P�=��)I!H�_ٲ�����3k�Sg�"*B�["ي��Z�4⠡�ln<*,y�|�ɹ3���*�$�(�D����]���lǈJ�=�{�*�EG�X,���-�s�Su�@�<8��՘4�[�'
�4�Q�}I��_�/�{6�Ϡ��%�_oI���|�7�1�M#�� z��2d��kJ�OG'�ȑ��&3/�4�T���릓I*rH�9����= �¦�%�����ŕpa V�n�	 �ٹ�����U_��\Ƈ���c�m��q�S�N>	,�̈́2	Gw$}�SO�m�Xw�H|�2[��q2P�S0x'|�^��3Ny\>3f�A��>v�{8�qi��N�����.�@D�æ����@yi�l�6B��ᵴ���fFhx�H�� T���`�9Wh���#�@�F��["4�}3-���|�*�q�v����m����zg����H���#�}]�{��}�ї��ڻۦ�Y�)�h�ز�׽,��`�o�{L�uP�R�R9Oϣ-;�/|����x��8�l�'s|�J��%]+��	Ϲ���ӛ�)5kU8���pm�����7*y�̍R���db�0��u���>pvt���0}���Jv����mt��n�e�-��]X�*e��Z���Kl@Bd�1홷LZ���Wm5��-���"l(��PdB����D�^�1�$�ȍAL<oԖ���:NX��kl�Q0�s�Vd�s��S�h� 9E������o-�tQ�ɟ���^^{?՞@Nt�B�Ok��V@U�|��a����xV�v#?(������뾋�DJh� R.��`�!m1���7�;l���ڒl|���եn���&P<����bޗg�8�R h�B_� R����2:��h������i���t�G��N?���$G)D�8��Ң���j�P�s��}��+)����SZ���D�OM���`���E�8�l������.|��t��n�ζ�VL6'Z��Q`.�P�����Z�;:A'��vZ�i��2$� ۇ�5U*
�eE���؟�~�B�m��n�Њ�t��w�ƍ��罋.��A�j
6D��̓8�H��?�"�|�ڔ�e�
A�R�M�l�[Zb"�U��E��]�9���/���_^#��qGK���{�����>�Hvq�6z��g�o	�3��w�Rڵs�9s�262J]�6_gT�?-���X�F�l�F!Ko��b�̥�8���K��孴f�zz�մ}�>jk�E��>6��;�JN<FY6F%^;b� %jjU�����0XZ�Txm�Rh�s������_�t3}�W��ׇP&�F�>.�1��O�����5�n?=��6�ac�h�b�7Y 3�Q�� ���T�c�0�����e�@=�3�Su #�����5a+��h�uߤ���9�)�i�����)��@E0D!G�ɘ�߼`�ct��B&c]�Oc�9�����B-R$Ԁǻ���w/4��U@m��q�[p09뙢c[��)�mٖ�M�-[D���J�mn�,ڹi���.��c���0�I�,��W��}�	�ܧ/�|�|�CZ���8{�{.��C��kS�muMH�P���!��p�Z�hV�R�흏�}w����ڕ4a?{��iN�ǳ�0�۲��|a-G4����~�	4&���#�@����5N_�\��ƪq���Myl�f�$���Oَ\���ܻ���茷}�*�W<�;4H��ͤ(���'C�x����K��'�&��@�������/�AO-|ؓ䔳 ��w��m��h ���&��ƛhr� }�c��?w��`o`�����P������k����J�ᶠ!ܠ�ٽ2�� ��#�=�xBt��1��:�^�n��?l�#.�O�r�?H�W��u?���~'m�=Des��z9B1=Yg��*u%�H�	NY��E��ʏM�i,!���:��I�7��SO~-�?W#�{�Eڹs�c�f����I�7�ɒ_�9�g���B.�8l]�վ���8I��b)kpƛE�i�c*E���1��_9��[j�XE8��Ly�%C�X�78�oJPݙ��yj\?�_}O�Y)�:�z*z���7T�U��`k�ZWϜ({�\�$G>�5M���HBH�:D�d먣�`0���Z�|	-���>�!x�������ӊ�t��o��]�!>�azi�+t�-�
\��_�uv���w�Ǜ�Dfe@����g1�<t������UR�I������d�r�
��I}����|�{�A��S�2I��$��ѳ/�Q�5Ё8�A�2��5ͪ�Q��v),+%�<�L4�k�6��5N���h��x��g)m�9G��%�̣DLM�[��T������.����O��$Ŋ0�W*%VZ�\�-ҰS�Jȣ��)�Q�>0��-Gcx�N��s?����ǡÅ�9W��� *UO��aT.��m4Qs�?�5}�Rx�%S�=g.aX�Z�R����xI,*UԨ�4�.]�˛�����O~�FH����Ul\������}?Nw��~�C;���˖r��.Q�p!O6*�N�fqT.��#G2�1J	�AcC�2Gt�>M+�ϓu��'�/~Ax����oЊU���'] �[�s9����.��f�_F��H�,E��)h��{�AĮ����*s9�[�ȼd˻M�����8A6�V�VP��;����յy���6h�b˴P�)��@ƚ��(�WPQ� OMt��	�$y�ͅ�E/��(�y�SbV�z���ݣ�Q�kK"P�WPpĘ�ǀ[��S��'_�]
��S�M���h|�H��/���=��V:���l��9/��1G�A��]�i���ITʗ�A�D3�m����,L�ru�xNDpn%Ǟ�ӅZ��_S7��%��~uۭ�ҋ�衇��2A����d�
���/�"�;� =�g���
��=:_^�:�2j`�QqMeT�PȮ8 ��/����JF�r�G�<����rx���ߺ�^۸��������p�e�`�|[�J�$u�p4!�9����0�'@iU�C��_�>tv�ڼ{�Կ�͚M��i��Mҝw�C�:��3(Ɇ��ӎ�o�������c�Q�3A��ec���q����a�-e���uZ��(6DI���?�G�h\x�����Co}˩B��ָ�F��O���*�}m'=���'���[�Q��_TG8��Z�(T�BCfz��U�}��T��B��^^6��l�z���(?�:e8"��u[:)�C<�3�F��w�UW}�����ܮ�2�
�	u�1U�U2���d���|�9��� A�M�MØ��Ԏ��b�Ҕ�u�$�g�V�;����gK#�S7�C/�cz�Z&Z<OG���rn��U��]� �LK�S�l4�S
��ej�KC��jl=����ﲌ���zH�3�����R	C���m���?CO=� m\���)�њ��y�h���t���'h�Q�iݦZx�a9�r����#�Q���"�i�fhxS�.C?\OGL��҈���Ӟ����v��%g	c|����	���߻�Z:��%�d���q�i'җ����9�]�F��yy�B�� =Q�F�/��6>�VK��A�������Lf�uu�*
����t�;�H��4"ŇB8f��c�u)��v�Qd0L�jlT�����~����mغ��:�X>�O�e{� �Q.�78H��+%ݽ{��4�|���d�,>�9�B�pNL:�)�T�:���
4ʑQ���M4��m�����N�Lں����}Ud*N?�8z�g����Bi��E�����t,���~���n��^����i�����<^{�G����̍�n FF�Nc������$͚��(�������?�>�dnX�w`L Wx��ixl�N<�4N��t����BrnFۤI`�\�
*�hCw
Q��I9'Iw�9�3fs�')�.H��3��_A�SO����O���J��r"���)R���k���ģH?[�i<���7�4$w$!��HS�ȁC�4�[�dg�7^X
�Ұ��穲�'���
��S,�P|l3��"h��z��S��|�1����.iaCS��*������~��_�#O>!<#�m�i"��z�Q�/��\�)�?a�7����4�h��{�;��s��m�2�����-]'t�����?>')ܥ��+:�%��	�z��B�
g���MLi��M��ȠđV4
�b��mc+|��1@���?�$[��V-��f.���Ȉ<�B���74�w/�2ݔ��2�퓟�I��&�&�}��l$���7t�����!���Q��Z`�OL�R�4IKV.�e�El!�z��W)��%iÞ}�t�ч��I�O�yףԷd1�����ȗ�2Y���C�a��"�ݡ���4w�!d�l��$h���)KSyb�6����<�e��W7P�N��K�y�iժ�)7	1�}����Ǟ�A6�qN{�ثh���V�<�܄�G�S���\�G�{��5����4����ݚ����<��y��u��ig�"F�`4�a>�2��#�
zHP�e��c���I��C2oB��t8�*�k��t�SjI�SaMU�D���������+�~S؆}0uy!��Ly��@�����a��5�U�V�Zdjb���H�X_h�S�	./8�JM�A�#rP,OA�)Dǜ�#M��Z+��kJۖsqHx �YJ~�\�L[�����54�w;�b @��)��D4V�<~��4cN��;{zپE�އ��>�A:|�R�Rؼ��4Ꮖ8`(R
2��&�c��Y9)�����1G��k�k����w������O��ײc�Nz���h�!������ؤSO9�����q����|��WBT&�!WM�
mA��p��?c�O�=z��.]B���S�$��ܷ��-���z�E6,6��b>,��5nߴ���H��f�RC��\��|2��!����ҲC��@C�˯T�ՃG��"=���Lghtp�88@�,X@��]�8Ω�dI�B�QC�~(��P$KY�� �޷sG[JsD ��8�Ξ4��5��V<K�^[K���.�Q��Ӥ���\Q�̤�	˃(ˑ��ir����@� ���.�#���!iiMK�l�-��_�$�kCcY�0F����a�_��m;٨�Ŵ�x���v�FDn��`�3u;W�aC�su�R�Yq�����u��9
J(��� =�7�z�x������J z�, ����A�Q����Jcģ���A�	�2�T�s�>�J�A"��Q��-�2���cFx'!$��)
�t��)��E,�DF�56�3Ho� n���a~��%����G9�x��;Z(ݖ`O��G_XG�x��m����i�P�h�!,�\�b�x�C�-��f�0]�o?�t�S��s�6G��5�<4��#qq����42�P�m$��e�����u������^��x�����[_���YL��T絘5w&�fG(&��^��^b�y2��������H�g�=��:��#(��F�������\���X�����!��<���~�KC��G��Hy�HΈ����0��oҖ�P,����1:��UXZ��G�]�s:�S�%dJ+{�s���_���"x��lޱC
�Ü^�x B�T��b��	X$N;c��Hm������"6�@z�T�-;vR}r���8�y��t��?Gs�'RrdaA�����%z���h��c�ܨ��#���LFm2-��}�lmcØe�:��o�B��iт#ؘN�5Z�-5h�ɚ5;����"э�H�	��'�W��b��h�04"�D�t�S��{2��������N=E�9Z�����-��Ų#���R��A@�5�婿7���Ԉ�Ƀ��L���d��Q�ڰ��xj
9��H$�aST����Z���̽ѐ_HŢ�D$\�S�P�T�ర��}F(<;
u�d�F8T-L�M���	�!i�Z��� �f�x�܀ �l�ڦ��Ň	 ��Q�k�:J�\������v�&�9o���+3���Ș <o��WR�{y�:�ըu�!��)s�0���7�zfAr�K�b�8�rujooa����Z�z5-9l9U�
��(��qNm6��é��o��a�dK�(�U8���-m�0��t�u��3�З�%NL6���2u�ZH���Mt貥�pF�Zg͒L����i��|�2B�}�9�TP+��ذ�sF�M�ECR4��0����T�g�<�����ʯ^.Q�y�zE�Z?l�dA��u���uj�=>hZ�t���V�4n��4k��N���l� ������
#"�|��)YBD�K�^`��<���c�x���2?f�a���\N�gϡys������ߢ�C���#ld_���zI0/���٣G���
J����]4��j�t�����:���ȣ��[ǩ�S�l?}���9=�G��A^�^--
 ����Æ��34@m�Ƒ�[>|��� ߯�$�4 �s��]�	u�������T���6$�QS�2F���FU$��<�l4�t�
�������T��T�Ӑ��������ɍ�KX�3g������<ed�+�v����ۉ��F��ߙX�zM����.����g��彳�ͯ:nO�0fU�aJs�v6�%�h�'F��By8B�,C�5�;�O�P���UB�T�KJP,�4�s;MUꞽ@�ۨ������R��vڸy�,R����:BT����U���5L�	A�1�@�!��%������{��G,ovm�E'�|�tp��x���9�z���KG�=z���%�`�jT�Ԛn�2Ƣ9���	ը�d8��0�'�yCe������������Ga��|�1��W�Ҳ�G���;��S�U38���4m�(��M�H��땪��!ՅZ�P��IHuv�Dy�����+���K��c�CJ3��x���t�o�g�z�>�"����t��.�� ˎ@�q + E:)��r�#�0e�:(��29J-a�����ܞnZ8���7FWϽPA;OO>���u��ӣ��N�:�/�2�}H�]�H�0�(;�rqRH�0;Qȉ��_ZM��x$�li�V���/�J��Y�T`�;F���ǣ�O<Nv��HE�Q�w̘���yo� ��4��!;��E6 U�3G��8Uj9>s�	[�z��֪%Jf2��Jͮ׽��Z�?	!�K5����9�����&��
���>jU!^��f�>~�B��R\B	��A�ë
�hp�pxbl��V�,<u�yg��g���s'��ޟ|S`ir����6�����s߃��>�ԅ�}k{���E�c�C�����Z+zR/3 I�9��95j��BX�*�"ML1�&%m�7�k"��0/�W������M_�ǫ8��(#��o| �jP
�(>���1E:��s�`Dgo[)�b�FT�D����?���~z����߹�lL�{�u�V���h����B��#��$�JAϑ�.4`����i� ��ڈ96>�ݝ4�u�ڼ�>�O��8ˆ+$�n0ns��$�S�Hk����f���Ew��0�->�]\��Q"4U(�tc��qv"�3ht�����1}��/HT`ʀ��̻|����WtȒ���=�N{�y%�D�2�=�ˆ��	��%�hH
���y������K���t�}��I�&�=P� pb�v�W7n�;o��vl���V�z��i��h�xo����B���=�ڹ�����2����}Ԗi�x���������:R)��E��}�6m�H���Y���G�֮[K���}��ߧE�(���	N�gu*�}���;�$f�%�_vF��A�;�)4�������c�xh,����U�ŵ����(��Z��-Py�.Ӌebv4bږ�Ga� ䷩L���J�A	~�00�F�$��D�5����3(��s6fS�ZU$+x��[R�j��c������{�g?��߿���{��ſ���O;z����ƻ��z���~�5+��V$Y��ٌ$��b���?j�WBsE�=qh�'d4� �}MA�� Z}ˏ��sסK�ˁĀ��=C�u��cPԂ�f�Q���\��i�&����eCԀ�����8]��-Z<��>��Й��@G�<L�;�����D,D/<��<N:eR	��1~�L,͇��
o�9h��8WC�*�E�P�MG��K�{���ZMR���S�<�g������(ɛ��SDL7�=`��P8 y�0 �2_Һ=#���*z���t�Y�!s���GS��Kt�1s!�a>��^ڲ{�?�Sڮ?��m�����8��K��!J��P�2�j�7%H�(�PT �ܠxW��i����,�c�>zn�k���k8e�EGtR�Pf��[������F�����cl%o�s���a9�ǐ���x�^Y��6o�E3�^N3�z�g�_Kw�y��z-�Ty>�-tĊ3��3�Jo?�d��*�|?��u��)U��-�)qNem� !�a�����:GC=m������ց�M�_��[N��ŕ�-�-�YK&�Zٵɚ�͖B[b/�����[w�Vw�U庿d|��U-�mm�T�{Ȏ��{�P:�&zA�xZ�Qi��b�������q�-��[O�l�Yύl������/����<c���Y���o���ۯ��No��t��/�U�	#�Z��]���!eXP��k�Ug�\.�� ��$z���Ñ� �o��5�ח^�{'����b�2��(�Qs8J�g6���+VF�@*TGt�@^�L:�;F?��5���~Q��.��_PH�~��i��X�G�h2��w���1�8��ʊ˖���-�"\!�T�Mx;d)<eU�H��(Hr��%����$Ʈ(���:�l('�jKwЬC�T�� ��Α+-��f=��!]�R�J�(��ˏ�t�L�GGh��5Dc�dv͢h,I�3��I�ї���ZRIڳ�(���|�+�����)D�8�D������sX[�6����>I��z�~�Q���;�o�"�1o��f���CǗ�B���(���)�/Á����/�.�Z��N!:�H��v��G_����O��1Zr���?'6Q��9t�bA	$�O�����#�KVI��vn(̩i~�Z8�C��(ey]�d�U��Lmz����Ξq��������,4��������u����E�=��Y���_�x�D���!m,_����Q�P��<�=����/��������_z�+!�H�'��#"������ҠcT����/�������$x}���F�������}����R��2`�Q_A�l�@aM�T��l������)�2�r���C
/��s��O=�N>�4z���%\!�h���P�ug��WԘJ����3�(���і~�g��y�.���}��V��C`Ί�k��	���s2x�E��O;�rPW���yN\��)����]JcS}iF���tuʵ*��a��-j�#�:`l�;�@�đG%�m��J�=����k`J�
Q�9�/RWGU�40ι=�P���u2�&��a�˛y�̙BA��;���q�9�Fǳ41���!J���옥8SL=���50���5�5Jw΢a6�����At)=� ºzz��)f8�Q�8���T�
�sw&�y="Ѕ��а��R%��5�s"�'�)V0-<�^��*]p�������Z<K�z��I��IJ9���ׯ��n��m�|ձT�$�
��4�9-� �iTP�᝛׾p�K�}�����~�3���C�h����]�a���<�R�+����Jn1� m�阽ut���k�1�ki����n� ��
��t�ĆV6�ޘ05,���qש�t��ι�/NZ��@}�G�ⴡo^{˝?��oV��.�1;��Ԁ�U�DS�4x���D"@І��|�*Rq��""|bN���p����+vh4K���741>I�����o�ɯ+0�S��b�j�,ʘj�˴,�Z�,�,m=s�o�x%=��K"����E��9Z�a���5꛻�(�ЂÏB��_�v�|�]4w�4��580L�Ni�C����ce`nÔ6<�hγ��3�%3$c��X���Q�H.[�I*x<r���)��Ĳ3@+�[	N�0���MD9h�¿��ɒ0��J�/f�����%_�TF�qk�B�8U��K�w�ΐ����)}&�2���;6;��G+G[���A� h�T��N�8�+4�����zA轵�[�ꘚn8";��r$�(,���5����F�T�5��(-[u"��N�ȥt��>��A'�r<��h��0=��Z�7��-[���]��ځ�		����C�^���K��I&�޻��}�?�����ᰞ�����ʳ���u�����>���v}�o������'�~V���>\�,�w��g�j1~�lL]#��,:88 �-���}����o �@Fn�:�ߛ1�g�v��{����O��ş��׬�}d��u����R`2����&�x�4�."�*�=��pX����3�^5�9�P��ا��o]��WِEc4&�	0t�)��psz��Wcm�M�oM�JN^(7�����:;��7I�exd��?͇���8MZ�ㅽ�ů���zY��R�AB&����0��I�5�s5��/��!����<d�ᎊ�|��($�E4�{Wk�ע���R!��H�V�����4�.�Bi3MU> ���DS��d�"��r�� 
�'*XH��������p���G�H�Fy��*GR(��z�HcE����lԁ��e)%ErGH�Q!���*��Ƹ�6A���?3��H�Ʃ�1��@`{���	e�$�92)���;:(��FC� ��2ez�s���'�~�~?1J�~��h�P��O���?�S��:���P�sTRQ�q2~�������N��R����޸�=x�O������1��:�����y[������hb劕t�+i�!�{�'�s�6�Ag�����p�u�SK�x00*�6ɑY�4�cn;bŲ'��k��7�uȜy;���\(WO��&3��;2d	k�L0HeVSH-�$�šsP�4U��~���� R���"�kQ��������	�w��cD�t��)kC���,_(�f� �Up���ޱ���X�^	�{ͦ0ta8��V�%��j�R�o�u.̴��rC�o#}h��&���˟5(�Yj�A��������h0�����U>���J'T'�R]�|<�kjH� #`#���w\K�8�VE`�P��lM%�T�>"�a}[2!#�m�i�v��P���1*�1d�Y�åSq�s��)t����oWv��xo�9��j&G~���&��H`��B.�3M��-���͢@�Qu�=ÑGA'x{�)��$FeT �Đ �l�Rɸ@�s�9����پ�8J�5w	U2�R+K�����J� E-a�۱g��,$��*�z�������un�:A8#�������G/:���K��s����m�~�_O9��#'��_?�o/��4Q�U?"�at�0�
��ٖ���w��&�x���-�x��ÉV�\2j���S���Mzs^��}���O?���6NMF�I�%W�aCG'DM>U@���z�/�@&]*G�� �hhI�kklPj��(�4)�=�i� 5�(�!�'�\�:ӊ��.lƆ�jb
��C0<I�Z����r��3i6 eN�&)�u���O>4�2��[,P7�̣`�UoЄ�� ��En��N�z������U�(����q.ORT���б2��ߦ�1�j �԰+��N��۠���2v���fH}2]�#DcccdU�y٘�b����{��[���a�G����(??�"0�u>�6�U�o|�F�.�BG�� rL�[d�!�i�Hu��������,��~:NLes� #�7�AE NQJ�ד�C�����?�F]

�0�6�3G>�5���":���0!�������'G&���x�|��Ay0�=������׿~�97�v��/�p�|]gk��M�/����Xq��:E�j�j̈́��e�?�:��{E�����������\Og��Ň��қ�:�9ً?���c�|�ޘ*����t���P�0	�_�,!:�6rs�[x	MOM��<���՜R���)p@^�B� �Hi�����W��/ɑ���0��GC���sx���[�8%%���ْ�bv��n_G~yT����<o���jA���RnpLIDb���������60"����^�82� ������{ "�%�D4������k��i�ib����u��Ī�}�>c�Sۮ��,P�-:h���5"��}�vm�dg��W�8:��[G�:E-6��<� �m��A�L�)x:�옢n�]��T#|�QWQGyբC�&F)����k����.��H�xDI ����� �L�i�QC�
�0�:)�m8�:CD2�in���S���U����6*�Q-���}o����| ��)G�秷�~�Oo�y�%+l�}R��T�t�u8�S^���4(�����M��8������Jw[��\èқ�:l���?��\��c�=C�.��f�pl�2��b�f�f��p�_���ߦ��Ԁ\�x��� ����l4��hQ�{hҲ M�!���f�F|!p�UZ8�+E	�0B��(}����<�h޻��!�ACZ�E��=���Ã���_P���m;h�7�$%��9,7h���T`#�
�fJ`�`hɷJ���sH��D<.EH*PS���L͠Gͮ���n���Ü�%������=R)�{9�6w�����h�� ��xG�y�4�iN,P��k"�j��Xs: h�KTTt|ڹs'�Ϝ�������9Z��	�V��6��sU�� ��8:�>đ��E��.`�(P� }X�� 2�.K��Yx��
U����6\�ѐ����� ��U%M�4Ňm��
ahu|��S�⮁�}_��}W^��~v�8���{�yx�÷ec�Ăx��)G�0�ZB�(Kp֎&[ߐ�bKKa�oXf�No�k���5��k�N�0���(�O�&�<$��
P�AH�=��&^�T��4�g�y!�,�2�Q�\]�D#��H�PA�!��x�Q�J���q���������aC^��_�K�8����'S�ӏy��WdEa�|���"hm-׌�d��8U\�˨#�LE��L:�&��Yz�D���ldl��T?'��M-�5��*t�N�V!��;N��|�Q��l�w�e�j�U�3 �� <EbM��rH~��
�|=c�޵7��?Am3������x�p� �_/I�X!dÞ)@�F��]^HD�00�s�u�sX�7pf#�2T���"JI{Ѝ���at�c�	�XM"�	Ψ� }-���Ь;�rgg������ƫ��cl�a�o���U�N��`��� ���7�o����g�X;/�á��d��_ȫ�݀P�� |n	}^ 57#��V�Z��	QS�AK�U֛�z�Γ�C_�HG� g������Vg��(W�9o�����Q@n|BrT�q�Z�i�KclQ���Aɕ'褣�Q����W���y��Ř`�7� Z2D} �G?,t�rp�� c{8j����rmg]mD��{�܃�=tDm��P��H�h�ӕ3�,�!��A�g$��zJ�y|�QR���뾐/a"\]1Ƞ"
��k˞��)��Kmca_�q�qt�/n�����G����i�?�j��IO�R�ԑ�S�M;���4DU�0�Qz�C���K�و�.C��!�H҅2T:-�����d�<�~��#�'~Qh��1x�Z��x����o���l��2�(���[n('�7#N5�p0��6��LC�
�D$�(SD�L�o��c������M(������&4�M��6�cH|��J��mbTȠf�MЙ�����a��/xPT
E1(~�!�BoӨI� �0�C�S�����,LA��p_K(+2�n�.�ΘE�������i�Ј�ě!p��T�Į;�9�S���nܘ�6(��
�c�h�Bjkk�A@S�UUu\?
�,��3��O�/&^ExL���
ǃT�ҵ�;��(�9jM�}^�b�Ӗ��Cƚ��Ddd��*k����i��Kǌ���O�(��~ϯ)�.
ťh��(7*20	�k��f����M1���aÒy~��`m=��L�"j�p��$�_� P���P��?�D�,�6�<n��#?KQjx�K���+�Px ���f6$]�5��AH�m�Q��-�X�M<>~OWg�u<_����Z��0���LI���Oy�ئ�*$�t����So��M~��r�F��ٽ����/��S %=���Qky�8�:5~ӠL�'���E���bC��Y}�!F����:�[E�tlb�� ���L�aニ�+*��`*�vR1׻U1>f8"`9��m7I߾���?���M��}Xt����"m��K��5��:
����P*�Z���;�3���F8���:�9�Q >E����!C]'k$�F�[��ºHT�I�Řf�=WGQ0"(d�QS�k��N	_����s��܇�z? �9�-�53�:gΚA�-q6U�D}�>B^x!�R���	l�̨�=G��$z�Hӥ��5�����#�À���J�C*��ܙ��|~Ē߱�;2V�ϾRR _��T]����	+�?��J��3T8bh�1�/�ͨ��jl(�i�K���d!����
a�^�������}+����5(��~�w �0�}�U��:D�u���Y##~���xӬ�6uqH/9j�R��ep������|(d��F���ij��A0Tu��_1��S�@��Mf���ڤR6'��m�2'�y�&J��4o�<ڴm;�"�P"�ѳ���#���8jf]�JU��P+i�P���!G�F�&''(�L����&������)b��:JlPJ�o��M�Q�HU�T����3R�H��$a�%�p���S����#5*φԘ<_����BS\�5ٖr�5dRؓ��%dʶeheHW�@L^��(79NN��k����*Q��G����aL�Bӆ���M�D�	�M����Y?�Q���f44����G��2��`<.398T0��pH��@U�P���Ա+Q#�ߓAҪDs�U=Du-Rj�z�|?���O�'=k�._vl��N��G�&:��{��+�I1f����
\OΖ
��[<�:5���/���~�9�N�hf������<�?�����凎�� ]+5�&�\�
��氠D�.|ŀ/P����(��kRA�Fd.#2 �$pr�q����ƫ�ߡ��E\��6�n����b�Ƈ��x>K�w�>�����U��h+yHW8��9|=6����.�Y� � ��P���p���٠ }&d���t�=_?XŤc����W������ �tmU_/��Ă���u16F�c�?A{�hX�nFq�TK^�YLe�k��Q�J�T+�ЖZk+��޿�9���l�$F�|�c)29�i8&MfKQ��Cɓ�f����:�Æ	��_�涤v5��/1]�&Z�&�{|��'�!"!j�d�ǯ��.!�I�\����@����C-������������\�`"!�X�i$��b��;�s��}3��F�^�L��QP& U[�$�+~Ty�7�M�O�+0h�#I*O�@�/9Q,�ۼ}',�^z^vl�ܸe�!�=�q���L�Ia�I��M�6��7u�[(��R�˲!U�n�)SCUUp@��'8Ln0,$o�Kȏg �I�>�G/;w�|>'�&������DU�a/�V�/���-�D)�i*8U!��~�<{v�V��a��ׂku�E94���ZYEC�k�
 ���B2VyQg��P�i؉@�M�&��ǯcP���~�����s@燯���kF�����#�6�����Fl1Bh��XR`-'a�o�d�Ӏ�k�>�ϨgX�ԧPS�M0ڃ'�Q��cah[�[�~�DB��	�����7�Q����WW��lM�`�����E{X���J�]�h$�ϯ��f��p�2X(�r���F���2��bWuE�������O>��[%�a��X�B	L��Qӎ$>��'�r����d8��w�9#K�U�^�t���1M)M^^P�"R�}��G�O���HC �"�F�x(j��u�1�U�+�M0�.ښ�[@nDb��zU�I��tJ(�ĵsπP��J���4����*	\��q���u�wО=#�ʳ�Ѷ��?4j�ņ������V)v�j!+a;9��*��������t�O�XI]�.��ӟ(��T-I�PoP�!�+VN?Qׁ�G��¤^J6���8e�2
�h�yU0��1�UwB��CѶ�:����YÇ^M�w`�O�faOZؐs�A������ɤ�G!@�T���<�n�j�����qK�ZM�oWI��:�@��\���5���/;�͈'ܒ���������'�_��+&v�ٳ װ����1���F�q്��+�Dժ�ԯ�yO�\Hk������~��g��AY�vW��C�֞�U/�q�H#;6um��Ę��7*�B%M ����±�(P�"Q!�S*ZF��z����aYj!7
�@]���ލ����Nݽ3����Z��j/�ps�Yx6\p�'b�xէ��ݳw��Gߡ��n����-�$���h�������Pͩz�Q�\G�z\���K��"�ht\SeB�����Ј�0uTH������'����q�/YEe�)��0�`D X���)��G�Hߧ�k��'�Y�R���z��G(Q\��?�����o`83CQ
�*5�	r3$�]��y*ֲ��2M���s�O��V)��2�����@T3���+����>�Z۾�}��Fd?3�g	K�k�~<�H-���;���o:���=���щ�E׎	-*
�fX�<��ö��3���:��ml����:B��c�5�k�3��~������K���ӏ�v >t�:?��/;%[�k$�NE5�R]����:01��D�9�%2��0v`��dJ���Q�	`nou���=
m��i��8��Ԫ�$S�"_��j�'��_� �AfȜ��[��eiI�apR����x*%̐�&o�w	�9���*#
ҵ��{VQ�FO2�RY����ɨ4�u�T-�(E������� ��;�~0�u����&��P��A[FZ�&��!T VLIQ,.;*��{�`Y�(�-�R_G{�r�/�Ɵ��2p�-��RUI9��ki	EeXu�P���a���R��
��ܪ���DDM����b�6��4�����4�(CGņf�W �(��=��q�k�S�o�T<����Mo�������N�ş��w�]��cN�T	�jJV��	�oz�mՌ)R���z��-N3m#�p�ƃ��kT0j��ڳGF�����[��}y�o_�dן�y(P�ˏ�:�Ǟ�L��s�N����Ê��iz�p)�=�7M�#�)�JU�Vxz<D�#0u,u]0D��c�/D��J|Lm��� ��>UȌ(&d	|��R�+�S�{W�ʭf�l*� sF�-T/MP!����>��HK}]$�#4�2_Q�8U��=S�)��-��@
�iM-���\m��\�?�
ɰ�!Gڠ����_���J ����q�I0���R�! ?��i�]�!}�%BP��* ��R�T<��J���VR�4�	�Vʓ[�TvXD@�Dn���_TT9�g��@'
d[1�>izS���W5C�Szے�H{Z��!�SW�!W���u��u6����1nKq�� 42�X������k��k�П�B��w=2w��ug�KΌ��)?"5(��Ec��aZ�������^�g	0˗�w6����QĎ��=}�����\s�y�O���%���A�_É|��ޏ���N|��W?��ӻ�-H�iϒ.��>�3��%8���"Ǹ|�* 2�T@KeC�Y�S��o��	T�4-�Vh�b��j��i�D&HP񏲧��xtV�Y�Q|W�HpNX��8>����)�p�D�����`��"<mC�`�JC-!6�U��ըܦr��<������i���`��׌F�[��-F��4jB�dz��M�*}�����u�t�Hu��ܪ�;���TT�3NsJ\�ݝ� �b4M��R��0j��R�#ԥ0&��R(F7R�P��]�aX�S{����a�2�f��i�Π @�}]��x�DRmxL�V	~I8��gh���$1��5�Ҥ1H���_����p"���3/\x������3_�7���Ï�3�/��,�[jUO0>�BOM�J:~׃jP�a[��31�U�t�H%���WK�Lw��6m���W���/�{�O�߾��C����X�={�Ğx�չ_��\�v㮳�.�76�oM�1b͋�H��JQL�����(�̤RN�ݣ�H�
�V�η}�0@�"��tZ-��+8��
sV �Nz]/�A�͘:Ԋ/1��C*GSJ�����hbx/�l��|^lo�����b�K6�F�b�D(|��E�Y��˿�̩t&06�V"7��4̄`j�=��p��N�����餺�:����B;������6 ��'�5Lϥ�ч@�y�`�l���¨G�1*���P��8��������)�A�܅�*��)k��seVGm p4�nM�8�A������Uk,Q�~���7��^��v�����I�<N�:{f����^��o��/��g7���a�@�w��ɪ�N�N��;lG�4�5�~ �k��C��u���U�P(n�Mm��I�"T��=sI��� ��v.2k��/n�{��>�������]O��{����V���z-^�.�F������Ė[���k����oo���3f/�Yn�H��9}]dI���F0fx$ S�ć��,aG�2��T���B�������A}"�3>Ў�6�@����xm��M��:0�% 23H�+ ��ү=�xs�1B�����}t�	G�w�N��vҼ˨=��o�	:�D�Twц��d#��F�Nꨛ���t!�
>�:��L���"��W[XRhR������Y�{�~W�<4mA��X� ��UB�W��e�ȑaE����������"�(�*zI�����
2&�Z�U�kyy���� W�a��$9�@�!|�5�auo8����Bc"��A���I
�!C:M�X��f�¼��JMj�~�����S�D�L|�H$�5��]��}p�6�VWs��2��3:zf�����K/��O]��K�.�_�6��?9�w�=��=3g��L�5�+P�*�k�0m	����a��f�|}S��)/�W5_�16����XWkW_[�\�w�o�=��[o�jo��h���֨�r��:�}�#3'&&[\��e#�m�2����Lŵ�{���j]��i
�����$*��_��d%��[!9=d_�-	䨣't��+k��␉g���ʃ��c�Rѓ���� *��+r�}�Gȡ7T^�w�g�.�֖�DRP��u%�cS���k��q�<�T��_�'8�d(�WT	ꢕ7r$*PW�v�D=5p�z^3��J0���U��|9�Dڐ��&p=�Vx�'�Rb�Gj>���Q�{�b!��ׇN�-�V���*��U�BX�>!^�x,"�{��5δ�J�+ʟ����<�?��pD�f��CQ[G���;G9!Nρ�������:���QX�\�4�2�0Ξ�@��j����uM�)c2�T�D��u�(zHÒH{N��띿���3�{�.���>���.Y�r��u��=C���.�􊷬߶�H���J���lS2�*�� ���F�I}%U�j�o�?���&���UKV��5�]
�x,F�&KU�����=��|�����ʱ�@=��z݋D�l�Ba3����Q��T�o嫪�
2"/�*00X8�+Q�_�*��kC��oEYж���.OP�����ψ���A
E"
�d���ȥk�����ܳ���C�#5H�Y�ӚϮ�ߪ�$u=͌�{ѢC�=�E���B܅��^*�R��7κ���Be�H/k�vM�3=�buI�\�j,��M%��SW2�pHg�R�{I�d7GQN9��7����)�J8�s6X�|>��N�x,5.o�
�.�0�Nk�q�zH{g�w+����@W3��jT�h:7D�Ar���}��J�(lh� %�i!���`^*HG
���H����k0��D�I���$ ���}}s
A��~0Xُ�dX��P��׃F�I��T޷��ْ�1����Jy�~�����;�/_�d�}�Ǜ���H��H$m��F��j�,N"�|�GV<��3Ǆ�C��΅�3;����A(f 4Y�hapS�@j��:<x�,�D���oNu	,�L]b� Q�{k̺���tD|�U$�Qh�EV2�!��0 ����*�`L�o�G*%Q�~H_<Β|�B  ��IDATݱ9��Q�S�,���(������u�;Y���p\A	l�s�ܿ`M�"��6cЎ�E�ڒv���uu�S2�D�BqK\�T*%�x�7�&W��!�Q�?�}a������N�������V�eDb�P�Z���i�bEt r�DR�s��I��ŤY�y-��EG�ӯ�G?a�a���߁B=F�Oa}(a8�o� ��C/��&&�lpZ���%E��b�P����$ @�]����Z&B�x�R�&-_Q6mh#�ҘBE:��ߛ*^�R�������(e��d�6��f�J�2���P?�ڒ�9 �����T(�Je�S��F��կm->��l4�x2��V*���6Gn���]{{[KO���
�k�ǲy�C���$���lPj2���F(���j�jB ��K;�ʔ�X��aV\������b�:��AȊ�0�?�*x��b�R���jx�t��ٲ#j�I�ו�1���B�u Q�sU����%�e��e(.UM�9�%wC��� EX�آ�ʸ(oM��D0��t@9�Y�����o�DpL�6���u�������l��U34�x`�>����6�����m6ms� *0<8|�rY��a�=E�{U����� :�$�|��$�T�߫�U$����E�Q*��B��
��e��;�}�����#p����pD!^��\��g�֐",�D00<��fd�8��S�1��qĜ
�hET��D%�xu=>#]PU�@?(�+�b�5Q0�\鿿���H�|�R47��kOԬ�?�kjj�˙jh{�����B����ez^<d�:Z-ʙ�N8��]2+�x��\��K�T���&0Ҙ+���ʦ J	M�����#X�#�<�j�{�H5Y��K��,ji�����5�	Q,�q���dU@�=�B��<��DLJBc�����4�ź�H�W��	�J�H_8TwU�)�=6<
ʞ�I���D" CU�}M0=��ÈHK�Ҁ�ǒa�R55�ې�Æ�r_��U��IHiA���F�U����	�<U䳤N#�GJ��R�%����c��\N!e&s(��a)�c��9z<��w�+�4U�C<�Y,dmQ��a QP�>R��f�ԎA�DE�EX���R@��p0,5!��Uƒ�}�'ӆ�h���1HjXw�0��Uz����<D3ftK=)���P�rD9@$��z�P�ÖN�8�����T�Xa�/�t�J�$�������>)*OOSؑ�Z|��>ס)��:a�E����F��Hn5K�N����k�I��1�U�(���(���)��8Ĕ*@�&��v���-�Śaj���W92C�ʓ	��� -�^Os���n;�%��릎t{T[���Ħ�h�,G�0}
����A��GBeJ:l7$�P5��>�.���l�G�B��c��0*2�䤥P�2]v�jE�8B<Kj+��H���tF��-�w�����&�~D�C�O�ڏ��0-5��(J`������5Nv�H�A�*�F��rY���[{��1�I��U��p��D��[K{v(CPWzI0EN�PC�:@w�r�߿ƿ�P/�e�nr2/C�X�\aRR����P̩G�B��J�}f��U��9M[�`���S[G�*��-�����ͦ�K��d�vo��I<�j�*�Ut�֯{�~���hV_��y��z�\���[������O�͛6Ю����O+�����3��;�]{�p��x_pB}IQ�?4����:���A����r�I�Z��a�fzJ ��;c�����k��t	���r_�@
�]$R���v����3���	'��ʞ��+�
�Q�H�RR4�D�J���o���|�fy�r��j-� N�k��0W���wx�"�E����f�nPW�ty0|��7o���a4�o��J�iLC�N�����p�F��sP��?bs��j5��^�.:L�~��>R5�p
9��Xi��&�ޝJE0@q �	GbRjTI'X���!0�י��DN6��������~6;>!��^�0���1@]��{B�`(~���>\Q�]��x���#���0�]�l��[�]��z{g��%b���˫)��q�0C~v۶m��O�Z���ұ�ˡy���:�sĨ�^�x"CW׼b�
����z�� �Cw_'���3�^��/�\j1���7�裏�����(=������M+W��9�g��ȰDS˗/���s~�ч�cOP�.�~%�@�#F���[�)��I��a�vK�QЕ���M�i��W�4;8�������/WwM
���*��?޾N��Z���ܓ��������$" �����3 �(HE�""9G�#
&���E��,,�s��z�S��~��[]�;3���c�����
��{�w��I�CS�m�_/��U6a�h��S'xE-nV]�$R	�V�	���b�v������E�	��=�u���tvqq`!�U��!!���$�����*��?��,�E�0}c]��r���*Ok�W�:�
�s��F��Q�ו��3�Ӿ:����?�F�1VU]=��'#�I�d�5�F��E|�����l�
P+%���^P�Jc��S"�(�9��H�rV�RD:��S�j}��di���{"�}�+� �z�}�#�7^/���r78 hd�YihlƊ�����o,\(���6ي�Q]��`�{���S.p��͛~��uC6i��=�;��o/EsC3�� �ԬR����S�Q^I%\ioo��q�QG����e����x��"�Dy;����V�Ϛ9[�k;z�0m��������Oc͚58��c�=���CQ^�R�6{�44��������� y���n�D��|*.!X:�����u�qr�0�������Y}���D��q��Z���#Y<a�	�u� {E|�D�+*�Q ���/�YZ~�hk*��)y�~i��`4���(�x�BO0aw�#�(�	=������i6�Jn~�8K�W� ].���=u}KE�����ǫ�cOw�AIJ���BsC<�7jn��d�3�*�2�����FǍ`�S:�H���;�[�5�T�U0����<-<���S$#d�KH�X./FL5j�WR�\=�И��d~X*���e�J�aO���9��<�!4Ԥ�����q�m�"�X�DV�tM���˪�ź�ux饗���(�ס��:���� �˼y�P_S+�������C
$k�k�x���*��{�}?BR�/��*�|�M,Z�f͞���>Z�ɒ�KO�S����f�wÆ����>}:��~�m466��-_.�/�q����顇�h~Tэ7ʪz�E��B�o�=����v^�?}*����4hKo�+n˸��<(z_K�,1٦����!׉������%$pl��ѓ����t�hζ���ۅ��'J�<�J��o'�NJFI
:P�`�M��Ec�Z*�;ܮ��g�ɐʂNA]�+ǋ'jv�^t�|���H��#���G1&[ �Z#����y���z����+j�E��:��[@�X�똬���l�rU�^�:�0�|zP\���.g'�B�V���Iz0n�J�ɶ�L���\]] �H�Q�2��ǖ��x���òU��M�k93���T)�х�+�! f��o���̻P�nQؤ��d���[x���ຨ=*ǑɫuTr�{y��Gq�M��w�e4T���2���{$L����g�3�9,�xl3�&֜f��+bHt�\v��N/��;��#�<"|�#�8B��ʕ+�^�GN9E���~�vK�/#v���������/Ƈc�F�g��,`��/��Q�{P-�!D��WpJE��<������+3.���T�?���N�Q	�Z��	��Qq����-^�4�WJ�d�@�F�]Vm�)0�\����֘T� ��S؎�ٛ�=�|{��<��{��[K�20:)%%|�h����as2��1$�(�9��G���X��)Jf��q���~�rT��4�v9�^	��~��鈇���P	�dQ���(IӘ��[�v��81[��kz|i@�oiĥ��x~�+��É��O�U��ݣ�:#������hI�����c�*C6�Z��6e�h,ػX�uO���x�r=4@�[^}�et+��y��W��h<��H�eZ7C���3@4��RImಢħi��L^�*��M"�jjۂ��O�7I���Hxr�:aQ
k�b)���c�;8�w$CT�{�|�4D�c������d2��<�����b(�O��)���p�������ϗ�h;��w[�mkX�S�F�`8A�)�C>[`p�S-L؟I�0ũVbǤ�$O>
=�\V����'�'ӊl����`%��ZW��Y$�*����{��Z���U	�tS�B�� �ᄚ3g� ��X�ޕ�+�;��$�����
���%40�̖"/��L�Z�BV4�$q���Kt*��kn��8��Z\MR�GR������"�w�:��W]]�}�X@�w������>��qY6Q{_�8��I��Y�<��^}]�c�͙'�׭<(����i�<B BE���(�I� ��Ĵ�����`h�c�Nlߐ���H���R�,k�,Q9g�o����m2v�A!���xASn�+A*�4#�Ŷ#K��Z:������ȾE��D�����P��:����(]yR�}�j�-K^;��Bj|"*@-e��e*����t��9^ы�}�N%d��Ò)�$�Y����!a��X)�C@��l���1��fFC<�����pEb�3�%	� �mn4��;k
��,�S�v�6�W��Z9Ζp���P�4�x�$)P+�Ν��S7�rKjQ{�Q�2�2���;��ų$�3~��q�:O��H�゙Eɹ��ۢ\>ű��xV' PKc�k/d��XU�+K{'Fb�}G�6*��1�m����	>Z�K5\zLno۹!�F�"��I�B3R��Z�!7g��T*o��l����Y��EƷ9�痨rd��@�	U0�,��U�`K�:������\��u}+Z��f�'f8-$Q�B�m/]�d�1�环BvP� oC�"F�q���!WjTR�aV:U��/�Tw5al�S�V(��3M��}��1Ù���%��P�u�<6�I�Gt;Mҵc�8���Ȩ��T2�%��(hc'�7"�]�t1Im5u����b̂60��-+�9�~�M���es��,L�Ӛ�:��bE���^�/4R��F^��bx	��^�!�)빅vΖT�,פ�`T�ͼ��}��e[C��7R~��AG6v?{M�^;y�s��T�"E��Ajc��6N�v��~�[�C	��jD�n1�$�*�d���jـ��͹�&e�hKA���4H�ڸʋ!h+�b�V��%�L�Y����4��Kcus�xGEO�i�hQ�(����4؈
EM�@7��}�58�]�I����1�Ni�q=��Jc���vNt֐p�r�|����	)C#u4��g����A��t�����(h��z*��$+�yL���<']A�o��r�c�B��hƬ>�.�X��Ŷ�[�-p�P� ��3\|SJ {�0�xdp�m'i8�RaTF�g{�ᶆ`G�J������D��ZL�����mL��~��mq
���\��Q�)y�⦎v��I�rl%l���nH(t���,�:Y� ��,�*e=�ev��$$ �Q-��[}
����<;����aQ��HO��Q� Xd'�`ͫ�7��!;��P���Zݐ��j���r�z��P�}O7���^�~X�Ɉ��<���J���$�5���DW�!��$A}�����!��,�OfpƷ���|x^B�#�d
3m�?k��0]�>�bA��x�I�+�G����m<����2�5YU='�:T7��qB\�:���	T��Sk�d%%��E)p"6tu�ץ@��Q4<��}��eE��W���k	ye��>?��f!E�7��K���9�v[�l��<��}O;�;`G����Fv��N�o�F��� gE'�UR���[��pb����Қ�7R�lzڲ.�iRI�16�*J�GD�T8C� J)
��Tji�{�V�cڄqش~r�:�.�Պ�j���Fn /%���U�da'�O��P�^��L�=��[	Kk`��Z� 7������J�뙴�"S�Ƅ!����){2�g��fBF�uD�@�i��'�elp#Ya6[CDB^ƀ��b`��&�Ly�t�:P�c��0���"Z���{9�{���@1�I�p߷������/���������Mث������|K.��O6cS|��c,��#׷)����ߣ��HPQ��#BZcW>O�#Z� c6'idNJT��e5�0�~���(ѳ�E#E��t�+����=��ջ��v wp�?���:��/���y<�n^�*j��	;0�a{HY������,b�[y�3P�xN��0����=�M��V4�ONh�2�S�������
�|��}�����BU�zG�� 们+�`����)����7�ڈI�ڿ��S86Tڣ�ڐ��:��oԝݎ����D'�=#�mkzFc�N7��54��U1���f�������<�14�Ka��R�x#%O)����D�G�v~���)4�ޭ��n�컋Q>�C�*L̓�xF̕�� �!�bj��m��U,��A��I�>��+ł��2,asa�2<����?Ӈ5K��*����@kK-���p�>�`��/c�%�{H55�:Q���Du*���!�	��8?4&�, +[YFB�=x�D���&���M �:�6��5ܢ��.@��[�}-�^㡄k^|�ͷ2�(/�Tt/8�=>�I'��_��W�`9���}���!�����WngO��V��/�+�Ml9If��ƪ[~~�8)����f-�T�߾;Sv�c�y0��2���{���^m�a*<T�cl�	�SJ1*]H���F���,�dTp��粍��]8�zYO���T�=N]z�WPQ�b�W06�h}�(���7�drD�F�x'r�j�?�D.�&�
�_yM-8�=��+_��<|�v��S@wfL�.8Ȟs�B۸���?�Fo_/��ㆸ[��E�M��h�d}����z�W`�rn��kE'�!�&k���`�J��bl�
F$a�[&%�ii��n��1�����S4lq�Z��עZ������`?~��������{)���̠�P�K�P�ASS#<ez�����(�I���ܦuO�H)i�l;�t:\�3�vv��Y����K�v�Tf@���80�������5(�Ο�h>\%/d��C�;�8l����[��h*�2�ފ�J�Z&zY���'�2(`f�oM
�8���ˊ^���49kףs]ZZ�p�U�'���Z4(1��nvLy79�'�ƵL��F}C�T�p�MD$T���p!K����i�U�}@i0YL�N {|߀�L_���_�R�D���t�}�l���?��R6�<S�B�[����DKV6�6����b�X�HvnM:%�,�Q^fUV���� �Z[���L����"(�Q�?<���qc@��c}4�e�nF�)��z����'��CG�'�*��O��ak=6�=JͿ�㝄�����4lW=Y9M{Iq\eb�c$�Dwa:�6AU�,�*4�b��o ?؋���_��k��)T+��;��{H`K��;��_�����Al�Ҏ���G��3�;��K/c�֍�)/`:
��H��;��/2|�(��v��6 �~�P(l"�=s�A*� ~���P ���(i'��6�\Ɛ�a�d�ў�I���o03U%E�s���O�c}��u�f1&eٿ�\�`a훷���]��2e��d�2�dyIE~���q�aCWb�[��n��Y���Ѧ�~��r/IĈ���K@��D��BCg�#�S�0����V6��<H���������t�AE���<"R:)�'#�ʄ��#H��FG<tw�c��U���3����i�0LB*�s�vD��@O���n�������$UyđGb��⶯߰�=h?�9iA����j�WJؐ��%����y5acQ�:7�aaXc�h�!	�&t>-�d�f��q|�4�|���8��>�gF�AR��.f�sb
�
���w|s���x������0�q�X��U�1{
1ӺV��
y�&ē�74p�����̓K����jx|{�(�(mG������G���CK/d�uAi��_?�;�Aw�A)�.�9>S��ƕ^,B����I�� `�߭�w ΍��*O��1)�I[k_�&>g���BD��j���*�^y����e�67��<.���11�L1R�8���6� 7��]�ѻu=.>����S���:*Fj0Q�j ^��nT�����=��o��_똬�@S}
�!�V�R��iV煃:W��B"�2N�-���z)^(_G7 p�$U��>��Bp�<�]ڪ�h����6&��4.�`IY�)av�,0�6im!x:[&a
��kB)=f*�$�?)/Bbv2iŹ����S:��x"���!����m���:q��_����_��=��HTՠ��U����똩��z&��)ĕg�"	�Z.R��S��xL$��*�2��'���2
>9���*�8%�T�q�g��Al�t��\�-r���q�]]d��N�z�Sƻ�ǌ�\pq��yp�;�;��Uz��b�$�K+�_ZY]�L���~�5�P�� �M��j�ԩ�C�T�(�Gn@c"�&W�۬�2$=�}8Z�x�}��x�a�޸�y�Ԗ��Ӈ��A<���xc��x}��{���鉤����۾��Mju�t��u�z�i���
��9�4g'f`��:�B���#��X��cz��I��B7ө_��x.pj�-ȓYY-�������J�� ��am��kJ���	XOv/7�F��;��ɇ�4ȣvtu�����)��a�L�؆���e�t܇p�w����L�W����T�[��摹���&c���\�g�īumTFo�P��e����66p���Ζ��|�pCa�'ŗ��sv-SրU~�!�k��}���[�?"?�b}�[rM���I$���6�UF�
^TO�{QaP�54������c�bt�*�9����~���f�v�g�qX�tn��v���,_��'OG�i�J(�[Դ�f���[&|>�JҜ�����ia�Z�Ԗ�S���E,�c�O%�U	��!L@�J� ��B����mAI�|(�����fJ���b)ݭ�Y1�
��[�}���0�NN����u�~6�K���oO�����̘9Uݿ>̚3��s#>��ƃ�3����ȵo��Y��ڔFOG�0l	�P��I�9fuXf!�4�����Y8;�vDh�mG��XY��%H�>��&n�m;ՠ��K:�VXt{��������bE/�G���P�9�z!0)�3�Q+>��jU��T�wYĜ�1�wm�@�uo�Q�����W��>�Q�����7v*W����}�Dgw����`�L�Y�þ�ʪ�=�=cۇD���'t�JCUB�����!K�F����Z�ƒ#��v8E�I1�L^���AQ�w�m�ՍY ����iKk����$�Q��68�5�d��>�mG({l[����]��PE2v;#R1^g����B�Ù�\��O>���P�\+�����?�����_�{�qtttQ&�Z�T��K���j��I'�<M��%m�ϱٵQ�
w���w0u*���6��lfO��]䷣���mE����+�ؚ�P���oP�����r����B0K���7�yEkl�XDO��r�j��t�}�J�q�e₯}Y�\И���#�����^��w��~���h�<�p(��0���A�'���^��I��#)ר�~I_��y|�K�i�*<��Z)�)֤A6ǦvsF�X����W�s��*1x��I~�:���cl#���m]H�s)��!Jw���V�`�ҁ��5��,S6��$��=��%�����)%0k�l��d)n��N����������	�4��TX��P����O?w��N<����s�AM]�t ��J��'���1*G�}�E�rY̨9�3�2�9j&;6�+��Xca�-и�q�,���z�L0Ɯwt;w�+��V�j�Z���iV�ȚF�A=��?9Hn�_�C����ACM3r]���܄!�}������8N8�*��gs%���)������~�gl�Ąs�״���
k�v
����EF�RQ3��d�R9���xA��T]*����#y-����A����� �b���C����h�F� ���<��7o��6 �yD��W�����������l���$��*;()�ց�`�����m2�Z�
s��Op�ko�w�s7.��B������������?��������!�O�:m���BU�JBXM/����%3�Ύ��/8 ���=
?��l84�4�y(�av<�\ZqF�Z������-�(��W�b��U��'M7�SP�����C�J�X�M��WWT��\�VtoZ!��_��'p�_V�B�A�έ�������_��a��`	v�s�'=��4�ʣ`�?����*��'Ǒ�B��^��	���C�WN��ecjP���˸�[���~�n5x#�8\Ci��:��t���Y9���$�ň�������cz2{^����aӷ��S��Tt	K	�3`U�|Ǆa���Td�UZ�K�n��\�V<��t�L�S�'F�'z	eX�jЫ~O*�pܤ)زq�:�̛��zک8���Q]��V%_��� ���g���ǞxF���-M,�$Ē�R��b` d�"Fgڌ���n��6����N���s�E�+�dc۹��u��"������a �p7BZ���!f��X�][�����2�SeѾ~�2�����GwފY�[�KMU%��+�q�7/«�aҌ����#��S5�2�EY�4/B��{���bɎS��-f���eR���S�)+w���
�V��y�8�a6᪓�\��=��l�*��C��^w���3�FG?'F�K�A(w�C�2�e��Q$��9��*�w���1��p�E�W]u���2fk{L��shQ!{-Z��2�i
�T�^oC�8��V�^��.��|�����c�����3��>�?��o~�����ŒE��i�4���@��d�����%78֢�2w�w���ێ�>��o�����ع!O��f�eï@[$_Բ�����*�Ӷ0�U~͚o�;ù���m��Cd�&�W�B�������sҺb\CV����n|�}����ދO��hhH��5�q�=?�Ï?�����9�E�����:���K-�(�B+p1f���[l��^�(���`��bM2��cUȵ�^�еu�t�c�	%9��҂=jD�,4!K��|�F����Z�Q.�	iV7E/VR@+���ύ痘��	H;�z��W7�����Y���V�R�n�Dʄ�+��צ_� �CC�n��x��EN�����(5)�D"�,��<:��3e��ptz��{�
�jQH����/������r">���޻�_����|N>�$����q�]wa�[�`ޜ�r�{s�[I��.�M�H\�Ä9S��~+�=�<����m��J�a�2Q��:���y������jPؿK�|�D�}x";ـ�m{Zz�g@_��X�h�ͽ#B�"���׏�r���ܪ<�����@}s=��[o���5\pΙ�eTU���[:�?����)�^���sb��@ʅ�:"�j~��6��G���3^S�Y���Ϩ���Qx�N	w���{�{q��G����x,�T��b�8i�?�F�,K	7�@��[UZZf�x>��bC���K��D!-��AC$!R��o<�O/�D=�O��ރ���?��Zȉ�G!$v���g��sߑ�_ÛtQ�f�/�صpƌ���uc�������s���)4r�h<���*wj�fs�*L�<S<�{�s�Ʒ/8;�ho�,*����I8���q����'���nԳ�{Qd�"C��tCz2�{��@p/xG�k�G_�V�z����+ky�qū�BE�ubx��N;��b-���vY�����\��j���B#�U�XS�x.���X�x!����8��/��G���|MGO7�z/���6T�LFU��T55`�X7�*BSЊnk�F����PFD:�*C�L�b��lE�W���d��f�
t�oE˸&�J�9-$��{{e�C��nL)�:$%�l�E���и�G �.GH`֫ދ�tvB��n`d»%�$�F�Ɓ��g�y&~�����?/�˲�=�,u�����n��BW�ˢ�ê���;�8�1��hl;;���[��I{q,�1:��hR݃6l��.�ulz%T(T��c��x�s18�S�8$��?�g�l<���ޥ�*/�K���1y�D�wϭ����p���~p��"�jR�T
}l�"�
AB���c�F�Yx���)�3�RvO	�x��3(1[&/���*����
�涎�yرmd��;�%��*|pԪ�T�l Chߺ3&�ᯏ>���ݏ�AQ[O���s��5X�}�4O��XM�x�0����QFGW�ƣiY*|R�V�ĠĔWB���5=(�'N�-:�z�$�R��F�Ύ���sϠ��>h�e����8�8��X|b�;b<b-��r����k���#��i*�.�n��=3}l?P��ǳY>� g5di h�n��1Z���Ip�`��j{L�S0Z��#����YT��g�t'~�8�������s��{��i1��L���S(+�@]u\
6S���ZQs6�<Z�}M�k�6uz�/x�ͷq�w.��� V�X��˖���?�5c&���X�l-��O�T���煍*��|`�Y���m;/�·����1Q!��+�ʴ�X�1��h�U�\G�4ץ����\b^�m"��F�yLM�ΎM���ܯ��O���0w�	R�Ea��>�Gj���?AF���텮�A�wRD-E�� ��i�U�m)�+!iN����Q���
U�<z(�I�U�='���҉�{�#�X��UX�bB�8Iy�� Z����蟔�����n�>��bjj��Ć!�~�%�U��ؐ��+�5VX)UP�͍��8�#���kf�2e�,H��H����Y�ǟ����&34�_P1�*�)���&�4.4��7�R�?��f������0Dp�e��8<�!��;_��PA����:��^@,��j$V�ֶ4�,_�K.�>N۸	�~&N���+�����{�+�������aG�??$TG�]�m�S�fH'K ���H7׈���%GFYt*��|�ݕ!#U�VRn���9�͎n��JhE�B)�L�8�i*���&b"���+��7�?�w1Sj�#7\��~q?~����9�<���h�oT�G�I���)P,K\�(A@-������5,E��3j�������4J��c��C��Y5)�b�Eh��B���.�m�ظd�u��NV-�"b#�I
�LJn��]bp���-��h<+m{��V�0���y&�*���:V4 ����7��i�&#���޲e���S��~�l�-��$Қ�g.�_�ם��+�+���Y �z��6}�\�J����c�)���sp�Q�GWw��+���}X�r�U5B�S�vu,y����~7�X���m���L�N�P���NoY�ۋq��'��h�1>,���4����qo/|��/n��j��x�С*����;��_>�Tc�'����n��Q�>-�3)4S^F�*`":�ٶ�!tF|��#�V��
�L|����q���_1��]��4E�Y�ld^f����_b�Z���ᡠ����္;2�#iI5��3g�����?��o並OI�l8>e�5�j����b)�����t ���b �L����nm%�.%��9fL$�&�q
�������gG�lS/{�����zL�ӴQ����Tw�x�y�Q���׬c�z�$G�P�{ɫPu��\*D�Qϡ*Q���"�['K�n���9~_����ܳ���-���������t3�����P>q�2*l�&�D�����*�
�M���S�e��0��+y)z	Ʈ�(erđKɹI�_�c$bR�g���Z�D�`ˉ��]�6�����!�IR�SI�t`�M8p��q��7a��feLr��Nb�n\|�wq��a��� V݌�5D��!�R \)���d5'��XK�) -5��J�U�$F�Uy$�eū�3�J�^2A�oG2y	��pu�Ԝ,.��'oT�#�v ��\���O���2�_|1>��ϡ��M&��U+��S��s��d��P�	�j�·�a�Hi1Q�[������C�իWJH�6�ݽ=A��jjӧOGmM=�y�9<����!9���Vh��:��y�>?�n���݉IӀĕ7H��t�J�l'�y�j���E)���J'�oCw�nqOQ�Ԁ\��Vu����6�X�
W\t�
�|��9����_�"���'�ӿ�T���j�L+�z�zc�#Z�V+�;Fe���;h]�"�<ʶSJc5
��=�b��a��059�����1�:w�st*��+�R�bW���@lF����Z�Z�f���n�j�ShU�e��WP���K���=�L���ѧ�A�2&����w�oO�G}�4x��g�b��F�C25j��0AtH�����2Q6\'F�Ԫ�@4�E5y.|_���ӅR����v���+;�LW�!ۋ1�cD���r�2Q�1��-��?�y��4�Z>��O����M��3����z��c��)�4�M&�v�m�0~Y�m`"����HpC��a��b��B�f�����Dz�!��Ec=���*bp�)�׿~����ᩧ��gK��~��@�������k�2C�S�H�>��swهz)?��!+E3�u2�@����9��g�$���P�(.=�h�y�)�0�-bƬ=��?_�W�:���^���7Q[W����'�|�=���"�l¸�3������s�THƣ�\�x���(��qBь�M��������>P�"m�z��ط��.�W�&^%5eѸ;4�ٵ�:y� �\y����G���K+S�YX�U�xu�Ģ 1EnrC��V�h��E��GUlg�q���c8�K��������\��a�Mm*�C��|D���`�>].5It_��P?�Ӎ�����$_�+�bX�M��J��n�Y����s�wJ��	7NH����������r�c&�b�_�iE��2s_�A�?�|̚5K��@sscp�,MԶ�,�B��%����0�*��ﷸ�(�B�5$v]?���k�ţF��h���K��Pn����x(6�|�}��$�\��[���52-��oo���ip��E�q!w� g+�it�1�����`Vy3)*����,^VZy��A���q����΅���=O��1rGp�Y_Acm�����#��OPS��	q�UU5B�'�br6���tǈd��6`�\Q:�B%O�h���v���c��uKaF��k������K��
[דTe�=;���2F=���n4զ�Elm�G�0��KaڄF�q۵����d"������{q߯~�����l�ҁ�-[���&-'��^�`[���~`���� "�6��H�P�#KE�0W����*��Qw*f��R�' ��凈��i�e{�}-����O��9�;
Ҙ�obC�PbH�C��ӧ�3ܞy�9���,�liǪUk�j�Y�{{���*�O�y�
2N91��Iʰ�?y^�!�wcsS���T��={7L�:��#�	p�M��Y����c	�H���E��"�hi��zY~�heU6n�e~Fڝ�{����oذ��OD~Jcu�+�M$#d�Kֆ���k+b���q�3w.ڷn���S�g?�i��֛x���u-�
�}ɕ�2{O�Jb���*���q���k���l��F�D�w�Y��^I�̚�tQ8�7��_��8j<�i�v�A�6�����0��<�>�gMMS�TfT��ڼ����4�
�j��}�s�����+0o���=ЭR5��_��n������>�V���Ő$�`'@&|�p��x:w��EJ���}�3X��"<��29��m��\rG�N^��s�cO�kX����̄p`�mn��Ĵ����8q���!�1y�$�W5�m�|��^����~����)S&�^ȪU+�	��9�mʝ�l[�9�#�MJ!�w��z۬��w���`Oo�q��o����׿��V��3a�$���gȗ��4�-��}�ײ|�r�<��9�;[h�^%0m�8�jq��ٳg)m��d�D��	6�Vc�]$��P�4MbP���VR�j��v#�kM��;��·��s�Acu�{j>���O�Z-zg|�<$�[0g��X����C�V�&�,����έ/%�� 6���u� *@տ� ��iU���:!�jG �56�\�)�8�_�\��}jpMk����K����s��ܙ��������g���[�����G&��r=��f22���jDK�����;�[Ѡ<W=��^Ħ5k�_'|PZ4,Y�X$������1a�R�D��q�KFĦem�W]K�
{|vr�8'�B���d�qe{P�ƕ�߳��{���O<�/^$@lKK������>/�1{G��N��h%�y��?R�-{6�֞��!bd���0�˔���\����G���_��R�D ���x�zL�-X�bE@��G�Xώ�h��s����=���~<O��� �`��B��KWa��7�"�'��Cy��>�j��c�Q��܊?��Q,|�m\Օ�=c&^�E|��O?�S�r�/y��f(�T60d�4q=���t")FJ�'��h{��ق��c0d�A	���4{>�|��JR(�>2b�CTޕ��?}-�RR�ͦ�5,�J�P&]ӌ�_3[�p������9P�{n/�����5��=�q��OM��E]K�0yt��	�E��G��'��+��	��k;���,y����/��O��|���.�����.�+�d2�դ�G<�8���X�X�����[�	���������־.'S)j	R�*W���9'���	��1�`B�Y��E:U-X�&���0��>�v���y����k�����,�4C������g=�iӦ�!;��Ce��АXF��?���x��'#�T8�!���0�=o�,2�q�HٿI�������\p�������tU"�Zjp܇���+1��ױq�V$Si�כ=o,_�}�r|��_ı>��9����~�c|⿿�kV`Ҵ}�CN0<�eu�0��˽��I�� ��s�]硸��/i��	`Xؒ�����И��
m���0�5�q�*u�q�xk�B����>�f��3���,�y��>�l�D�n<
�w���RW���vA��ް�!1G5)�ɴz�q��lEsCZ-H���/}�4|��?���N�s�W����F����U�U&��:n�{��s��P)�%LaSϭKn+v��i[R�I_�&'(��X߮�LTW [:���\�ӉȄa��I"=}_��C��Q�a��z�^�&��dRL��xL�+�_@j-�XO��KĜ�v�;��PȺ�B2��Sd�2��*C�W|G���Nõ�^+��u�]b�x�=�������WFCi��d:q����g����%�P��&=/���H�M���8�V��L��;^��k�����?��=u�l��µ�މ�q��C�������ُ��w.�!�x�5L�:-��X�v��Jp��}����9�摝2�Sh��6�N��X
�]iPke4O�y7&ul�9I��PGp���ɛ�yX��M|�}��ݷ]�@\W���z�-���o�k��V�9�C�ƀZ�8�:���7Q�\�!��Y�V�b�����P�uo@R��+.���=�?�~�����SO���Qh�ڕ�ɱ8�,Uy87(�]�Zrgn��#C��4&m��å�|΂����d �B���e'F���ɕNW���y��cK��/� ��v�u�N�C\;�}����6����X�����"�|��i���5�����_�������"`�F��'�e�Zu{��R��a��œ/�ܸOX�M�L��?g1'	)]Wx+�*���
HU�Ч�T���xN����{��8�����O~��~'��G�IVP�t�o�i_;W^�-|���d�<e~z��8��+��?�Sf��x�	���ň��1����`(�ێB;�s�+1}�El;���1�G���k^JYǾ~���N<O�Ț{׆"G�,G�:���X� ���q������|�_M��~�����џO��u��F��T�#[PPT�Ԅ��Q\X��͓n�r�3�����X�C����{�^����G��Gk[�(��Uй��3��lo)�Wv�����6��fCN�44(6��x\@˸�<������PDڀn���yD��-f`� ������)W!::T�+Ad�0��*HRֻ�S�a|�n�u�mP�PN��#b:��)�bc-z����{�%��ᬳΒ��x�pڐ��E��"N��(��[�S�Y�N<;����wt�. ������w�"R<�#��Mط���L�\à��I�{ṧ��K.�.^�%���g$繶�u�u�Tx|��X�?�(���g����⺫/��u�����0g������	z����l�O�Vh�$-_�Ro#��\��$`il�ג�w��Z��ۗG��چ�Lv����w�@ 8������y�m-M�ڴ^�H1,[� '}.��\*��ދq�&��[~����_��j��%����;6�;���S=��G��G`��R�eX8-�:�d�s�9X�V�3��U�]�S�N��ԡ�0ż��/��s$\*��At��Ճ�h�ڊ[�~vEe��Q
�"�R��A,������z�6��P�a0\lhAK��j��Շ�%*���Jz��6*ao&�t-�<FyשTRa�Ca8�h�b��lh6i��bY<���´؊5j�ӣqa��{O�I�Ʀ創���\�3L����#JWc��q�S�Lq}!�� ����}�!���K�m�\z���2�MX�~=�j��=��e߽Fd@�>�P���|��������S��Q�2QyU]R�ا6����/	]w�R��i$9*�~ƒ�Snx~(_�J�w]�t���e�xV�<<`�у�2h�I	$GdG6=R^����t�c��X�8��C�#�0�����J�7��[����s��4��a����LE��*��2*l�RK��H+
+�lU+Dy��8�+_���/����cT!��ݦbͺ5�}�}�A���(ؒ�>�E�UKU;��z�p�$��g�,�b�[�M�$-6(v#�;|���k*y��g8�j7�q�(�L����IL�@�ل.�x�%�#,6ạRT�+<_�w�o����d�,�F���()��z)Wb4�7mD�=�ZV�gޓ��ǜ<y��#���%z9<>q%b!���������h��H�y4.d���e����)A\���#Q!H��)���j�e�:�<�ǵ�y��Wa�ve|tMQ��iX�|�Z��V��0N<�XέQ�S��f�~�yX�a�̜�-�=zA���f(�L�o��n(�YT�2h���`DL�r���T��j���ʷ��F�3��Й�䡼��}֑P��n\mUB&}cU_|V��\���G�~���c���܎�qS��U��H�q�օ� ��ܞx��ZeTL<8Ѓ���S�r*���?��p.����ǟ��i��8Ѡ(WN��L���4�czyѾ��;qK-�w��Q�`e:�F��	7��c64��T����W����V��ތ|fe���a���z�9F��Cr�Hc�xa�2D����ʌ��v&g�������~ѫ�GQ�J���[��=��Ցa:�� ��؆�3R/e90Vt�)kX�5��P����W�̜9uj��hGf�_��f&s:桦:����jLvK��s_�����x��Qǈ)�8w���z�۸�ʫ�9����e��~�1������/~k�/Fs�D����Y̗�g0[�5VŲf��{V�S6�"����~S|Ǎ�w]�1��wv���v6oĿ+WV1Pʐ$�\�ذtv�ކk�w)����w�e|+���?q�E�!U�,�bT�g�j�
�dL�>$<[w�`�B:� �߉�58��_Ƭ���~��~�cqy�N���j Q�4.ujS�x�w ��
}���s���)Ki*�j���q-�!���1�G�Ǣ�mB� �I���3�rWM{Ԓ�Q��,�4p��4�=j�Q�/-�C\~^������N�gd�ڔ���9)���jN�[�'��A`�	�ѵ�)��R���p��/Ƃx�%�;a>z_��j/&��h-a^F"��*���jA�g�6q�x4K�.����{����e�غy3�� �k���=�b��l�ҡ��)��c#�������G��������o�!.����z�*L�mwi�n�A�Y3�mj�$�a�JEJ7"Q� lwn�G �J�$��;��H-r����Y�oX���~��1cj6m���)mx�O��+�FƋ��u������SH����`)}��r���0<����58���P�tp����g�AcS=Z�M�Ǧ���f%v�NW���y%��҈��4^A(�5j�r��k�}�	oWq��Z�$|_�r���x(a���Y�Qe&��0�1>��Y�X�"Ɩc����Ņ���o���-l8�w�`�a�KP���f���k��"{�0�Ǟ��'V���+j��H�Kjh�Ǧ�i 5Kz�D<*�M�P��h��l�i���پ@�Jh^���vL?��{ �mMR$���[y�>&Ϙ��+W�K��
����śo�����y������V�-S@�k>g{=��*=��<��k�vg�Ds��$�ۅic>��k����²��]�1�8ŋ'57�w�J4T��]�9���ڃ��z��t���V���h?[6m�ٛ�Z-zT,���Q�����AR�C2RĜ�S�O|9
]~���r�:���fUܫ��Ne�Ȳ�_$*�p~H��lޥ�M<�T�WY5 ���R+XKK�T�S��N;�km�lvB�C�  ��mQx09��ƲO�DܞA��e�Fx"��Ó4��-w�~oe�^���,P�qmV����u�G\����FdJ��6��˲e����My��,Ş��F�j��mr�y1���M�6��ai���QJ��U��7���#�
�4=^?��T���Hإ��lي��3���[�a�X�>5V7�Eo\�4�n݂��&��<�6}�y�o8���p�����.�.���$$�x�/zD�
�g�AX'��p�����޶��Tm\NL-�N"��u}y����N��ܒ)4M�Q�� X�I�� ���"��y�N;Ft�+?ÓuM���a�"����p��3�aSZ�7���[q�������	3�O�T�FĢ�U�2q�l�4��Zij�R?�5*�U[#���ӐN�p�7�Ǻ���K<^�� �G�$��<���6צ������I+CBw�uB�r}딡1:"�,�'ZB䊔M>kL�����T�}��-�w����ЂN!P���9�Q�M�[o!̏a�o؋�G	H�Kx�?���r�z���P�Rb��=[�Cπ��aO_�n���S�pY�_O ���g߳,d˻���;��C�@|��jr_f��Ѵ�w�z!O:F���&���J�ȹ�����{0C�%�^�{6�cִ�X���s:�T��{���8��p�uWa�����O������C�k�,�� =AZ_�qF�@�Z�[lRD�WAሑ�iԦ<T�����]�z_��ϒ�<Y�0��q Rw5���i_�ř%B�)R�Y6$F�-�G��(�cJS������N��N� �b�Mc���s�Ux{U��&��x$�I�O�3�]�:�G����8���f�vm�a����u<��c����P�V�^_RuRb�-H�i�"�X�2�м��P'Mz<]ipyy# ]��	(�+*^aڼL6�i��B݈����<w��A-2��ryü�|�T%��f��dc]m�`E�X�:tK�a���H�d �i�JM.�b��cEE���,���}��ԋ��k�-K�F���;��ic��c'�D��ɨ�+�Pk�R Jy5y�>ڰ�N��I�$Y)����5l����RUϏ?�����hnl��ի�٭�8�1��tnQy��u�a���q�'��������󔐬����"��U˖��u͵u�֧�q�2V�|�fL�
eTι�2�u���\��X��_�d�'��O��'s�|}�?�E��uF�J�4=8�dT��Z�ڶ��5cP����a@ilr��)��QD�Ͷ�AY�M���-�:$��w�YI=ݭ��x)�n��0�-{פ�`��Ck={��⭗�ũ��.����ѓ�G$Y��_�=<������ii�_��8�m�hō�ZS1�D��Q���~��#�<?��}��f�r;�o�~��]=��+w3�?��3c3d��8���}��r�v���ܒ�&�x!6�q#���'�}CS�i����O,鍓��&�������m!�%�q���wuw(�*��2.sb�C��,Rس�ބ>>3'���}�����IS��a��5r�x܁������ejU��"?����@B�=b��1���$��f���&E���a��C0��K��Z�Rߠ�+m���9X�q��Jr��i�L6���7�ʇ~8^|�%���<�:4�e��I�X��q�L�X�kձ�M���k�����\w�Z�Ʃ��U\t�7���E�<s/���U��_Ђ`�xu0M�"��F
n ����0���
������Wn#��)�	||W�ÎT��um��u*����I+C�Ŗ������~5�q�B�,�/�|�1�;�=��fj�֚v�Sވ�[���ˢL�j5��9h?��}�z�/�޻�D��|5�u�f[5�A�T��`�eKL�� ��+�M5��!삇392:��el��X}#Iq����0�R��� ]+��s�=���dqԀ��4��X�kP��A�?Ca���LVD�C�+!�W0lM��>z��D�dc���4>�`x�{p饗K�(Y��\uϠd`@��^l޲I�j��Fb`Ȱ_5^�L�sl��h,�T�%+��O��@;x.��,�AC��X��Z���6^��Y�J���!N���#�b+����IH�/��m\�V��mS�a\S�܃��7a���X�`������3�@Vy@,F���p�������&�@V}�CyL��gaƇc�b�	�|��	�3����@��_���.�)����M�ñ��U�f\�b&����B7���{a��Eg���%gU���o�!��W\�d*��~eh���?�_��{��㽢eM�����	57�2g�{���#����F��l1z�A�����<�GLl� ���9�R�-2#�?�e���T�J�� I8.����1�P��y!�!�5F�}4�BcS�Ҕ���l8{�������~]��IF���#VAb� ��+�g�����"���>�Ƞ�����0����� 6kBτZ��r��9ꨣ�5
<�]�Z8 ���S��J	�:���q�7k�9�Ԧ�v,��� ���>X�+���:YƜ\	ߴ���ǥ��9�O�<I����)�����BS'�.Ӄ�YA+�_I����"�2���W��xnܰC����+�����8���㎻��˷�y�|�y��}/\����+g������mlFM*!F,�L����.�����C��g �aln�8�;ՠDH���c�ـ�O�XyH�޶��a�u���=�6t�d�"�ED�����ڍ�\w�5�=k��ʘ���ŕ?�mSvC&�#��2�HO�O�H�T�B������1>��CѥB�^�,_�XR�9�&��,M:�VN��5NNBN���wN��U��$�~J9۴�F��'�>�@VQ�^B��В���پ:֨xҔ�*nݪ[gR���o���r1}�L��a�����Oeʔ��s[�����ȆAdN$ݝ/�E��a�� ��8y�����ǬY�0�K�5��t�Of�J��/�ɞ{�y��	Nu+,��=',�B��۰��I1&���l�;y|�s*��^t!�n����u�ى��JЖ��W˸q�����>Ӹ�_�V�(����"�����(����\#�K5{J~�o� aˤ����p�u�Ļ��O|B��A�O�d����!�P/;���F��S��]|c��*�o�I�nf���ŻP���ľ���lj149BEl���\��M�d���C��ԃ������F���c���g�*�,-0c��\~%�O�^��~B�n��Z�WǔϫcR�(F}�TD����3p�կ�yZū�X%��� V?��chD\��	�
����ش�w���G6"��3�U��)\l[|��y����6�x�Vb�=s(�������:�n�ϟ�g�}V[�y�HkPyh�-e�y��"�-U�TV��>��o�Y&�~''[*��$�u5QI�[CL̂�"��:>3d�=��x��4��O��_�b�B���x��6�!)�ۊX��K���噇��N
9���JvK�,(\L
�<yM܇��F��ϴ��!�m��*��I?&O�1��4���H�Q^y��iR����O��Iq���S>*��W���s��ukW�o�x���7�2\�S�YR�F���H����o�,��{);�8P�o)Ў�|0���n��ۈ[�]���ܖ��ju�U�`}"�����bެ�8����nù��诽�v�z�_��eHRU6i6#{�����גDSu
	u�ښ�U?[6��Y_�
^���u�:�a�Ŏ�/��L�j����j�oQ�%��j�����~�u�H6�+տ譂ej=��<)�{r�н-3*R!�I�<1Np����Z� ��=cu��,h�15ɹ�vuu
����F����s�����4�k|���χ��tR4-A����&�&��\e�>)ΰBW��jٶ	�������
���vkl��5>�"��帧�-�K�AK^�n\6�[���>a�����*hi��/�S��Jr!>���^1̆1$����x�+C��H������Β�f	E�x�T�;e"O����3O�m�̙5k���MCm� �߿�Ғ�b��� ����xk����D��U�F�����3�J��o4�-$����r�S�u�T��)�iO>БVO}f��ؕ�a-ȣc�@+V��$R=�L~���#�{��3s��&O��7�u�9��6w�f<�S�LeԊJټ��:|N@Y��i��A]<�ݦODS]5~s�/����2Йf�gQ�|F�;Ӝ�,Zo�H٨���=��V=[)l=���-�r�O7ZvO*���b	e����v�sp�p�	�Sΐ�j���0'3W~N�N�^���� �Al1'$��U��-^dWh���ǣa���z{�|���2�6#e�������_�`�����':���>_?�#q�g+���xn<��x�j!o:W�4,���,Y���k���e�	!-����yS�ֆ��зa�z�X������6챈#ٙ���yQ��}�W�e�2V
k���d�z.}�j=��S�m�4�w�W�|�"����>N���H$��͕S4��Kx�h^�㔠�
��qweڸ��Fz{{c���"0�j.�@�c~�zI������h�EbE��l���͸�4^_�2n���kϩ*�@$��o��WeP���is0TP�U�BjR�x�H��H�z��&MBZY�)[ѫ&Ͻ�>(�Q6g6����X^�3�VvJ�:���dr�ρ�z��h�d��l��އ�P����HPVoC%���$�C�r;��Vޚt��RI��S8�w<af��50؇�Ns�Qx��W%�i�#��oz�(fuD�U�u�s��ze�PL7j�M����^ת��>r_��UۧGDG2z44GY��� ({��g㩧��t+C2~/C0{��-33��@Jb���p��שk~K�s�Y�K����V�l�\�<��p�d,��^�`k.|���3<�����@�=	_yM���Xy�y�ɸ>��[�C̺V,K��\MU5F��
��D�X����ŋ圉���p��;�7��'?��{�C޻?^x�Yy�q�����W�t�<����BZ��l�B}[�t���^z6���
ӝB3�K:+��6z��ۓ���5q�t��X��xİ�"q����e��~����g���O�4N8�(�tfd ��ڛ���7���
?R���R�M�5�e���8b�*lJ���Ԧ�KS�E�2a<}m>6�v�L'�M/bnv���~��d�̙�:NB2��
����+�N���`�lp��6�`�Bl@2 �1饜6d/��<7z4v�g���㏋^?��#����_�7[[# ?x�D�����ġj�u�ËG����?�IB$j������i������6�����e(�H59�,¥
�H�<�@�1���ı�#���?��G}��� o��&.��
e\��7�$����bϟ��{(�_��e�1�����F��#~DBazR܎8�}r<����/	�(��Yrk��@?uwSi�#^�%�kqb�X�b�ҥ�k�j�6s:,�O��;��-�=|��'q��G�����W��u���":=&M��$^^13�,�������8o׆<�k:�c[ڷ�@��<iV����<䆀�zͭR����m��i�$c���fӅ������^���P��La��ufpH��R*��f��XS�b�ie��L�O����+,[�Xt9�w j��B��dFA���FWꌩ��s8���^J�Wj��)�eFǱ�5���GeZ6;a�q�r��2!~��{���-^�	��Lr��S��J'��TiO$E磿��{�r��	�"^��l����a�>�G�P��Nn\�t�����C-��A��⩒^>L��mhh��������A�ƞ�G��()��N�X6p�!c(FD���� �v��um?��,��[__����	����_����Y"yN�m��°�H[�D�ƍ(w�<C�oX��K/�!u�Q�D8f���k�����3�j@e<���dˮA�Tx/��|�q�q��s!�1U�e�y��g�y�g�Me��Ad�����\�����%3v����O|F-���#�5XP�]%R�B�c�iZ4D��!q�E=r�I�pw�A	�k!&� �����^�,�bA[|^�4�V��Ul�I�cp�:����~���ZlP�ƴ����?��+�aڼ�1@͌�Vg�%eͽ� �"=�,��_:��m-��s�<��?b��E�*%e�x��6d�
�v44ta	�6�LN�+X#ya/����P���+d��Jϕ9� �K/���ȍ�!��;�S��WK+�����F��Mss�Y�����֞-�aV����%�c67�`�{��������������{��;e��9t)�TPD����|1&���X���Gb%bE@@$H�a
L�黷U���~׻�^{H�5g޹�5{������r%pJ�"����+���qeȆ`m�Y��;��N�b��_n��&]m��=~cETMl�,k����X��hq�2���r�i�}�����S�ICc�
',�#���GL̈�K��u��D["@�0�B�6Y�UΜWѯ�Y7��ݪ+ed�6zYE�R����l��b��@{��h�./[7o��[�'��X��ߣ�?޹����A�;g�\����ur�K���_��Od��9��q�;��p7x�L	��.�ѽ�%
A�HZ(��-�R��IX���0r�p��9)I_��!��H��$�y�t\{��\�Y���|��ګ4%8~�y��M�U:�g�ds��{ e�n�8!��,�����8��Sf9�r��˃�'��\!��:���8�Y��	�{K�y?����93�����x&0E�&*{q��ǟT#��4kXx%Q��j3�1������Pa1S[t�k��>���eѢE���U�a�&=.�J[[�n@�9�R�.�+����t�R?7�y�����I6h��ܕ����筹:�/~�=�5k��o�Zz�9�M~`�w<D�����]�1��r�X�ب|�r˧�s_���<w��(���4i�B{��SO=�m����X^��=�����B%������wml��j��W�>>����E'���<K	�y�M��<XL�wfO�Fs]��QE�����ٳk�ls
�ɍ� k��}�|�{?��G/Rwn��W���	y��ge�=�1q�t�K��E����Eä��h�%�&�|�T�(}A�;��8��TS�Yr}�� uZr��=p��q�������~��g?&u�N��:0-7��q��4J��i2"4�S�g$yP��P�����_�h����&ɼ���W��#kW�p��Y����"�V,������1��ɒ%oWAf�uG����y��A�x	�im3ua銳�Eم�,46��`c���åy≥�(9�J�_��u��+җ��El^�E�LR�'�a5/����lZk��Ui���G����������bHw TR\��y�O^|��Ѝ*�h�Nk�ͲA��4��	�$����+օ��r��Ν5k�Z$�?%'W_�n��g?������kҷ�B>��`1N_�c�������D���Rz�e��G�)���N;M��68{��	�����P$��¼��Ik&j$����w�ּ�B�>�x3��m�㝵�_��a��_|Av����Q��r���z�Œ�8�N���p�,�g�^����a�/�P=B0Le��$��ػFC#�n�NՊT,�Y���.]���_��2�ٵ�M�0y�|��_��qӧ�HXY�$�Q�5)Px6$��IimH�'L�8u�����i�v��sE��	��j�.��BV�׍��4^�=�l9��-���W�n��/S7��Ft`CW#n�T�e}QX!L���X�߶�#qo��F�P��,"�'� 6���u�L��lzsk�,jp�M1�yM���<��A'�{z�t�!���_���R�Y�>V��c�e�A(� �0͂aS�zq��i�f��� ����d���q�R���5��vA�2.�+��SV�~]ǀqZ�x�c��:�����G�K�-[���>���Z�ӳRA��S����E>W]u��#.�bGBh ���TRN��L$�14��'#W��qQ��XaG[����m��NBS��ؠq��� ��ħ(!����#;�o���]$��|��X�Z�ƣx\�̝!��������r��K���)O=�Lҭ0���Uc(��R�{%����	��W����RR4Jm��C�םP
��R�7`V���ǔP�$1A��|-f�}2y��YG��{�9��S�7ا
��������$�k�!L^&����\AyM��=�N��3X�v��Y2o�LY���겗��7�d}��j�rA�|p+�Ō%����w_%S&Ғ�]'W��K������vy��r�����n�ݽ����HM���~�|����D&jA�.���Z���Vk���gc�a��p-���\���>��3
σ&G�Ι3O�a,��K�X�$h��@,��sr���o��n B��y�e��P���?��ү�����K(����tr�w�������/�m�vȼy��[�Ly��qO�w�����&���A=������5���	6��b>@���߫`���� ��$��U�e���*ۯ��O.��?x@rnn:�y�I2���OL����g:���tV;�rω���u��UA����{e��7e֜�~=䲒tk�{�k����^�F������k?$�����}�j�!��D��+�PI��4�=�$��e�.�tų`w׀k�/��rv@P��Yga�Eq�څ��wIi耴C�?�Uڝt����۾��2\��Vg��8S͓��E �3�����,�`Zܢ���ҥ�(�M�g��s�ź�\�/� ���t���~/l8��;v����k�����)o@��@IR5�TP11D�&m-�^�:�C�7�^�6pN���������r��r�3q�>�U�2��^p)X#|�h�j&!�چq����[��:��C��(yM[n\�A�:k����XNÃn��Sr�q\�xY�����s/jR*��she��D��_�4
~â�{�� 2H�c�m�꿓����U�y����Pf��ٴ�]���ҧ���J�!7Ϥ��HW;�\�W��$�#7}T^{�5ɻy������}��z�O:����"�%@�Y\�M��� ��@ ��RN��F�^��%�r
��(#咊�3ˣ����I�&sa�P�C����&b	ٽg�����*0/��B�^����4~�䔀�����b�"G��#Ç˽~��]j�cΖ��P���Z'$���;�ӟ����G>|������_���hnrs��Vw?Cn�$3΅C/C�;7�ɂL�s�J� ��"I9�qx]j����'}g?]h��O��J����E�T���Aٳ}�|�+��:�����u�7�My���dܔ9nQ��l{x���m2;��d�O�t�a�ĩ��|��N����S���{�hxPS���
N�:�����_,_��u�	޽��n_�;R����PBE���U�@C�En�fw�k#X%A�*1�΅�#��.Ԑ[L.�c�k�Խ�V������W�c��N$�������/�ABjP�H43�8���[ezE�Ϣ�G�Qp��c��rӷ�0M��cĳ�����³?��R}�:$V�sֳ��:��R*F�#���Q�φ��g?��t���s��hP��-E, b;��mw�:Xz��)
m�ơ��,-���mɌ�f�³^8>��KO��@�V���7o���cV�e���jE7�뮔J���h�gް�dg��%����V˙��,�eæ�J�pϯ�<]N?�tg�>%���Ge��u�Գ�H�����{y�7u#��#����1%�aA%7B�Ж��<w�-.n��\�	�C�t�/�?��?��'?~���ץe���o~+u-�$�&7�7�057��`�*�i�i���M�c�<�u/u�IHk���[�"&����� ����GА�����\;Th��E"]1������\6�n�R���ґ�Gv�L��0���G���� G�CW�.��9p#X|�?�W��&P�J�E�&���w�����{�7mI7'״g��p1Z�`Lc���+hkB3(!���\p�Z��(�ɳ{�Z!H�󛜱 ��ܡ���i>�S8��#p/�۸�?��_�O��$r��sϓ��d���jq��w��h(�|�-���׷�����zp3Z`����Y�4�uuy�,��^zA���%w���o�GdYz���R� IFR{77��y�~j��z��2�Y�[�l�p÷����׾�eԠ��{����ÏI���j1'��0n�Ҍ�	�$��e�L�}A	��@����6�1]�˰����Z2mki�\O�3�Ҳu�V��-��Y�&IWw�Ի���?��bRfϘ-}CE-pb��
� a�4�a����㏖�''?����2a�D](0����;00��}�B^MI������+Qh�ƍ�%y���1��G�xJAK���b��a�&V���D��km8�U����`�p$��{�u݆_�b�
�={��E�^~�媁I/+�]���T�� f?�����>�ʡ���i�b.�lL<FRK������?W,��Ã�PLM�_b�4o�j���!�%����X|橧��'�xB�پ�8Z��H�?��ȏ~�#u���k�\<?�M��9�~�Z~�U*�qX��I�_�.�D�:�ie܃�FЪ��}q�T]�������iY���y�!�ͨ4�-(F�g�q�
�Ӝ��T�������|�U��+_��["W]q�<��3�:n���N��[� �ĭ�EaAj��X�tyt �"~��B-�&��-X(	�I���n���,[�.���g��?v���lji��W��_���s��E%��:?��ř�ݒpB��<i�c/^t�\}���_�>$+^[&Ӝ���u $!N�2�B������{��s�.���/��/��Pm!f,Z���U���
��{rKCƤ�L�� K9:��0�
�v�M7��j��L`l��:�B�5A�碎�sY��,������5w��b��8c�mL3�����>{B��d*�ӱ�'��<�w$c+#�x���t��|��,.ϡ���Ca���0��CP�z������Zr;w8����^��)g��v��<��c�]�m�}aU��g�YJ7�Ho�c筏�j�p�VЈ�ĸ�e����wP�_��+��i�se�Zv ����Sa��#��Xjna¶_Ĳw��q�*c5k�L}o�s@�^�'�R����6����٧d�3�Hp�U�sE/,�q�,F��t�\��<�P &@ٿ���sʪ7V,���+�}�I�uq�?P������|�#�����J���;�!����
�"�!h-�QHgS���h��!��햻~��Ѫ��,k�D4+S�F[YET2������"�`#�}`3-�8��6�n�dH�T��ϧSe�,�E�Ba���Kji�0��5��0�����K/U7������,H�fd��;���2!�L�K� �sȎ�w�P/�p謞�������b�͉W�Z��m��Xp҄���I�u�Qp��fE��.-�N��k����xx���IǝX��{�lR;7��c,q}�\A�;��c��od��:s�u윏��'�xJ���Ǹ2��#Ӫg��p�H�sg�q�Z�(��o�ݭ�U!����������y�t��5��Ύ6ٱm��5�(	v�[�����Q����7� k7l�s.X"�}�j��'w��i�( Oa�����)s%�h��C�U��A"�R�����#�F3�0!U�մ���$>鸣���iٽ2����Gz�	�2Wz�p!=H�C���}�%4��QNv�I������8S�J�F���`;AE?ے����ի�t��g9��݄�s�>ݸ>7U�F���N�����QX;1-��ڬ�z��w���Dh 0�-�/kׯSBp1d�u�C�<�qIj�\�ϻ�3o�.h0�!4��z.,"�m�w�Pip�Q��	�>���	"�ƙϰ <�ߴ���R)��PA�25+]���Z2뗏c����5B����ⴣ����{��$���`9����<5 ��>ZT#�y�1��Z�n�k~�a'8:U Y����1(�����[�k�z׻ԝ�җ�䫏E4��Bࢋ.T���qo�Fu�B���Yl���#��Eh�}}h58��	��v �'�x�u��e]9�]������t���%�0<䔇���&*�i����s�+�&�P��Z��>��Tc��;�����$)���T����BV���q�ے�Q~����tA�Yp>l�=�-���nz���0w��G���od��Yn�:�br�����������867�dʄN��ÿ�V�A\fRZ��ޏo�|X��_��i��nc�ָ	�[�e�p�*N͸�������9Z	x��~�3_aq�ǟ���߸A�x>�ˢ)�����r�X���cA�)�_b!L~�fe��7��
�,Οc;hQ���d����:U6^����?o����yeܷLP�!��"��c��\"��դ|+����1ՙ���S����݊�)�K�� �����5����;���x��n� R�*d^��y# ��o�&���'��?�i�/�q���ޣ.P��AH͛;W�;�<Y���Z�8��@��v�ĳN�燔r �uΜ�r`�����{�|�Ə��u�+.����J���I[c��h�s�0���a5h�zW�U�3r�%�Y���:3�Lޙ���"=�t�����2y\�\r�`�܆k�����lڶKf�X�;��J��0�4u�Y���m�OI:A�SV������F�jLR��78�R�l��X�Μ����Or��[^z��h���-b�Lb׸KcG���g5Ⱥ���T'�H%)�К�$ A�TC����6��mX��I�(����(mCkV*䫵ఽ�������s٦�X�$.,����Ȗi��������Ÿp�������^� 3,�UʇAaI�DA%}��Yn�(����4���*���w��;������\-�#���/|^�?�8y��?��'�T��|q�~Ƴ��B��q,���.w���-J�q��<Z�{}�I'ɝw�8�&�>D��w�,Ы{�]o�s�������9������Kh�c�@���τZ�%p6`}XO�˻q�b��ۚe�]r���w�in�w��w�����"5ne�)�*�E�H���Ĉ������[v��7ܦ*:���A7�<��Cr�?}M�L�Q�-���~�kim� ��9mn��|�3���rԌ�2н��n�=x@ڜk��P��9Aљ����$��	z�E�hJ�_�+��l��n���9��8����bU�_�R�1�=_T�$���P�l�:h/*[�gN��X��{��sm4�((b�j��瞋4�	DsG,+U+u�{�rob{}�g����(�,��x�$��ݛYf�X�X��j�S}�kT_�>��e~�����p������z���sh��0�g�j�E����yx��c�Lw��!@�	a��Z����:�jm�����@�gm�J!� �%&x)@�(���z��&羸�3g)0/H��X�����ʇ�����O��/+.�3�qV����OK������ܥ�Ʋ�D�Z7%xƂ�s�,ψ�j$l���������O�d�ʀ��t��N�y��������
Y�q�L_�H���Zj��9���)E[��t�묛}22Ы�7*�qA�H���׫C\�X�gn��\w��`��WW��]�uw�]Ο4���%�.p��`��s~��1���È���������UB�E��_���B��$���?><Z����!�z���V�Il�e�b�����6��X��n�R��'z-��+R�~�̀�F6����8hi��׬N'�Ls��Z�%Χ
��c�L�Zp���uu�蜵9Ko�U�=̼5;e�]��X��{�qd˘s\��K@��?��~��auR�~�)'���ŉ C�P}K�}6f��P�E� �x��s�vo?�il����6�Z�ʞbCܱY����5k5]�T��F+���Ν�����)�S+��_/��Z+��E�|@/�0�Ӑ�D�bG2���	aޣ�uq�i��B���:�h�����u�8�C�8k6l����d}�d�$Ce�3hg9UA�����D�3�q�%"W�&<YO���m��ԙr��n�M���]�u��(e��5Mi���i�Z�i3czG �����l���`��d�����c�P�5BQ��6!����V~of�6�:-k�5r�Ŵ��`G\8�-��g�1%�j��Ð�����k�����x���M�����?~�n��g���xp(>)D�F�\D��v��@f����׺��G4��g�&O���2п?d�V�'C�k^�|��_�f�'0��7����\'�6@��k�Ѿ?���t��F��k��o��o���Ϲŝ*Dqk�j��/��Mr���W�����%�_"�u����'�e|��k�����޷��-LDwPV]��5�
���q5�R�+7&��2Ι�)�oΚ1Y>��k���c���e�^�9�$9�CUp��&�Z�eΜ�Ҝ(J��؆=�U8�Ȼ�Nf�1x>u�J��$��ߕy�f�E\Tx6������+YL��T�۔��mz�w�� *�E���eѱ�(�{��߯B�eJz̀�̿���U���7���W}�R�l�b���(�VPI�d +,.���b>��qaT��)��:��SkC��0R#���jc��b/[w����}4�dH���-��=0�hzT���4u"�{<)��}	��|RS�������N�6E7�믿!���^�̘���?<�/����P�Q�z�����(iM�#Y%����Jm˖M�Q�+ÕW\�k�,%(�?����=�(��X�����K�3� �i��5Z�:��-,9]��!�I���#bY*�뱎�l+j�TI��1�\c�:�g%Q,hg���t���Y��e�	�����'?���	n�d�����
���))�5Wr}��]2���LԄ�r�&�x�Ӑ
R��NJ��[���ߦ���_i� 	2M�JqT���4�q�������L���P_�ÿ;t!��>��)"Ҳ@443zh@���eA�:�%�b�AXFo�W-�ʮT[1՟��-�&.���6��'����[����+�ǩ�Z_5��C�z�m����s���R��ߨt\��� ���T�;C0H��h,F���;o�>�z�Y}� ���p�i�^�ZB�P����$����J���M�5&B:���Y��/�������iӧj��N3�<�2��ٵc�����/��lؼEN?�$9���ѥ/Ȕ�s$[JEK��v���_�#��p$��&5��	g5�}��`Kc��h���>�a�{��)�Ǘ.��Ǟ.CY�H�u:؍h�a��S��ٺQ����i�*8(�2���49�v��=r�ssn���nr�ڲW�	�J�lZ�����T���LC|q��߰�_*�8&���po��S�����i�g������3��x��G�T�\�g}�ڂ�qq���(��{&�pqh;�n6:<���Z¶�f�Ƭ W�qlq	#�fl�9���)�3W�h��r̤:�l/'�O��w�3lL�kA�����U���+���N)���*R҂��BWo�=�\u�U�F��A���E���֯�s�9_+�qGʯX�Jڝ���f��Cb&�il�E\���F�B����N��t+V����G��C��k�Ȧ�[��)Jcs��<f���IB ��D��m�����z�y�f���0Vl�%Y��\����ڥ��9�qc%�)��4�{p�x`�9��o�93'H��n)���?�W�:���;	��
�����	-���Ğ�$?4"M�� [53�"��ýښ��W�W�`{���",��HV�vq��Ә���ڛ���wLZ���� �@72q׼�=�~�g���t���{������n��`�\����G�˄�5���L�y��`/���,��su�7���?o�gp��2ev>6��v��3g�֘ �E2���Q��B(�I�{`�\����9c	{���)#�c�qǄ�"s��\�MLR�!P��LAf68�#+�DvG�bW��,-J�ݢu/H�}�y��	�NJh("��,�`�g�y:�jk��\���K.��.�T�n�%���M]{�;X(d&K8ZKEл�q²^]�m[7�}��'����j�r9��䴓O�^]!���	�"[H�d��-��a���yΓB>��4>���$u���M>�Y;�퐋�������vy��u�l�&�~��2\t�Gc� �*Ȝ��2��N}�.*w�&!��V�#�@� `�_���ϔ�S�$N��7ֻ�4�ܴ��d���7�#�&�_��N�f����R! ����� ,�����������R����o|C�!;�����A>����ŋ�7��������p�ftoA�׈����s���0xeh)۠�@�UQ�P���_1�}x�k���1U.l_b�y/d|���΃W^y�lٺ���>�<�f�G�Ca0���m�ҥb�;Q���˜�A�RP��)H�3�<8
�c�Ay�hT��.�XXCT⪩O9\X�=80�da�-�*��+��L�= �P\�'߄���������e˖+��7R�׹I1�pI�x�)�mN_KIO��kk{�s�4I�u������{�y�<*N�)�`���H�JJMIC�����-�&N�g_|V����%�w�>#r�Yo�'�xuC���ۭ�LK�"p�'Pw�z�ۜ�H��`��$�2�6�u/a�rRrǦ�r�U��Gn�V;���}�u̓�'0z�e¤�rp�Niv�>Y�%��"o����ؿW
#�:���`�{N�O�/|���MN��6'�	p�~so�on�h�i�������\�31Ԥ�"AG��1�c�rm ����׾�5�䢋eά٪�z���	�%��6 ��pX*����yx�TƠ�Q.G��G���=C͍&���[�wuL$~�蜉��6�gˌ�(�'�1s��]�Z`���7w����T"�)-0���
�����3z!Zм��U�O��`�.�*L�Z�_|-?��AC���%��5i�o�N����WWx �2�v<f���]l�
c�.=�3�����
��̙����ղ�{�������;4q���e�_{#�Z������KΑ���ha��~�s��	�r=L��d� ��p6�>b8�R)[*����(@����� ܥ��L��h�e���I���W;�mݹG~��;5b�T{�03���	P�ե�'	 6~��W�0�\��3ϔ[o�USe;v�����2f�c���L56r��pF$J1_w�u�Êk�}  jh|@l,8,ȉ1SqÈ�`�[����^�q� �̅�pW���0:���N-��kw^�0m�7�.c>���8�/�/D�b�tl4��5M'��}Џ�bLX����W�7�C�����+��:~�PP�@6�sE����LX��4����qO��bm@#
��\^P�l|�G��y�q�}{V���C>.iu�� ��¸ro�o��&]��Ϸn�n
!;;Օ���\��������&��E���dٟ^��/{�"s~�}��>Q�]�DZQ�ܓp�dJɎ�����ڄ�j)��TT��lvH��':[�e�n��mk���Y�f�s�yҟ-z2��}��,���L�4CV._�%R"nFl���8Y}T&�k��Λ7Go͏�O	w�iS&5����Y�V����K��cC`�0�<$�Ҝ���=v�1#�C����uϊ@B�C=�B�x���!���Z�Ĩx�=O-Adߏ���¥Ԋ��:��d	o�븆��Vڍ2~��j�k��H�B.���Z���H�!H��{��_+�~��)F�S��g ��z����eN��QH�lp>�z����袋�[n��|��[���?ǳ��dhp$�Xn#�)3�|Pb$�rYSO<�T6q��o}�[�A�r�x|�}�������c�]$�],]n�y�i�/_�'���M2M�����{;%���r�0�a�˓	J�M*�I�ݙm�RN��&65Kﶍ��k�+K�~��EӲ}߈�s߃2e�'�:X�-�������yc�sZ��Ʉ�x�"}s&L���������P�W�Y�\��ʼ���à��� ��9�0�.O6�JV^��N�?���e��e�m).c�0�l���:`^6oܤ� Ƅt�w��='��;j�'�t�Wvxo�6t)�u/�e����O��=�x6'.x�B�q��Eq����&�����ј���e3z�R	�<6�XR����È�V6&(�504�,���}���J�����������g�x>\ �C�p�5����=��s�Bx⩥�z�:�x�G�l1
,�v46�'��B��-��<�2Ѱ4,h�5���5�V�ԧ?��Ms�}����N|����'T���{��r
񸣏�����sI���e"�z�[�\�8d��)$=e��)�n�9�));���%g�/�m)��K�Q���N8U����ztc]RrC�2�MP��?2��)*�o�[S��&�O����ߨ�	�1n��\>mV�	j�#m�ūx�G�N⣉���+�¡h�F+�5��9�h�*�	���:	n�Y�b���ll<���b�װZ������<�@�8��{q�J��a�|_�	Q/c|y�a�|��� �ԧB>R��[cn�jYUc=_��}K�VU��Ô�I;�͌�a4��;����=�!B������7�����&�2i���^��Q �R�!�p��-<��s�ů��Z����L����=���������nH��x�$Y��;ǹ�9�����#ӦL��:��λ�f%���F&�R�P��ѱ��|��Okqy�L,T�t�6�PɬiSd��)�]����oH"�(y	��c��_�餺H-)im����6�Ƞ��9���}N���*����Q{��t��V;wdc�)�X� �5`MB�p�hm��#-�9�="<B��qpw��p��d!�	&�6rrJ�l�͹ƍ��E�Ec��g$�m)O�?���j_n�e�j�rs��� n���<Q��X:َr���Z<	�w->Ÿ���ʁ���L�-nN�J��+�v��<������P]���<�-�1#���0�u�����ԄoDB��X+����3_t�%�#�h���Q*(����6����,����{�i���q3��Y���d���2��x��W�zi�u���&�O>�G��Y� �����u�7lki�M�֩�;�S4ny���w�CꝰI& ׅ������X��u�T�"� �9�'Y���}rˇ��E����18(w�ĩ��7Ua�wk��Qs�u2�'Cn`I-vtv()s��W��3z��),X 7�x����2��؊�L��ROJ�"�o�UA���3��h���6����{+�Ŭ/�#�Ⱦo�j�����2���`���2�zi�s�Oq4`Mg/�m�a:vÄ�	8��R��^O	K�g��vX���?(�Mޗ��q���1z����?9�ߩ��X��x�'CQ�xy��s�%�|1X��&0���kv܄IOQ��9����R�`:;2]F����N�,,�n�A����-B�s�%G�p�UZ��59�����w��xn�i�ޡ�T��%���f��r/�'��qJ>P?��jv�
��r�£�7�6��/-��^].�=U����M�n@�M�(S&vʶ���e�O�[���U�b� A&�N��C><}�T��غu�����[�*���߰A+\��b�B?�
"�A�����q�U������ղ��F��>��9̕�C��I�R.��G��'��ӻ��jb|�9m�DL��+���1"M��qN6>U��8tޞۀuf5����R�u� � !N�U��`B��~>���k��d->����R�E,Q1F5�f�2�c��.���ME08�;�B(�eh��B�lp jq?���� <	�G �臄 ���W�*�?���e|��LX�/��%�p|Z�4���UǊ��:X)�o&O���U+��+�4�d���%������k����JS]F��������ɭ_��9Q�u����^�%�gd��t"O��bV�Y0W��(��Dk6l�T�A[#*4;/�*	��7N|�=�O�W��'�d@��jp��3O�@�J���u�{�~u;*!�����T#��H>>l�����x QvkuaZ�6	�Ҥjn�d�MiHRV��zO58Z�y�"0�S�OK�E`�n�M^���zԞ���bG �cC3�'��� k`�`�t���^���`�ޛ�1��I���h�lt���L����'z�4��-[7&��h���AB�p�;�-s�X�x��
@c�S,��q��l�wAl����q�.Ec%#9-�L
Ř���I�����ݸz:P
�ܛo�Y�8XmR2̆�=z7�1l-���{���K���g�!}�:ιO�]dR��������$Iu�Ό�*,�¤�I���o���}Wɼ9�e�)�΍���OH[G�_P`R��G�dҸ6�2�]6�Y�>ۯ�9�P�`?~���lj��Yg.��S��0�ЗX�^����>��f�qX6G�k�>E�ہī�m���=��f'h&>��Dz!�˻g���퉏����T���7 j�*�S�0�>�N�4�m	��F���x��6���Z/Hi`N�u)�ԧ�&iձ5a����:�K�x_l�u���E�b~,������qךU�W'|>rp�4����8��U�j��~��o�m��*�7@v���!c��q�p7S��48�N�t)9615P���Y+�z�b��DbP��A(�}WA����p�	��:�����GF���@�����]{k�2ޣĸ.`��N?U���;Ze� l��H[[��5��#U�+�wm�&��DV���,>�$9��� �Z�C|P!��2��qxc(�\*�H� ��fe����no��O9I��d�^�I�z�y�>�x�JQ�<����NtRyPvl�,%��=H���7Y�+W.��a)�2v:��;����mQs�ȍ�R�\�	�>�������q� fb8��I�]���:���vX{��E���+��	����FyI6��"3�zh��<B�Z~�v�(��w;jt���<��Ԃ��<�(R���RƀT�v��K:�q�tqu6L�n�2��Z�
i�@�q"*P6F��)����?)��		cq
.�YԽI}{���&6h`J�������l�$��p0�6����︕\��x"�Ye��e#(�'�q�y΃%I���'*M�7��.�?y�������`����_k_t��2n@z���uB�,\����"�M���r���A���薆��L�2Qz�V��H!+��eM��fb�o���m"|�SN9�nA6m���u�C���⋊A���>bW�T���XԘD�,~��`X�3O9⾷	)#��P�v���J�P�ބ����X�>�L �g���:**L't1jL%)QJ܂�<'��,��X	<�E80���ު���������E� ��b�]�]�jY_�j��_9 [-_��ɕ�ߍ�S�����:��5J�����D(L);���H� �f
(�B� ����}��x}��ڹ[����ڦ�!fE�'��'����٭��ЪĢ���P�&���\6���G�xS�mCʪ�rغy��]�O&L���N,m��J�����0�x��Ŋ�W�t�B����t�Q��ʰs|$"j�X�:��8�m4�9z���\G�4��vp�����d�TZd�����U�>y��/P&^�pfw��t��B�xOw�x�[�H4<��Rh�t�wN�����>�46/e�>ݙ�oi)�:�5�5�[�,�x�@5�&��Zʰ,F¤wq2;�=���ď�,�Ֆ���0�8~|�B��:փƴ�Q-Z���!D��L���Iv��,
�v�3x��E6B(��.��ҵ�lyL�\�QVMa,�B�g�*�c�uu�=�^�,�͒��z��٬@,�~��I^��`�u1��n(k�7D�v�wxŘ�b(�3?�8d��`�}y��/���2���K��љTd�V%���}{�ʬ�f���{4����oѪ��Ҏp��Tҗ�'	\�|���@�\�wHKsR��Kϯ�e+W��)S�I*�7;K��c�������}��R���4����t����[>u�u�|��Ų ��i!_�/~�4km�=�,��ٵx����t�p�`Z�O�����4��-��mbs���i��wF-~���+��+�'Ű�~����{�~���|�@��'~7�.���,n�����5.����ԊX��{���N��/׶^5<��N���#fKa�et��B��A|.#��*��D�$���;�]`>	;�}qA�B��"�ߋ	�l�aF #f��;�����l�oЯ����N�,Ex�G�Y嚥E��>q�;4�������S�ۡY�>Zh�����Ep���ľ}t.���ϩ�B[S�vwo����E�2YWˉ��YiVw�ڮ��ǭ�cN[(�w���Օ��Vt��(� ���<�!U�nA����@��&�t~�-[帓O��^-�c�gL�&3�L��׮�gr�G���Io ���q��;U�N�0N>��ub>���|!��+n!��I�s���sN��4&�	6W�����i펑�f�)U�Z�k��5�1ի&�b%+o�C[+Q�2DԚp��X&_�����/7!j�m.�i�M��a�0��Q�����Y��1 F`B!EJ�,;�q�Z���R����Fgh|XT�x����M⸕j����Uu����Yw�����l�y�����hod'Xx~*��+6�S�T��5օkbH.���XғX�Q������=ٸ~���8�_�
�����ٚ��#�b{ɒ�4�C,������ߔ)���Úy����̓4�I��|��䢋�ʈ֓v��g�%O=��4�'�����(�T���\T��|e7@E� ���Ǎ�zgEL�4E}���v�h�N�@�ҵo���[hN�ΕFK������w���jf 
6m�-۶J[G�׾	��)��b���)-��*a��LD����Te"�~�L������ԍ@�i�A���ԅ�Л�t��
4���}������Ȓ;ܽ���EfV�� ������ǿ��
<?�[I�1�4�)ϯ2���w����y�h��0��S�&X"/���Ɣ�,x������;˄Nq���C$�����
��X�R� |)4��fH�|��X,��C��\��vL� 1amdM�X@=B�*�AQ�����I�]"R*�h)	ކq'��)�S�[c>�
.X=ԌY�ϔ�ٝ�?[-�W_��<��1y�5��DJ������d��蔤����2κ����F�r�xݺ5N ���N\��O��zĹ�'*�8�=���<D�%��Js����7�K.S���	mR��/͉�.���ܑ(V֭E���:���+���ޟsZsg���2�T��)�&�Z�����\��wLj*��!�����u��g�30�-�Zy�ִŠi�|�BKEG`��+ǅM�D�4�� �<���b=k�5c�C4�}�
�g�A--k��[q��iy���~�t>=��R��Ym���7B�T����L�9�X<��q7�q�y�ii��m;#���(C�.��|)\��U	�b!��\��-F�^��+_�����J	���߫Ȋ�*�5v�I���I�%S�{�����G��������',�5�����184��9���`}�Z�p��Z}�����>�<}�)]Pa��<Y
)@=���� �7�2����~��Z���a�pe)D��2G��k+����\z����%�Δ=�6���B1�>D�Ow��RI����L�']�����m��ݫO>���L�u��Jj�g����^�{�����[:�����HDs��j^3����}
5��ώ[��q�P�$G-�{W.@s{�ƹ �&��0ri�� "��\@����3yփ���&+�OK��6�y,�i�'�҄7F��R�Xp����B��}ރh��HxF~0��f[ߜj䨍�w߼������m[wh���R�ٽWg����l�`uu�V��\�RA*��N-�4ZH$$>E����(� 1����T9�ISbRJ���g+z녞�V��۱q�zmn>y�D�> 	μ�]�� �b)�d=|�#VU&�� �͚5���c�>����ʏ~����x�>���ܧSn��k�P&9��m�&)���ŋ����ߝ�H�F~r���fy��8�9�L%g�IGK�tGdެ�m�KS}J֬�ଓFM�9�H�Y��?�$�t�˰�`�Xh=��ݻw9-�5�?�A߆��0���z$�רR�qke���as�I"B�����Hr4>R��/�^l����znh qOC�=ި����A��?Y&kB���|�"k��J^/�,�`N3�+7����0!E�È��-�l���������uPj�M�3��>Hn\xnˤ�eeTq�`���J��(q�^-�tK�A�ZG��;V�0~M��5�{5����B����DP`)�~�����p��gr�	�U)��5ju�5��e-��Q)��@h��y&P� ������
;)��.���ƺL�n�
�.��*q�Y�^0_��Ovv���R�r�-�B�X(�������2�	�y��k�"�DBcȎ䕪?V%Y����ɺ5���W�Wtl��q��X��d���E(S���n�V�^-n��|eǿ�Ԕ��;��<��N3��&���@��x�:!,137�b`1;j�+# �{�sqn~�,�\�m\�^���&}d��,Nb�<�Y��}��,.~ǅc!�&�ce|9p}��p�b��Y��|{��W9��[I��O9���9W*�Q�(|�W�u}?������\�V�ٞ`��)_�g"��fˌ3PB�V���L�Rh���m�[O$�!t�Cyw2� �O\�����_t�j�7�nƟ��o|�6Up!¯�248�GAy�2Q�V	σ���MM-�(�%B1�8a�7��
<n,��њd��urÇ�In$'㜢��vI�!��6�&��W��d��c!H^vl^+�;_Z�1�p�Y({v��ޫ�07ٱk��w֩2i\�,{y��ޱ]A@~�}i��}$e �{��U �~�O/hօ�:e��2X+~�5�iJ�� ���w��#��GyD�����h,"&S+��gSs�$絒��u��8�ŸP,xi����)SU�q�g�E��T��2h<Lg>��jSƆ�D(��{����n��C&�������/n>?�s���-9L��ǿ��cV��{"�G�(U;*,� ��cI�W@�+���Եd��bL��N3W[Kc)m�+�=��_`�,��k�x:��V��������:��sT������|MFkKSxO�9d��<�7̍glS\��u� �\:��Ev)���(������ʸ�e��Y2��no�J$�Uiɪ�
�z��Tȫ�q`�fy�M�����m�d��M��(�t��k�(�����];�ɠsY�� �:N�#䃯u�������4C�DY�����P_��M>!���!����Ƒ�c��]�E��XE�����������.���ܲ5�1ƿ:��}S��d���]aҷ�|�ai]�b�P9�/�[��ͽ6H�e�J��ΊB��!`�.пwkh���$Ŵ���1�$)��6`I�3�s�ؖ� >��-�r��&&@��*F�ح�-	c7��F��9�k�����o�W�T(J����:IJ���p��;H�W��S
�A��@��2�N8[=փ�%��y�(���Yc�μΛ;YDM`J~��_�8@��P����_�����o)(�VJ2
�
+��2a�$U, ��g ��Pߢ�I�S�l�ay��e��;c�\r��;�L�#G��I74�D2Y̎�˓q�p�L���W��C����帓fI�\Z���69wg�l߼A��6Bu�$f���'���U�!1��ĉ�Ry<�#9�0A������Nlw�-��w4A�w��H|&׋�!�&�2�Vq�j���L���Fx;��3bac]ph�4����z�Ø`eY��@~h*��r��=��&Q�.�q�4������y�����)}Z�z�Xǁb|��ŅJ�������	�ì&�?Ðp$�AѸ�P�b:⿐��a�,�Z�Xsl�C�ް0�z@߰�PTVD�ra�7R�b�Xg���bhjm�h)�Y��o�-8ԕ5U�ҙ`,�?s�P^X?@3"N�dF�{�d�������,�7g6��Rcȹ3�qXJa8d��Tc�Nۄf��8;��ɒ!�u7�V�%���on��fL��{w9�e���6�(,y�L#�A��>+�ב�Q�C����l�&u�uc]#�{�S�@'6^#�Hf�$=߱6�6� =�4��K�"{�
7_������7�.�`�$�m�NXCh4Ĥ8����9l��-�Q(*���k��:���6~QU�;/�ڎ��5J�`��^-H�.���h�h�Y�P(ۏ݇�	��/_��6�#�rw*7|X .ɤT=��A`~�lm�4����D�����	sI!��w)ЌP�Wܓ)�� ϰ���կ�;�n6ո)�U[ؤ���Z�"RXzm	�z7@����sJ�q������>�9u�X�o�Z��^���� �s�v9���A WQ��en�RR�z���il�d��w����g�-�gr��3O���E.<�liki���.m��)�
�	��!_�H ������g�'���Z�c����� '��t�&��e#0h@��l7�8m.�.1��0-�g
��P���g��#B&K��1"������lH��-w����ɚ��a1GC��:c�3�8��!�F�������cNQS�|D<���0P~8�{s��(�Ώ��(s�0��vY���k�f����b0Rv�*�� l<�]�b+eAT�/�����R�P����ײN�Mv]�w�ۅ�U\cE\
������Ua�a�8���ϧ΂�y\U2��\�JsK�*]���`=��X�_��>ֳޙO�a����i�>6oب� ����	�R!�,�K)�V�t�=}�iq�[!�#�ki��XȆ�k��'Əs>���Ha�,�f��I��Db��d?e�$���&���n�P���I�����J;�����k$V�1 @��s]6&���c3���L��o�����}L���JF��U{�JF��ge�v_���$���'�<��C�K2
�z!��JH��;����o�5��0�f�V�'~ą�wi*�&+ɲJ�~:�T�룸!����!�D�E��Z�8��#�ԏ���%�����4��jD�+�N����K�U ���AX��e&N���,`���A��xg��S���B�]�oB��<��3f>����������U�Ni546I��c�]b���amڞL
CG��-�
�\
�ndh@/Y$m��˗��W7ʦ�[�E��طW&���LB�}�U��ˊ?�ަNW�~g�\x��Q ��4���bCW�0a����J��洶�ua�YϠ�?A50�nX
2;��`�|�Mh��׬r��i�xp2�I�G-�'��ݳV���@�2l�~a't�Z���H=��iҍ !�̢乌CÄtQ�-��t}�,g-W�nXEXi��ݡ�Xf�C���!��q+#��ĵ~u�����JWo���"���v�U�ݪ��k�����8B!ր-�H�(���3���`k����&����Z��S�|�ȝg��"`�Sa�:�>�Z;����%��Jk��b��(Nk��a����-*V�X�q�ed=�IMӏ�>S_z��Ƈ�B)��9�H�|vDNq�����7ˆ�d��9��iQ���Ƥt��FEM����n�fM�����~XE/:�8&��y��`-DiG]lU�Yl��{�t� ��~QTH����0�ܛ�0iy��$^�F��o�FU&@���8�q�QS�0+*䰸8��4��5>�]<�Nr�W+'0+��|\*��A)$�ֆ5Ê��Pɕ�uxD�p%؎�G���P�7Ŧ�,IQ-����jRQ�W��,��ĺ�1��g��9[iI�Y�z�N
������?Ќ@�\؀>��	0�v��B������@k���7����=ZT�N�zᅗ�ɧ��Ftn�3�۷m������,ʫ��"�]d��Ya�ܢZ(�Fge�e�z�?�@��0N�ςK�*�҃�m�����h���غy��ڱSN8~B�����1�i�q"��q�ܜ�3e��ӛ�B�t�jH��h�sNP�KA�S>?�Z��_T��ē�z�R�׌l����j#O�ņ#^B���x���}P%?�/z�0�6�:�$;x��5i��M-�Yy?c��I�s��=4�ĵ�7k�.�m���M�@X`,*�_p��P!���!��lhIb(<�UC��B$ ���T�f�1N�Nj�7����M,��bQ���a�٢�e���h7,~���j7��?=�Ұ*U���e�ZD�����j}��HƎ�{�q��t��毿�W���ʕ+�w�{Hv�y0�)@����t#�Vp�KȀCESqL�(��E�t���]��R�o��������Q4��1��L���]B�D����u��`�m(��6�|�E���}���k1�G�<����eK:0����h��}�223�yH���2�?���3NS3��f`K8�HUL}�2rN����6"�r�\e /n�W���N*��X���P-�b��"2(�gl32L&�q� �O;�b�'�xJ������<+ca��^Ʉ1a<���h�P�w��z�F=|����g�VF�V)�i�z1��I��e�"<I)�R2����D<�c�XO|j��:[�Ȋ��1\MA���k݀�)�(���� %V�=r�-�(q֢E���n�Y����K/�F�#��e��>3�V!`hf\w�w��d��{����{d�Rb��e�K��5��)��ױ6J�=>r�6-/2��if�͉��\�,����9}����g��ݳb�3ҝlN�w��l�<��n��@I���	8T��P=W�4��YuVE��t"Ĩd�v��v�Mmn��`BH��C1�:7�i�8��a�����*`��,�w�;�Ze�����07�|wc��4�O�3����Q]�:c��~!�Q)˽��f1y�@���x-nسQ���-Q��E��<�0�����`x����ุuRm�z��i�u{_Ӷ�Zgo���]�޷�e��Vf}%��ڌ7w�Q�o�SjXį���|��_WcP"1��=��3�|��8�r��>6,�����n�)фR;&9���>n�3��+ڜ�j��k�Bu�]���:>nw
	lJg�����c���I��dq�	��( X�y��\�|qD[�f�d����Q� K�o���~��`��RÓA����F�8�`Ѣ㤭��3d��U��m[8~a�bEⲠ���Z�-�g�S��@L�[�D)��&@�dZ�6���ӓc�_���V��㶙�{jq��O�$)�B��VK��[ސƗ��<{�l�����-����?����ػ4����G�MKej�8���ws_���Y�Ɋ0�p�%�t2�Y��1X��اw�8��������/ڥ2�Pn� &�%��	�� l�[���wl��6�G֖T�q��$�&�.�?��;�K�g�@)]�IkXV�|͊���H��cCs�̛7W�;����X!L �4��=�
�T���C�<&=}4대�.�f
����S�_�ŀ I$<*xѢc�o2�w������{�뮻4�o)dε�`�l٦Fɭ�#�6vGcC�8�&Cҭ�b�a���p&1�5+��Y��S��{�9?�W}tz�`³��]�a�."|IsK�z5m�Hm(6Ʀ6KMkځ���n��4w*Dg�,� ,�`DB�AR5>�^���X�;������	��|�-?�{���]3�N<3�~\��(������a�m�c��8i�U3�|��kY)��Uc�T��Cas1c��fK��o���&#�\�bP���j7����<je�����V	/���Щ:N�������Z�����c��' b5X{ƅ9b�q�q}���lwB��?�1-�=W���#l��qGPa�Ι;K�:z���m۶ȷ�������B)�>a�`�;%��=��e�8ܽ�K�l��w���cÃ�m�|�~5�������� �l��W�Tü&HJ��K��E�+|���<������AW�ȵ�}�����e�eÙ	i��\K[�o��(����ni�����4��7�E�&=��3�x�dc��u�A@����~<>��AZ�'�ɹ��Bf��ܷ`���P�(���9ʍȋ�P��lQ����o40��P��Z��[�<G�j�����~̾�*]���!ݰ�;���_V�N	
�Cl��z���#�An���2�5U��`b�i���xZ2Y�9ikkQ&7���r^(Y�K!�^ye�we��"˝�B\�]�}��>���I���=���x�%]ϰ�X���:^�M��L��k�c%`�7j�J�#i�C�॒w	xPk�����iU�P�NV��yD�$����+�u��	��"V|��Q��|��֦�~/�-i����9�0x��ڹ���(&��aYK����hE���
�-z��V�'���w��u�-1W!�m�K&X4d�h`e�z�{)-@�
������|�*X;Ƙ�e�T{�cWa�H�%�Sbt���W1�'�e����q<j��Za�v�뚅���"O?��<��c���BS��{"��es���5��;{�[�#&�bV8?�8�@�|�k_�g�}>�p� HD �/^\t������(n�2�t����;V���R��>�4�AiB��.�::�W�s�oO���"ͫ���	?���ù�Z���M*W_}�nZ��.�ndFL�1�31����w��3�k�r?����ea�5]�B���xKcFU�.�,
Kl���e��
�,:ƀ�Y1��gt������f� xȐq-ƙ�c�d�7��5I�O���kV?�&>F^��z�@��*��S|��r�k�O�����	;g� ����$!�B����T�#�R��\�t����y�&�(`.�/_�(Z(:֯_+>��S�����Q1)��w�s�\�nïIz.�Q�I_�F�����}�5�������4�Ƹ�QB�<�ƍϟs�ۏ\�8瞤��!�w�nY��w�}�EV���@��o+ �8�2��U��k��ֆ�G�����<�2L=�3Ѩ~0�*���ZX1�@�aC��]6�@� �>�ƵP6H���&���Ρ4����y�'�U�
�l�k���Ƴ��X/�ec�c�`e�3ּ��-�����
�B�X�^�co�P�泀[k��aӆ���g��|���D��H\�ǳ5�b��j|�Ǐ�u��'c�W�oL�W�\1�^��u���q����>����t��~X���á��&R�gU�cRvf�����[�+yx*�]�eꔩ��%"���j�2V�T�o�tv^��C��%H�
����Р̞1ÇK�cD����ϛ+uNZNtR��ZiRB�"ż�x�E�UaŠ3�A��{6�l,��f3����BgbZ���zH�]]y�]!�6i�Du��U�f�V������fW�* V��-n?,L��{&��(�amYͅ!�� a��Tp]Hb�S�|~$��4�gx8��c,��9�J�n����QY���/��/V�M�{�.I��BӠ]��J����@BK ���>��H9cc�U���]�Z�^���x���O��2S��4W�7��辽��#���s׮7�=�fڌ����0�.�+��,W�N+Ƌ"R� ��c]~n������;�S��o�UP���={��^�A�@��o(���$��$�v� &nRGm�������g ۷lՆ��f!h!Z�<|60Qm˰�٬��=\�jkSۀp~ �VY������?u�|�ZA�|(
交Uq� Ȕ0�&O�R��f�����9n�T���:�8�e��&ͺ�;Q�:���6*L�2Ɲ�%�6��p|߂׶A-�nV��y�����f��Ap{���+ߥѫ���,���]z�G=#�$�)�F��8�%+������K���w�̟߳���_-k��:�j�����'�}�w9f&���5��P����L��$B�z?�+�7EK��{��y�3mP��U�0��x�E�X���3�鬘tOOϑ���fs����RW_�'��c7�XsA&Ez�e���@���m|z�MJM|>gi^��q��`��4�K{Z��|}��������M�W��y�`���ײ�MJG���G���V��>�?�^���Fg1�߉���^�,7K��T�9��"�"�ڍ�`�X�Ǌ�L�Y�3BB�-��6k��'�b�)@h3?\��*d�2�r��T�Lr�AZ>ř�!��1�˰i��9�dhUqּ̺�)�. ������A���n��4&��s�ŰVSֈ�
ˠuI�E��Xנ�R!W��>vΆ�ZB�K��C�	�
P��J ��h��v�L���A����5t��.�fiA�:#���(��W�"��v[^��ܲ��~7�GN��V+��K}&��.%���I桀765��o�b.+�G�z� i��8�O;j��̰$FH�i3���#s��=o�t7B���E��9߁{uCaZL��.�*MXK����P)ˊ���¦��Z笎�X1���C�:6���ZJ��I�k���{f�X+��ڛƳ8q!�{hU2��q�X��(!X�p��i��������&Dű0X�^��5{�9�Uf9�7���걶�k���bc�q����hJ�T��H��n�Q#�`H]��2�v}�9U_ׯ�r]���<^����f.�����b�z}��rnk�P���5B�o��vMa3����戺<�|�(rA]*�Mґ���u)w3)_���(������p�]չ�>�:OON�ь4#Q	!	�%� ��dl��\6�G��{��������1`c!PBB	�,�&i4�'u�Jo��:ߩS��#q�戦��N�:g��^�[ߺ�>GdF��Tn���;���瞝<�Ȏ�*_e$p�G(�|*�Nr������>�N�Ќ�zQ���˭�H
%o	t�
��\�n��a�C�U��t�o�X�\����NK(i�"��̏V�8��!�)��+?[�VZh�RfY����y�2�|]�X" [d�)�($~�w޳�@�����m��ӛ�ė[=�G]��B'��酢0>w)Gn��<��ۼ�NV�s9%?|/���Fy�H�3�̋���%�u����]���X@��gu���3p-kɿ��HT̘8�C-��$�qn�Z���T@��C�ڂ[�7��g�����R�4V�̷��v�f�F���W}�3S�ʃ� ��g�c���a��mf�� ]b-�J=
�DY�A����z{2�G9kX�&W��$i���G̠y�F��م��DpM�l�ڻ��݋��g�4���~R(y7$f���k.�G��G��x�I����.�.L�Pi�*F"�
N�.�b*
���K����<�JT���Maf��m|����5L̸�PJ��E���b�Ї	(1/u6dL��"�V�r��vb�:Ǹs����w��aa��:eHo�0��)�q�݈63Ҷu�v�=�+�Y[�����4�b:�k���Z3��k��J٦�x��@1n����ӟ�t6��Ub�tr�tG��W�)I�XI;����PnVC�P|���y�F[��֬�:
Y�@��"�I���T�o05��R�Vu���ie�r�Ji
O��rNQ��
	��n��(�'�����f�J����>��l�pu&�u�n��u����-,Q�({�B
�	�|�U�\
����_�B&~"9��d��n5i|�'NƵQ,d���'���^�H������������
�/��~**��\me�i9��OKi�	����ds�������hZF���З2N�>��#�@=��g���{0�� ��7�)��%�Ҋy}gKR̒�"�g�R��?g{��U��uƞ�C�O���H�����@s�Z�R3i�@�_��Y#{mGڸms4�N�s���޾݅�3�C�+�~42MY,fAW�h+o��x�̗LwW��\��ޱ
��ǩ�Ŕ��_�`����ҘG7W��h6�3_/�m�ꦀ:���k�ȍ����l9U�-)f��D�y�@q'
_�Y��"S<@�(������{���3��^)ݗZQޏ�y��I�ǬZan���Ï�=;w��E�ųs�n�V��h
I���ws��s��m�I��(_ɸF��1��կ~eX�|���<��J֞�R[�Cޢ�&���=�y�J1�����Kܣ�Y͕r�	^������Xr��0(�?99Q�V��+�2�7P��F�}��#Beqe�ڙxv#0�"X� ?�fr_�E�T�u�����m�@z��8���հd��qx��b�m����^��̊��׹SufY��Ntd���p$鏝1kx��:�+�b�u�ƤsĤ�$Y%VY���A��`�aU�y�P��o�T*E�pp(�b�N�D�D(�Y���0�ٻ�\���^���׮3� AY� �q�Եb_���MwK�l�CR�d�w�Ŗ�D�Ѣ�і�j�1<\@��w��܌�r����8r~t�q�@�Q�(�ի�8�gl*]�rŊnq�JBFsk�����T���D�t!��O;JغX�Le��ʒ:��T�
�<f��W^y���,���=��9�Ł5#�M�U�(���&�Z.%aՊ�ស�F��3V.���b93��� 0�-�@���
�*(�Y���\1�fq� PJ�ǘ�"�&7�x��ً/
<p�-�w��kK��;�(8;j�'pҽ�w�ù*�B�]������p���NkA���^�����<7;<�������j�ؽD5)�C
�rc���c�G^GAC9�ø���/͠��W�YJ�@[f:Vd-� �=4~����7�b�� F������x~�^5ҹh$��E~�:�nV,����[�E�+�3)�ȭ��0r`����g���M7�����[��a*�?��8S!e������=��Vڥ��7>�m�q퍊�ZI1X�fMyFs$,_��y�C�h�e�@�*��?��<�qd���ɤP*5I9NdZ@���eǶ�aeܱ�_&�&m'i�hB~�I*T7ퟮ���V�E��Z)s��)�|x��4z/�5O�DB���n� x?�3,����`�8r�ƍ��ܾ�[����u_�M���v���I�P���M�3m&�����9��I�u����~��3�ƌ��� Y98�g~sO��Θ_��\�#��BO�	r��`aX�ͦ�� �r�_'FM8a�C9�٢E�L�㪫�a���x��g�]�Lsq.���0n���W�Z=��ӥ�{�x,���͊�,Y��@��~�`�5<8z S��"`U� q�)Oc�SZ��-cmloMey��B1s�Z3ZV�-a�мpKTxP'V�g,���/yi�햟Y�?���f'S�)N{B8%F���h�J�j[)	1�Z"��{<�ɰ˃�B���L�t�$�ɳ8�s�,U��t�)f��qj��y� �E��B��h֛N<�8���nd�ZA;�*F�c�h��5���+��u{p�e�FҪX�^x:W�_��8����L��a�E��!0�QѺ�\��X�tY�z*�a���J�t���kO�PF�C�Q>���������F@���S��?�xг�a�u�~->&K5��g�:�恃�2�Z�M�������IAc������-(��k�Z�K/�4��e/���l�֦ Hxg|C�;R��b.h���79a�7����]{d�ܑ����On����S?d��l}W�Ы��dȚi��z՘���㏷1%;�|�Rg�Ȋ6�6��Z�����v�Nـ�0��~����-��V�O AᆘG����#zS*�r��!O����G�B�T
�FӍ�����a��˭ee��̏o5g��V���������8!g�����c!�X���	E5,2�ĜˤsB��u̕޳q�er���?�V`��t֨h�P Z���c��fh��� bH��?~mرk��l~��o��o�bO�gQ ��k�q����`dd�!_9��c����W��z�`1�ׇ8�����o�52��q����f��,X곝���G�����������L)u�����ӟi�c��3S�g�m��b\6<�6�4
X�8���~@Gy��Gl�G�p��e��-n��O�|w�o��e��gà�w�]e�}+3ʡM��(��Gٻ(;	h����E��6wI����@��-�bR
��YeV���1Ѕ����������Z$��0
�N}�4��J9K�D�@0H����Qt��3�@�����7�9.�(ݬ�_53׵�OJ%D����!��g�J�u1ӳpp3�6ĺ`'E��lO��U��p�I1~�ݵ�i�<��X��-	q>�
� q,z��nB#�bC��%��g��Щ�t�~6+>�t�0I�R:?�RX�LN4G"�f\tO�dl.s3de�0���F^!J���ocɘ�]v�}�OC�&�X�Y�l2{�ʧ��0{�r�qj���&��pC���˶����-_�ǢA`�p�xd��)yv�T��`�"� 3Q�w�
E�}Q���nׄ�������g���r���l��,���5�@)U�_pB��e����<���f��Ĭ{:�IO�M���B3��D[�^��v>5�q�
B�Hj5�k,h�*�D��j�vא�\P�k֮C���l��pJ����-%i�e�)��㎷�! I楧�g ~�������qA}�_	_���M���L�L�J_o`32�3ͪԍ&QJ���3������H�J�B�a{��a�ۚk�vh������ǃWs�'�3��|V�)�F-�q���tp�ɖ�ߴ��<��1��Ir��B���f�t&G-7��$q�Wjx���bN^�iW�O��n6��"Y7mJ��;W��8�m4������XP�J�h���Ń�D۽c�c!f(*�6R���!~�9�F(�
m�<�Z�g!�^rT-�T����f��С�N���i�@s�}�S[ ���g���+������[c���$�/�L�
�y�i��e�@���g�c�0>���������-��_���D�6m��C�c���.x7�=�A(����,��Í)[=��V��SmB��o=?0���4��d�ȕ�g��E�.)�D��`z�9Uf�{[r��I�~��(N�{���u���i�����:[�ڞ#}��#��`��h��R�����Q P�bn��T ���Tפ�gt� 2칎#[mܨ��������iÞ��p`ϡ0<8d��`'L�>(倹\�J��Tʥ�B{@��)�/Q�Q�МI_�e&=�11>�)^O���E5s�Y��D��"X�w��ۢ����K��J�3���O�P��g��$>AmAa!c�ȭ��a�������s��/��^����k<���o�+��o6A���Mi�D��	U͐W��9�?�qU#�B��7_o���p�ڔe¡V�XX2��Qʩ�j��͏����F	��V�܌��*��t
iV�{*��4���*�>��y��+P�ȴڹ�P�$!�q��-������7@�A� ���������dn��&�ҹ/�36s��Ac�|=�qDJ�
)���at"�%a(�z%$���l������D^$0�L�th��|d�
�0a�Y(���-]�i�f��+H	���g �r�xڬ�Σ[����ʯ�6u*����/���X��@ ,`C�0y��s����5��a(��G�x����UW]�5B�b&K��ʼ�6^�j�e�H���y��j�2�I3[��AJW.�Y�)�hG3�Z�w�dd@�qn���GJOMM���R1,N;5hA'm���J�q�BK�Sұh���cAq.��E8�C�t�pO�����z��}S�dM)�4,���Vn�����T���|�)�d�5��{~i��8��(�m�T�;�qd]��S,W����������K��R�D�� �۩d~�:aJ-�V��u�H�yB! ����g�`$��yv=&�r�\]عk�܅]��c<��ҫ����НnPބ�k�=� �[-�3AIOKa�<I
U�T���-�Я�LQ�07�t��΍�0E���g��4X>jn�����Mo���m;L�׭;��ԱH�2`܃����W�Z��W�m�hF�F`�
��h�*%>��K� /B5�]�V�h'?����]�z"Y�(L6s��~�#�YT�H���#�}�u[� T��
����;�Cʭ���/�Q&������}(�s�9˲=*1����c鴀�SLc8��>YKR����ͬ�b+��YV-�w�ғ�sax�;ߙ��e��z��� �GT�4I!���;86D!�]t����0p�b2�wl�Q-�Lv!8�/.���M�>�-�V��њX���N�d��-�����?���H44���=\�����?ܹO�s�l��6�%�,_㖪eP�<��3tf\�`��.�B���g����bSB<����B�v�8vg[q1�O|�3��E�8]g�����@�
{�]��T�,0dB�,�{���%��D���I���:��2o:�\���������f<۲eK쳓i�T�Z4��J���_�&�X����Ăۺe�-|��OMe ��xٹI��Ek3���.��l�R2������%k��GJ���B3���Y���B)͋���6X�E�*�g�N:��vL�	�[�f����ژ�L��vx<�H�5�@P��9�������l���A`YD,DP�"o�B8�N긛"�ܺE�;�Vl%�g.��w��z3��i�81��� 
傂+���;�8���G7wu���ªU����N�gcq��gZ��믿>.�kma3�K�,KwA�ӷ���)��Н��B�ӊ��k�*F�E�D�E��;�?}���cya%�~�m�A�u���ĊĶo�LL��r�h�Z�-�f-Z��B�A���M�����	)�)��0�7��dLM����;�����i���H,	���B1��p/�n�w{6ΕK���5/��\�\��4@�Y.(��|��|�6�Y���{a�Ɋ��u���6�b#طo1���S(�a�'���w�J�j�,����w�e��3��L��/��S���<�X,���jX�-J���wL���\Gt	he�d!�������G^��0݃��C�-��v~�!dq%�r��*�� K<�W\a�v4Ɔ��9���F��	n���W{�Z���/|a�=f�p}�)X��"[�;�i�1ɣO���\��y�^Lp��I�!s䕺O��q.�)�&����)<�2\6��y���ȗ鋥.����s��<�(?�3��Q��Ž ���a�x�W���:r]��M��6�|̩3�럛M}��V�-AV��3�p���_�e����9:z�����h5����r�3���kG�sb,������~��&�`��L���p�H���2S�5`!��[���A�w˖�V�w�g�u��q�\��E���ۋ�,��5x+sZ�����s<]��͔T�ktS*����8�L���J�Q��/� �1:z���?��8N�2�����xج�l۶��XV�8&�EW�S��'�t��@t�J'6>T�b\I�Ej���s���\�6�T�Cm��\=���-��t����k�ad�.��`�A�����3d	�|�	+5@�,_�Ԭ�o��4�6=i�d\��3�%-��z�~`b3K�TIc:�3�7��,LI��̲��Go�V5Y�;��aqFl�3�ڻˬ@s��8��,U���Vq~3m��轎�bmXL	���i��m���%3��rM���=`[#JI��hV�P�U
Y�ұ�p|���&��2`�Ī��"J�V�p˯�5�S('唏±%�L�A�=�c)�N��|Zx�U�����5�&zgv�3 {8�b��r�����9�|A�v5��P �A�gǕ�;AcQ��k�k�r���X��<E{��ZI}�-�/|���������(�P��w�vE�seP�)��I�241��xE�2
,�������e�|a�0,R~�WH֏*i�⼩B�N�O����eY�}Ȥ��*ͭ�e�,)�PԚD0�&bT�R�C ���}�ӏ��٢�7��{
�lN��2����^JI�{��q@k��εa�%����]bP�gf�'����Y�Ppd��G��B�H=�۰��3vB�4p9��p���MG��!A�Pg�ﱲlv)�����s���-�f����二��J)�D���I���8:��::c+��J7˥mgy�9:�!�Bf��+��������jK����rgtA9�]��S�E��v�W��#{�e�����`р�Z)v���Ê}M��}z&˔��pV�F����	�lK��;�ݚ}�i<��&�w�M� �%�%�2>|
TI �m,���L���jC�%̺Y&w�{��]�(�>mMsIP7S����ۀ�w
Yʘ��s��$E��'|��_���J���k�AuzI�I�T��R7��j�бnq3t��B�R���u�pnܨ�gSOJ�r󨦍��fR�76c	��P!,Y4l�:59m���Pv���h6��U����<�WƼ/�׽��	�R�(b$L�����l�7\������w�������f��*�\檮��^O�,��\��u��g�����xF��S�|� �q�3��$���L��]��Ү^�KV�U�j��R!�P�xx�x�N�S�k��u)�BА��
��}�_���,�-[<��(?���5J�j
�x��k�2G�8�����=&+մ>�Fc���%�=g<�0�?GH-�b�'K���e�B���8c.mD���l�=�@�����e���|�����N�Ro�)4j�ʖ���a	��u	��]O[&M
p�ڵ��(R�9�7�G���ޗ
��T=�0V-�=�!,�֠�/[��\-���ҍ�4e�'�n:��"��r������<4� qk�,MX��C�{͔�Bc�$��ԅ%����v��~� ~���a����Y
�Y�]�% �����(�3waX����;9L�0�N�  ;�q�"پc��E�=}�`!R�Z4��)�~L�L�(�����Z�_k�5�ps,
����t\-�+���peX��|�g<&Ma-X�ȞK�K�HV�@�lLk�=.ŷ�؜	b�y�K��B��{�( O&&S��"�|�2By<�e���'�t�qo��Dؽg���{��^l۴gt��`��zY.�UL{�`��l�do�T�=��𲗽"�;�Dv���2�A�Y$~��#��J�eÊ�>�)��.���;��B��|�dN��u�{����2Wpj2�sԈ���S(`l��f��3��������I�G�1V�Ze�.�[�l#��5�V�D�5�23�6��A���(	^R����*�v�,�P�:::a���i��P����NE������{���-�G�Τ�Q�X��BIP5z� Hұe,biwv��k�����j�M��P3�=��;>h�3Ӫ�Qի�T��}ÆG�E0?\p����'�E�C����W�M
�ߟ2����]Z�Tۥx����U���k16Ĕ��u������cmVg�����2D_�
�o�M�\̸�{z�k�8�u *#�Dd���?r��	ף���Ŵ���gm�b59^�'c�7`�T�v&�*g� C����.X��(�o���ݺ���?��2Ҟ}����B��h�$L�#�6�ɬ!0h�G{<ԣB�Ώ~<>���Tư�C� 0�)��/��3n�vk�`�4?^�YZ��RH��k��-.�G2��!�k����r�3�ƍ[3�T�Y\������?�<���ՙ+P���\>��J=
u�8QW�{))%��W(�"Q����(��d;��%�~b���ۛucĢ�P�-o� *�7�6X��_o�N`U�v4Ξέgip���&T�C��B�
uˡ��y�\�*�}>Oڛ��7�d�
�/<�-)�U�wh̉���t[�b�c�~]\j-�-۞��VF�iɲ�Qq�Vϓ���f����l|Q<R�FyYK-�1K����!&yec٧4Ʀ��|M��b9�bWn��¤�D���6�jV��B�P�~�T�<d1j�$����@lAx����R'�|����� L��|�Ҽ{��T��Ph��\܅�;���:��\(���O����?�d,����g������l��p�H�86ۡ֝�w*���ཱྀ��$���l��y���0Si�3�U�+���~;�zF�e��f+քR�K��ٝAcu�kĝ\�'�ݦ�Gj�x��d3Kej�Ѹ�p-�v[e�<�SJY�&mq���ȸ/	�����g��g�91�Ȕ��k��_#E�j#EhÛl5h�]���p�`�7���=��5��и������.�˥l��S��Qm��u�Dޭ��P�0=#U�R�_���$!�,1bTڔ�{jD�R;�
%�[(�(�b�?L�=�UH��A���1 hߡ�P�7Je�1-�T���­�l�l�fV2��n}°)|)H1�5�1�o��id���@�t���>������oW��4�B��w�U���/�2T��T��w�8J;�ҝy�y��˙b�d�לĩ��b�4�Z���������K>�g���<rߝ���)=Y��Ϝ�p���ڵ��*���^��  ��IDAT;mJһV-��UK��SN����/~���d.��@o{���[��Iu&�/����̴��S6A��qb�7l�7+��,U���=C���v^�և�oLUM�i�+��[�\ ���ΏQ7�u��pB�U[+m�C����!;��];���5G*�4OAtd�m�zR.��D΋q�ٽ�`�s��(���ph�@X�l�W\��f�z*��Ỳ�,GRmR곪�w��BT��B�I[��Q;f��6�)M�fF�Ʌ@h;�O�"�+)]�3�s8W�p�NKH,e�BjLU��;xo_�;7�R����
�z������bka+������������K����Ѝ&ܙW��fE�qQ=�/���-Q7: .@ѿGG�-0ݫ|}�L�[��=r��2!�%�ŉ����J�@�le�4W��d�/^�S�*�e�{����ġ�����\�B ;'�<ncQ�*�9��m�FE�k���h�S�,2#e˄�-u@�5�-���i��]��%#��?/O��m��5��k�ڿ�ͫ��{Y2��Q��4f���`5�'=��G��B�8GŶ��O8�8S�̃a5����_6��̃>��烯�Rx&�	c� j͵p߲e�Mȸ���:-ck�2��ivv��n
%t	���C�K�yM�}��?6��A��r?,�2�nU�J�)�ØB����%{�{�o�w�v=�XX%�iZ�-r-v=�~��!��>&�:���>hN�G���.���+�!��p����^aaB�����됒U(��ܫ�K=��m*G��@QG�|ot4�dJ����)�)~O�
�c�L�����-ZSq�mDk�20�O��
�m����D�e�?�d<�(�N�ɓhl��68)_͗U��?h�N���i�0'�ҏ#k���8�uӔ��ٰi[x�����K�3�<��9�;h��3)6"1�cB�EB<%Oa���@�:A �\�5�D<2�U�b� ��Z�Ϩ�(���f&�y�e�_���ܧ\�5�G7+�[P��Uw@�z*ZC�$�ȀRa��컖_S�W5=�,��`��ړ�>�
�5׹��K̲d�Ն67�	E򶷽�,B��l�A�>��t�(#a�^��u���P�(��7Xp��A kG�3�e�������5˼�p��t<m�U,d���[�=a�Jwq��>���2%YodhZY~@�zG�����ͧ���8^h�� �z������oɧJ���̣�W}?}��C����g�z���f+R�{G�P�.Ƣ��?t}8���9Gl��@����i7��VK3���� T8�%yp_�(ũO/A�l�ξ}#�a�~*�@��P^w�u��p�(�p���O5�6���ĔQs����?]śX��@���t?������@���2m�c��f�����5ǵ@ܾ�u��{�^���?���L�UW}˪���Ƽ��~�,�z5�����.��m�!��U!���R^A���{�	_��Wͅ�e*�6�9�^�o�Ay��t�u_{��Jԋ����2Yǁ�������St�� ��r��Z�;���a2r�WM��ʥּ�k�kxD�0{�m��H��(6�oG�����1o�]v����p�Mنm��}{�)��ѫ�)O����*���E�Î=#!ZaώC�m
&��@U��Dŕ��ԧN�7Zt�iT!)aR���J�\*�<�	�b��M�@����>碽˻��:]�N%�Y�ǺΕ�9\ܥ3^��Z���v>KY!�+OZ��B�~���ރ���yP 0�[�l��Z\2��7�)J@\���8�#aqW\_��8C��Y��U>ǹ�wg�%dJ���*"�V*��;���b��Za�p(����;x���ȼ�7�x��1�� x��#���y�y��n�EҚpY�ār��K.�,��Yr%��l����������[�#��EU-}�L�R�RT����u�,O���5+����7/�n{�T#��1I�/c-���[�PZ���NR��Hah��)e����n���4S��0 B�@�u�!�B��bnV�Zm�����@��%���o��9�:����"if��w�x�\��K�[G���|9�Z
\2vZ�O_(��d���3�,h�+cC�XQ"8Vcaۮ�0�'n&X�|��qFy�Ԗ�ü�ȱ$�1��o!��ӻ��.�& 'B�)��gy�{��n���	/��yV��bR''�� 1ߍ�ِ�VӳЭ�x6�;�:�=qV�QX���Ք��q����[�9lN#�s�(�J��9��:�s�����M�+iΖ����F)��ӦT����p�}{[����V��C����-�F���<��J���zbn����>1NY1?l�ذ �����%�r�MV*�� q�AbK���t8�o���Z���w��+%&�	U�&M+A�6n�p>�&��w������#��-3�y~^9<�u��v+`��"���G�FfL�B������b2�m�M�\K�\~�pp.)ze3��0�!����2�*�T� �$��8�b ��y�I�	��12����;Q����;hx��)!ރ��Sȣ�
��澸O�󱍏[��@T`���=%�e��R�)��)�nj6W�c�s��\��њ��S4�y�n�"��#_���]ˮ����5<'Ϭ�c�s��}޼y���ǣQp���RR�{�w1Z"��`���xS8�/�:l>n�R.v`h`�	��5��i��;���������FK�p�L�Z�,�/���X,yd��pM:}l� ��\fq<���p�:�z��HZ;���Q�2�d�m7��3��i�tSt״��#@�b\[@1�9,Nu�e#h��K�hl���Y�jr���<߼y�YX7~�>7������B3�Ey���g����{$
@�����.}�:ewEap?|2G���o����1�h_!x��j�kG-�4<����@1'�������t���>�,t�F)�V�LH��ecg�k^�:7S"�Q�Y�b�cɻ���Ye�8_��gW�Nh-��(m_�)5�=X*�0ǑmE
��(ZW�E�!̛�(|�?������m�n^v-��!�_i�F�W)ƌ�����
l������G��ȭ��;DÇ�����5��U��p�j�d<��S�h��8��ov���������_�L򂧝=_�$E(!�b�� -�>kO����T6�[h�gs��˔��<�ղl�*��?���O�jj=;e�{B�j���z��Ǜ���c�h��٘k�����P �ҳX�v�cd��l��856�G��	�h
m��}���fLfQ��H�"/���+�̗>RŐyʍVw �I
�u�3�w�7�|FH��|�w����8*󆵧:6�L��7�,��u�Ǣ�:�pq`����Y��;�ɟ7?lz`W`#D �سL�2�����΅�ɮ����F��A��ת�����nd���SLe,$4����d���������P9���TAѼ�k���.lI�g��:���N+����|�)�0��jJ�M��j؁��,󓇭��q0~^�_�L},��W��҈J)�������}/�^j_���9��#(�}��LA1�ʪU�����ʯ��%&;X+����-�����%� ��I�Gӷ�P��Iӫ0��"�*mi������k�6���RI�B�c��6�Z��bWD�����I!i��JE)+�X�f-��doY�|��'�����%���7ǧ���I�(�B%j�bO��zKF��M�Ukֆ��h��h�%_����B���(�;��OŬ�I��&��@Y0�_���[^�|����lw�*�{1w1������ܳ�ߝ������c�Ob�&���rݔI���
ȵ
���- �8�lp��.=��TȌ��Q$�����)�qws&��y��X�<􋧜r�Q0���d[|N���Q$��?itP,@���Cq��q�SMLZ�S�&6'�^����z�%�8~��~/�؊M������֘�������)����>w��b)���;��NS���'���� 5�J10WKGCe11U�26��S��@�3�"�Gs��&.椔]�T([1�^~_�]6s��	-@4Ev���{�R��d���o�O�]�vƖ�����}��f�>0�Q5T�Űc��p�Ono����a��=a`x~���3��`ⲇ���}�{lc�n~5Ke��޾4�T��=}qB'gYN#8�
�����\q�����|�[êc�۞�j�F��m���T�z�t��]�Z�ZJ���e�#k6�IR�V��
RH��{����iG��9�X���Bq��N�]=X]o#�&�䱣z8��v�q�s��}��B��k-���ᤓ�a`�JeA�=
�g+�N,C1�B�����x=X���32��
� �	��Q����p��ebf�f}��mP�Q,xLwK�k�u�=���z����� ն�r*�B.r�dc_ws"��3 )	�jT2\�(�%C�6�U2z(N�I `w+��j��eujz"K�:a<�Yz ������*�+g�|K��=���[v�bb��r^b240h<'����Jq�=�b2�{��h\�7����M^<���[�x�ƕ�8�{w�q�df*L��W�&���)%�siN٦���G )=����e+ç��s�/~Aزus��K/7��o3m�oTy<8)CvvJ�)'D3���Вb��{�����߲ �����C��c�r�IQ(�	K���{���`��ˣJ\���U�Y�:U0�Jj�q��IJ��l�k�P����W�,�L�2�g,/���ܹ;��X��gܠy`�WS0�cNK�����,&��%��N�V�7l�Y����+w��[������w~�q���Q�i5y�������=��r*H���������뮳�B]t����~�3���{.K2;
�'w�}I32*�H���[�v�;��+��2q�l�����S/��6n�����"Wܳ��1[�������Q:���	�vL!�X��
���G.��j�ʁ�}��N-��I3<;���ct��,�i���BTfG���	J#��S3�e�m|o88:.��;w'
0�5�����wZi\��sP(\w���B)�;�H���RH:��sm�����:�z�����F QT��� c&zb�T��3"�)ټk���֣w����y?G��+�z�UB�/T��!d`.&��Ց�X(��4.1;���>da����g�~�} XN�\�$�j�X���\��
x�/��C��1>p`�}�3�iܿ�6=n�a���A���?ϲ}Ƕ�ɜ~���\6c��M�8

��5eɜ�\��7��\J�O]Y��a��Ũ��,�
JER�Hn/+��
c<�E�2����yĢڰis8x��Y�B���@9����2:I�s�d��ֆhK��h���X�w�u�]� �+�6:�(b�_V����tjE�8�
�$d9�b�z�`5�[�(<��k�c�og�y�	��_��p��?�4'�G|h�]�Xk���(���<��Y���z�-���e���)����p�Vk��M�63�ՒT�����k!�&2t*����{�����!63	Jp��[��W8��Z�b�!����Şt����xP�`�8��;�nc&S0�߭^�,h�@P�,pP�(q��U��qDi���/7�F��EqN�����O�Kpxn���b��{��y~ �ǭ]g��s�q�	-[H�s��=�m����h��Ȕ�H�*��t,N�䉠(ϱ~��&o�3X�(kPvֹv�D	�rh��;�)�%9�k�-��b�2�QG�bt#�V}Q��3��G���?������/����hUh���KsX� sg4��c��z���5ǅ����W��������C�ԓO
����]��{-l	C�l\��R�A8{˥�]j�㩃<��kQ���n��<�V1��DE�8�H�4+��+�N�#�;7�����f�Q(fY*��ˣ{T��|��ˎ�gh�.�����B�U�'��Y��p������gѢ�,��ȿ��O�3�w/}�KM�pΧ>���},Këm�7�t(������{�1����\���=�l��y�$�!M�K�7������YR��k���S;���8��,v)~E�ڕO#�[��k��{+YF��h��}i;��l�q�o�駡�r�"ǢH�98�98-���se<�k �l�33X�@�i�ce#�.Z���nPfIժF��p~mC�2�����/��B����EQC��'w��}�F����yQ�2E���%����,�����?ݸ%�F�w�I'��7n�̢0�}��b#��{*��ف�,Y����0mKC�j>�B�	W!�E�S}Y�TZń@�s��T<P6[ ��f�1�Ri�N��E:_�b�����U���5r���l�s`��С
����f|��UBa�����]��o����A#0\\�H hX�BS���JL�ae�p�8#���͎M{S��Y,|�%�g(v|*|7ʎxɏ��>KYs��������h���kԖ?�ž��y�ow�k)Ѻ� a�q�(=�ӎz�@���a�xǪD���<p/MAƍ����P�!�R�ˢ{T����:T���Q�ȚSF��k3��K?��q�޵;n&�L�VI��k�@3)%Q�+G)�b,��B!
NP�>�#�²�yaj2��d8����]��N9ى����096n���Ã�K��0S��$�h˖/	�}� &�$s�!�¾f��`!YJp�ó'&��XA*Y:Lw��MGfe�5���Ͷݭ�eҙ�Q�$/�y�>u�g���4(υ@�o��ݻwf��ha��rb���IȺ`1`��t
���E>弿���UU0�!������;TP&t2{;���c7$�k�C�b��}�/,5�������?��#�~y����s]b#|�� bNk���O����Ou$i�8M�]�_���������L.�{4*�R�([\Q�%oI�FY����3g��Lc���\�b�e�H( Ǫo�'o5*��[���X�1Y���М��7$���Y�˲�TGܓ�Ro�:���L���}��<�.OR0;,{�	\��ǅ�i�#�w������}2�{���6Ή(�{�f'm���C�4��]v�	��;��}:_�ͤ-���fl��u�o�Ik\MP$�T��?Wo��wuq�z�B{M�v�7Rvy�g�w�i���g��=v-�bU�J���UǤx�v,'�q�=��z
��(�=�y�=3;(cB|�����\��1V��\#+�SP]�σ��?���w��.�aU�����Dm8���~�_��[��PU5�b�=����=ͷӠv����N|O�w#��~��鸎�_,(hq��Ma�V�P*g�=B�2�(�9�es�Ŋ����ͤA[r�ztϧ�۰
f��dw�{d��3��1�ͩ��vY�u�`��Vl���a*����tRC��^���@,��t�%#QL�S�~v�=V�<9�|͚�F<��?� ��	����?6��w�����#�r�`NP�(�j�Vd��-bQ�> �7��M��7���Tj��1�)U���Z��9��[�	�W*�ߘÜK� E �����o��=��P�
�xVvi���&u��4*��U��U�{3�A��4g�����=0������J���|��*�,�8n��g2����G}̄�F�d���
�crb�֚5������Nx��4÷����{��R�+1 �Y��f�s�%RGì�8)�w���@{=q,�ˌ��y�$S@�"��Q��aMA�(P���o����Ǹ�50�,N3�j�W��z[\�w��5�yM�7<h�[��W}��>�o�	��g�<��S�2���<A����cV���J���9�6���m~�Ԛ�s�m�ЭO�j{�j���0�#�P�Ӎ%��R1Tz�,�<��^�k�p�ɧ���`�zMF�ac`����TJY�6�q�{I2��G'ɯ�)��a"M����Z�by
�*d;�7���F�J���uYXV}�*)1.�p1|�װ� �aU�̀`�J�YXj�!�G��
afJ)wh�wՊ)S��,��ȵ����W_�q�If���M�x�m��� e�q]��>�jU%�(��u�N>�����M����g��E���2���d�q��m�dVe�{��%�vƀa12ޔ� ��b�1>d�\����C�峸G�&<�������m�PL|'��(��RƆ�S��[eX3���b+�A��5d��LH��~��w���8W��m��Y�NxF�/���c�k�ڐi>�qDJ�c�����L�w~O�N
�S��|���'�ݹà۠^�xf��a���~�'��9���M��M���g�[��P�:_l�8th���{���+
��'�d�%�@�Y1��k�A����BI߯
M�[M�Q���7&�w=L�kL�x�Q�t�=3񋣙���R���V3r��x�f
��*Vbd�M��L4�1>}���.���}}�k��ZN=F�l�8�	�?��Y���<7��5<�3c zl��z�d�xue�o�%K�Y�`��-f]�C�w�s�u��$\y���N	���H���ڙsɱ�ZL���,��SA37'���Z���Bi�|�*�a���p׬]m�X�\>!���\�|���\��8���Y���rc��n�ݠ3O?=�ܾ=�î���&��X�-b��x{�b�&�Ħ�D'E�];G2��v@%]�����a������6���@	MsA_�X��� ۨ? ԛ4Zܝ#c�/*ԕ����7�����s/|~���-�� UF�[4���ō�җ�����R�Ţw�3s8�?7O7 �EV�2ڕy���GN]��� ��r},��C�Y��<�Y����W�2��{'�B"�I�]��[���q��]��c��9
Y,�>b�	BL��C�?xv}au8�*3�Լ@/I�����;�SlW��]k�v�^	�%4'c��0ߋ�,����� i"���V�������r��rX}���[�)���V>�����I�%I��$�Qg�F�5sڥ-΢���<Yf���
;����Q:koT)m.[�[�LL��u8I�%Zi끌��J`�����T>! ��ރ�f����lun��)ݸqSt5O
��O������RO³�����
�ڴ�� i�M��D�h�$Ԭ 
�x��9�����;�
/8�p�ׅ��a���>)��&-b�F?���E�!L�]�KOŃ�
�}b�^/2��L��@�"�8D{�)�b��⻶n�fd<B��:r���ro9�ǘʚD���N�@�!�щՁAI�@��c�'@���y\�8�C�T�q�J1<Ⱦ�41�24d�_��V�,-oC1i�n�a�ƅ0b���\�s�y�R[�|�<�
\��@��z��ܼ��o�y�ˣb�>��?�:!������Z�^��a%s�,�F�^�QH�i ;W��$��xP�^����ƹ����tt����f��|�I|qO�O�g�[�Zر��p�Oo1�eǎ'm�ڷv ��u���d���^'���Jw��!�$�C־7u=]��m��A'�vY��P��H|�xv�[n�`��������ۚ�R�7�F�}z
/������qE�1-��J�Uc�t\�(����_qi��}4��5߱]h�$��x>
Cq�;1<J��lvV�:�띘�tB�2�������.�������8�x�i����T����C Y�C8�X\��/�� �B����������ى;�[��H��p_`�a�?��ӌf)�CvF�#bf����U���^�(*�kMp������r@)��؇�Oo�݈�(�{��_�_d(�/}��f�a�t��B@��8����i#��xm&ۉ�2�ʹ���v������G��['� ��UbU����E���f��Q<�jjBZ)\of�+j�,�׃�������أ��|<�e�ā��a��b���3���4��4��dR�T�nY�㎏��!K���&��Ӆ���Pf|h�?�f��������V������0:֌?��U3Fr�R���H[#�jv�'�Y�k�?��*"啥 g}i� ΁`��_��W,����8�
ʍ5�����:�R�Y�$�9�3u����c5X�
�aaq?,j��e����LD������^��`�*�'�����$�����r�Z�kZi[r��>8�Q��߅��g�e�ރ��Y�,�m���8�����7�pCX�~���Qj�����c'��-�~�ϓ�cN�v�nK����d�V!�L��2��i��;�щ�yڲ��J�p�b�u8^��0�Ɛx���?�z���2���L�/1�YL���G��=�����[��$ؠd3���]O��m|2o�L���3�M�(�!?.�s���&F��	wP|���(�\�P��.�.%5��n��BaVt���B�wR!# P*�CC�����z�������]��֬U'Cm�V��|T�'*�1�_�W�ų��e�;>�z��`UvC��gpò�������ɰgd�Y��G*�]S>k���}a �&γ��~�<���|/�O�V
Q�"��V��,^5��,3\;*jż��"�r z��3Pý�M�m<��ĔJ�Ag�a��<PZX5�(p�耧1����\K����'�'Tc��Ʒ3�5,�%�W���R�W��(��K���i���3�޳���������G���-"/�ߜ��k���Qr�9�	NyZWv�Ȣ�*Ψ<Ӷ����F���L����	.䘙�a����� ���;w�k==5m���=m֏R��4�Y����ǀ��J��̭[6�%�< O�`�"�gja咥a��at:��@��E�5�.<�qd
j#e	5�?����T�g�l|&�䋏7������z��5�����;�vl�;�f��D��V�w�x����Y���gG����١����j���ѽX>��DW�q[�,ʵk�5Y�����-(41滑y��a&N8�c^�t�q�K268bf>�8A�ϟg��u,��'Y�b*c���*��N��y���,{�q���(��Qb3�����8`h��g�ein>'F�����)���F��`V,[���E��{~a��\�O%��c�i)=��b8�����O�g�~�e��?/�;���Q$jfD�=�Yڹ��&:F�
&��/po����F5,\�������ʕ���EjA��٢-̆��d6X@,N*2��hY-�ҧDWie|f�t�hZّ�27�!Z�J���F���xʉ��hu���aŪa��-f5��QGT��l!�vZ��D/i,��A��kD��F+�,�Jo�d��J��"s��BhuG��sQl�5V�9��?�[������#�Px�{�c����<��yA������G���(��2�[*4���*��j��XV-��+�����S�D�����xسw_���GC��p841'ะg���}��������ǯ� �K^r�	�Ȅ{����B�&�˱}�3���p(~��T���d@���/}�X51�Y ml�����ܗ�B�29X�`���}Sf��jR� J��#�(.��2��r�bH��U��@3����CjFwSV��U��tT����L�(�}�9�!��R��LJ���)R/����
=z��_`X�{f�)"�,>� 6�!���- �Xd���R��tu*���	:����oxC8f�j�Q{d�)��z$M׳�f��=ֶ��ޙ��t��av���iq�b�����ϵ^irj4���)DR�7o
�>��������Y���ԉ��)� )x����}QyWk�6�jo�����J�8�P�Y���3�nݕ-��kll(�n���'���������� w򩾁����þ������x�ެ���p8zY�z��,ڍ�/8�#=�ڨG��T��?	�vX�"�!K��捏�{wG%2i�,��f1a���E����ހ5����ɪ�R��deAb�=�Ė��/|9��� �%���<)�LO���i�+�s=��}�F�.U���-V7���>*�k�b�֔W������)J��@�?#
�/S��5;�aRR8�s�ֲ�/��	h}��zͫ���3��/2��:�'��mD�NVs�B�CҔ�8f��kW��e#�e-Zv}�����ݙv-LR���q;�>X���?;��h�|#�>�o�=s���Bx��h�����\&CS&^��nSh��jd��L��Og�ݾ'�˛��.��Jd���n���J߰ɺ6�y�=����� ��O�iq���,�\)�8��\V��B6@���{it�C���x�[^�_��y�\�3�>KLL��2�;و�C��X-V\L�LvK�/���'I����]�m�U(Ī�	�l�{��W܌��c�D���LN9��p�0��00oQtg�;�(��w{|CXA��&*���!G���������^�{��N����V��!�	S�+.~����� ";��m[���G�QLtY&Ti6���I�XTb��PX���}B���س�7�;��E9�T�)��>���Ju#"m��\�?��?2�F��m��{��|G �0�� �M\��xJ�/�(�l�24�8���Pm/L���b%�e��gh�v�޶c� �������׾6���v߲���U=�8�@&5�k��x+�<�{Z̧���5����mn͕HY��Ն����!�{z9A�p��gY���{��RAg��%͌s'O���+sG�� �&8�ۍ���+u��g�qώ���419������zd���ַ��~��<��c�Ĭf4m��`����覕!��X�Y��˙fG�B�N`
��VY$>��|������Ѽ����{ ����	?������>lx��0�_\4�8`�<hn���}�_��𲗽�ӯǮ6T���O�"��4�t؂R��֔̈́]�h~�����"mv�k���eehV�$["�(�g���D�P�"qb2:w�c,���166j\�n&WR��q�P��d��ŴwN�*b>��w�Ӳ)���JCnX�/�mx$������2Ú�.��=~�Z�Ek(2,%���B�|Ď�o����7�r���w�����x"�n�Q�����t�X%�aZ��}�� q̶�J�V���ub���E�}������s�]iU�sy�&�ⶑ� ���6�T�I���J�����i�g;�S���^�[��6V9��T5|�3�>�я���?���}�Ct�6��@Ū�L�H�9Ł%��d�|бC�r�w��m���fӔ��}��!p��} 8LR���U���|O �b��,:��Ǭ4�Ǿ�	�x���T�Q�];��-��	W#*��V�I\����RO�+�]��<6��d5
g5>`�V/C���̄��;���SO����E�����3�22B^z��A�������00������k�e
:���L|�a;��PƋ[�~��$%+nsH{݈�p��w�A�T;��\���I�}j,"���P�2;.X��(P, �%�\w�-�|����LkŴB���%Z��UaE<X��4>�A�����S%����c�a�P��x�z�9q��F%z��x�p�L�*��Љ���כ�{ktXJ�����+Ԋ�9�#��9\@��)fG�C��(�+��"�x�I��cn��0�X ��AQ�I��K^z�)1�A �W�Ǣ*ifǻ���CUr/CC3�w��*M������i�Aǡ�8���BY6?�È���������M���(s�f�	�0���4���C_Ԯ�����n���NϹ��_wߦdK���q"/]d���g�����ؠa��$�V�=K�n������4*H��	O�7w'�ߺ�6I�Z��f�Q�(S!�xV�YT]<}O���'6��@��R��n��|V*03��t����Q2���9�� h{����DH9���Tq~���c��5�gn��g���/S<*j$�811Ն.V���I2�E�p)�rʰ�1e#*x�o��VN0o($�H'��$3������9sA���K �EW�-����A������.#�F\�4����Щ\
͆�_�3+�]�l�>� r�9��;6�-Yn����۳k�m**���`S��\c��=��\�qB��Y�z����l���$�4��A�i7S��j��y��w�PJ�T32D,L�M[,��5il�H�8g8ZчF'�.�qk�Z��תgJK�C�Q��Š�I鱷�HR�1mh~tGƀ�Y>}b���]�����AX�bq���f|�P��c6������&d횵�8�W��Т��i)Cy
�#��Z���?`Z���ΙgG7��b2�Y�`\�����"%��=tp,���k�E1el!�܍�=Y]�r����,\�U�*=+��S���}� ���ŉ�C�9��`�I�	��+޼���'��-��<B9c!���{ի^e
��,l./	u���
�B�L D��H��H�k���O_t�gR�)�A�ł|:G���ȸR�t
�YS-�EO�:�e� )�b12&(R�
�������ghp,���_n����E��qMڠ(�P��<d��ݛ�E [x�+^a�����c���]b�����UT�S3ap��PK�a��єm�h1O5o��,����0��P3��`�7?�de[H}ڦ�|�.�{_ɸH(Hھ{o μ?����V&ÓZ�#������6n�^��p���f�pu
���#/��;����X�^�7[r���?����M�)�v��;��kB���o^�.�Z�zY����t�Գ{��.%��p�q�᪈&NX�Z�h!�>\8B���X�s���`��j�{а&vI�m�S4���y0+���W7%�$�[�P�w�����/|����O���r�w��+W��h5�[���O�Sx��|gx�s/����@����W{܇jj+:��0���RT����i_���JfͤG3�+q���w�����G
]x���j�6IuN��x�?�AA���Ӿ��G���\9�*�Giឲࡒ@�P�m��i��s!�9��mo�>�gb�j� ݿ;�+�� C� !�##�\ޣ%�ڃ�zű+��X����B�����u>�;�C�&�����d�"26�R�N�d*}�z���58Q�D�?��`�a�o�`�ՙ�q5��#���/yiX�|����1�]D�n}B;�ƚ����^��-�E�wx^#@��8�[A}Y5�LX�W��L�F���Pn��0X,$��t���Ղ�w�"iG��$�%~����]�|��[�5������!.ʌy"�P���C���gҒ��l�p�6?n�������}^|1�$����mR̅�d�Hj�u�*��k�؅ЪX�&8���?�ub8d��F���
���UvL�<e�S\�����#��f\6O���RZ�#2�R��{�wd�V$۞x��Tj����̶bi��0�oO���G%3M�����+l͆�j��@Bg�m������M��i� �)���p�C�3�q\8f��}�cQ�8?�a/ 4���s�}v��~���.���y���������u�/4E�6��]�7��4�,������X$�C�B��W�1��MQ)��t����Ä�#��L$� �ؘ��� �v^��	�"X�uX\��-��x�jz+����v���f��1c�!XM�U
�Vh)�Y�����|�JGL"��Ҡ�A؋>����Y��|���׿��x��e�7��A1`-Ⓗ�W���%��q!N�eA�����7���?��1l��[��ś"�kd0u�ݔ�o+��/��Y�c�����&A�����ʺq�}������\�X�[�m��D�_�#6�p����H�=w��:�#=Q���W=��F��Bn�eG<��$+�d�2�\M\�E����D)��cV�]�F��D�lʽ��T��R9)�m<��x�]L��&�Mg3�Ch�C���*yE��d78y}X��ч��(��=��5�G'l1�bU�η�]�\*�k��~�	#���w۝�v�v���g�6�hs{�8b���',X��OP�� _+����b|F��FD0X4���̌z��AЩ4;��-��U�Jv+U�
�gp%��l�ef��b�[����a
Y�����XPq-��W��5���?��u���g"��g���=��_����3�q�E��(%�0ɭT,��ܽ��e��g�GF�Y�`8.����9�U|7����o��02�℡� `2��f�f|,��6a�}�TS�B� 2�ho��C���`q����&vB����:���f`Ey�?홡�3?l|�~1�̤����:!S C@��3��Q�P�C'�Z�;/��D���B��Yj�OY�F�oհs��p��%�p �;8��cW�<�p4�G��ax�[�������T	W\~�"􂂜7s��D�j�[6RX��q]�w�z5}q�t1�q�b�ƍ^��~��-�ޖ-[}�3:�SO}�	fk;dq�:�L�^���,x�� 8��'7��ɟ��e��@��a`��ܺ�n�0y��,U�Yߟ��*�.������;b��L�f;��X��!���q�8wx�^l�Ӷk����+���e���_oi�C�����}�Mozctn��0n������(L�Aks--c�O���L���8;K�v���=�L� o���������~~i�o��7�r����|�_d�䌤���}z��J)F�ǯ�%+պQ=� ,����^��-<� ���b��S��2�E�F̑	��ex�{���'w���Ht}���Le���QY5C�nD��qT��Q�$3�ZR�-�L�;ε	l4�'Z5E��������R#������֛n�f��,�R�6��'>�s�s��y��x;�\�n�������I���w�Vp֋��)Pv*gQ0�� P�� v��r>���%+�;�5�\c�/�<�h���m�	�U�x7���:T��jf���g�KivY�&�ɏ��~,D�{vt!U��s���!�o۶�oÎ�(�>[$ė�7YR���t	���[c�w��<�8����D���011bdd�ੁ�
��Ox�}߽��ϋӱ�^�֠Q���z�����h��eZ�,u�s�''����z���5;4����[��]�K�><ʫ(MYDQ%�o��c���D�~:�`*��o@a�����PjQFk�j!/ȝ�yAZ�ژ|��ьBX�$G?ph,l�8���+�q�����L�p0qK�,�Ŵn�z�Q|�+_5k��A8��� wv�k��7��󜚝��l�j鮐��pUֆC�Q(�iQP" �g�t,�yIu�3{���Y���_�d�-N99�/1(=�0�5���B�8T�ď�o4�Σh�G����l6��P�Kk�Y��bd�
�^J%��k%��2�j��8)>�M7ߜ�9�ᡇ����~�5�f1�)G�����kAYR���4�f����7����Y�u��%a�^���9mbj�c)�t.������G�"i�ɧ3��Ӵ%S,P�bN\�YG�����������|�)�D��b�R�����İ���[�LŹ�V\Zd��p�dғH���N��l���
כ#�Ck�<�ҧ�y�e�F'&�
�+��zlU�79�%ErLG)[�V�z�Y���n���
qEW0[�#DИ�+I1���)�v�=r �p���kV�E����}�/����'��¸ q)���HN<q�M�ott*�5f���?�#ߗ%��\�J�2�fJ�Pj����d�F�rb�a��v�}����˿/~�K�`>�_���
;v�X�� EfTb{�V��L��aP�E��6i�K�pJ��xJ�6�=�#�?�����xz�̬kp����)�Q @~�����_�zx���nx���>����0o�p<�A�^��Q�{FG�MaS�����ۢ�zC�
��i�>Kɋ��[���~�'���|Tj,��ʔ���ga��|�+_n���|绦@��ǌH�rg����"�ܹ���U���j�k�ī��%io%�������	qS���_�]�������U�V���]�z���������N��x[��n⼅QW-�J�R��H:��v9��B��Ւroo�H����:�h8}�Rj�����2����U��OFA?��O��7�&�>n}���}a)�uS���F�p�������o~;|��
K�/6�l}}z��
+h:�ZXAN�v�k��<�\��N$u
l-�4%N���be�5'�UP��;�� �,�B�p�z���^}lCX�bUܹo0���_��������N:��1��t<>��Gܛ�[vU�c����W�%U�����B` ��k�q����y�UQ�ڠ~�O��烇�(��\��3	iHR�RI5���iw�֝�?�Xk�}��*�u�|'����Zs�9�?���?������������ƿ�WN�'��D���}ޛ��7;���K`�YR4��=�V�{e��F}\.��A�=�e��-��	���f�����[� ���_fk�|x�lܴE�{�=�ۿM�g���2�>*���VS�M��NS��v:�<��sM�6񳒇m�DɴB��Ƹ���eҪjuMb9��P��<��ty�?@���K/����F����0Qe�n<jm�]5�=3n>F��nt �ͨ�S̸P��+�;!סJ�U9g�V9z���~3����a���r�ŗ��� �I��q���sΕW���_�M�>!�;G���zp�>�z����LO7{R?U��3lP*���H=̴�)�kږ�2@��`�1KͿ���"HQqE����%k�m��������{J*R��"��������;���At{��a_��*VqTc�>g�&���t}n�ϣw�pg�ndZ'�X6dң��z�Zv���iѤ�H�F�"A� u��ʬ�.}�i��<B�r��%��<p���4��!�@$@]k׮��5k�-�Z�Ŋ��ѧ���E����y�ҚƟ��xZ��"�;5m&nLV\����[�"O�t]�]�EO��=���X��O��[d�{�#�^w݋�!E.ɶm[�ƽ��rc�r�)V�����B)60_!�TKT� F!S���X��z�+^�u������;�����������o�,�w�����J�6�R�ݧ��g��*1���J�`֜�,��IІTNca�nV������vR�R��z�A�s�a��y���i�zB�u"p������%�����1h�w�{��ݛ���d�T+�?np.�q�����_�q�O�������S�M��z�R�1+�`��)�����F&�=�z�����A�.����=������	# ��]Dh�V*�s�i�!���CO=�����^b� yp��,�O����}�r5_��<�.~��!�	�ј���k(Q��`���悔QIΧܹN3c�k��C����.�8w]�9<�補c�<�jf����Ytפ����Z��C�o݋�3�K��Q��}�6Q{��+�%;�?�ZC��?�?��?8�{�����H��%1X��i���Z�^��~9|�ԧֻ/q�-�ju9��)�"6�P�&��hNfvt�F��y���L�FT�)ߒC)'�11#W<�*9��� ����z�&�je�踆�l��1y�ObWS� �f
j��a����L�j��ǰ������������XL7��䕦�3���ɐ�MR�a����S��Վ�Ϡ�*��jh0�0�pO0�<Dv�I^"��q��6Mt׌
Wceő6fV����c0ȱ����8�kC�ٯ��/�3�y)����˘����J�7�ozӛy]@"x*ݿ{�]�B��9��os�U�f�T�Ņe_"��������ܭN5�g�0>��j���_~��7�"���F�1��GA,aq�v�cz�:i��t� y&ĮK�,�k�qAQa���r��,O/��!�c�QIA���K�ґ��i�[l�'n�gy�].;v�/�<t?�RR��AC�:�!��q��I�������or7�J���و�NTs6��	�j�)\�Ehp�6��S��B��x��­�0+���R����%"�]_��� #쁉2jR�e��6/r2�x�h�xm���O@U�תmsؓ�����3j��6�^pq~��vǧAU�C�&S������� z��AV.���8|&� td�}��~�lڰ���qm�
�f�u�Pn\�L����~��{�-_$�> �rk�t�c���O��O�W���%�{�keZ&�\Ag@�'����u��kš�h�����Q8��,�v�*a̭����z&���睛�鵵}כּ�E�lu|�9�[;.�H��-�r���{C`�^���9��ꂉXO�l��q8������ߍ�?@�&�͆,7�d����vx�˟-�=���0:Z��,��8'�x:�{�^��w��M�kDiz�n�h��J6�j�^�o�A�g��,���vM��\�"�_���;��[��\ �������3*2�u[�W���q��j}JeϨ+�x	��J�K_�-/���`��iO�>np�Vp����}���C��}w��s�bh�.x,��B|��[�"���7��$¯|��tC�_����~��-����>��~�� ؊�ɓO��9�@;l�k�/�nx嫉�/��<����#_��W�v1˗����3������8�1����n��� +ۍ�Q��~���< ����#��G��"��r�ʍ[����>(}J>Fl�qlЯ۝.�'��@�d"U�C9����䞹��xp"���ŤHiht�G�A��p���Y}jF����������X���5�ng�0P7�玃�;=��}b�#��sH��qN�8�t8}�g�������(�e���� ��I�/|}�~�^�.��خ9��Fŭ��M���wx/�{��!��u�ƒ��S�߄��:
���>�0��o��I1c�LLxJ��c�[��!��B����l)VM_��!��S�!��F)wy��4�ۏ~���o�!o|�k�.������vht������^�_?��O3ۄs�܂D�I ��\"B8�pB~��~�� �����_~�ר�r�3Zk7�gp>.�F�F�0cy��F�$ŝ3����3iM�c�Y��\�u.���7׼�D��,_< v�u۹%��[�j]zh�C�QU�1^Q���nn��;����8�1De�s2�s�#'�E�e��o����N*��ʦ��-��]�z��x3��WK�DԺ?9!����M^��W�`�"@V�N���ŋ�����_�=��R�2��s2ux����:�+��bZӳB��ah �j�_/GgrN������ơg��m����XD<֦X���j�,��4���h�s�ؘ�ݴ� �.�!4�(��Ѽo5��_r!�����>�7��F�`B��~��F1d�6o�DWLf��B�_[�V(�eY^0���s�k�6��/e��7dg�ۍ�օiʶZ�Z �_�q���nz<p�4�cnN���إ��VM�_1��m�"�������ݸ� 7Fw��Rנ#k����,�(�r���qv% �"E��ɘg�`ɞVjS�E~�w��O�����}Q��=�M������]aN6oZ�v�Yހ�s�=Xϻ�\{Ӧ-D$����f���⑋������>�&��R�J�3pb �gnM@r�qI��:�f�vL�y�t݁�h%���h�nnV(��8�=#��c+�4��_��Exn���j�BqN�]��i���+����a�) Q�*������7>���c�� �~��y����B1���lڰ��Ȍ\~�3߸���ɳ���.5����D:��O:@��~��σ�X��CLX�;/�I9��؄4�O2�
I�K۶m�) P�G��~�K�d565��gg�I�ݼ����]�χtc�� r�'� 75�ƤӦ���gL�&s�-Ͽ�2���wP�y�oC�4eA�i>Ǭ�J��%�ݡAen��8�i�,��2��I�c��6|v��Y��[/u;��-����_�C^t��r`�~9���ik@�.%ï���5Y����_�
NBUu+�c�;��F'��jF��.]Q	lq ��i�v5C"�l֠�Z$�9(s�xchq!R�`�?�y��i�Y�ӯ�)���09N?K?ǴM�;�T?�΀��Q�ך��ԻT;�{�L�,�BPdP�a@�a��G��M7}�m.�<E~���q9o��k��k���a�MOΐ3�@+081�֯a�I>!c��,����f��ͥ293��� ^�����������wG��*	�	-@�qjb��~O� �+�g>"�H��}���n	Л��d���.�`S��r�3�������=l蕀I�͘�H42�2H��S1�T�µ'9ά�}J��(?1z0���@1M��wI�s��y��ط�f)U�ϟ�����/rë^/��_�F�5��$��ei��~l��|��ۨ�V�ͣ���\�0�j�YV���}:n����!�UŮ�	���y��sU֟�]$/SH}��F/���`�����0����E_F��q��������2:~�y��0D���*���*&�dw��(F䅀Á8�2(ox��'�~�����G�������������hP�C\�&ce�'P:'����gg���x�;�)o��oe����fyd��nq�a��s�n��'I��KV�����|Ź�߹��ַ�K�~�N��P�r�EL��@u̬��2�K���{�����/:7X7��ܹbSw��ី��I7�8
�>c'c��@q����)��fZ�%/v��xp��a*��z�9w�+gՠ0m\�m����i$9���OC�
p$�
w�1g�+Q_f��|��r�k_!�>�������t��);~C�\.&7vD�Q����s<
�KW�E��O��ݜ��j(��K����kL�?��?�.������&t��{�QA\�x���c�N�}5���V�~_�ޅq���=�zXq�u\����v=��lZ������3Z�X��(�C�����Ē3��ڙ�В��}� U�EA@(�@����w�C>���c"�Le�/A0�.����o���x7��KKtϭ����?aս�e�m�[�m�&���;�����{���'�y�,����E�����[�!O��W�n�9Ca�t�Fi�T�3Bo��È:���̺<E;�rZ�L�;�F��r��J{"��:��udz�&yb�!y|�>��%/u~�.�#���]H�9������+�	z���|��tf��<C<� Ĭ��D�`�zc�z�-3(�ܸs�{U�p���a7Ҥ
L�	��>$�E ԇa���ˋ�mHL�&��f���&#�I��U��{7�c5��}f��?a�����M�����)��	H���]�CW^E����l�!^��#�(k����m�0|�C�x��h����B�Z5�vO���Ĝ4����zx��rb����V���v#�lݶ�U���o������� ���m;�54�r�k Ku3=��N�J�V�iV�7�;�G�����+�ݻ�&�u�Ԍ�!�w��Dޔu�Z(���;�Υ:��s�,�H{J�TNs��F�� �	1��ߠU�3�P���T��l�X�{��='�����(��Ԛq�)-Uǥ�����E9������E/��o�,#҉w�hR�[��a7�D+�ʅ�,��iB04�ӃJpſ�8���smr�'�PW�:����
��?�AJKb�}�k_Š3����<kI���8,K��z����b0ᵇH#�����(#4<��yG}��"�#�	m,���ϑW��U&��Wog�����b��4�Z����^(�v="�������z뼗��K��	c�wh��s�]tev=�Y��qR��X7o�O���ʼ�S/��%����+�﷝��1�=���,c����2z��c7G�v7�^	�n��4��BX\�5k�_�=Ɗ�44+�i�1�ٹ��K�2>!�?tk� ���&�w��S��,����$���A��K�(��q�y�wq��P#N%�5_��D/L)����=x�lq���C�q�6�?�_n��W�G_��y��������9�T���h4�`d14Nz�5W�Z�ND��E�z*�L¿�F#K\�.ϐ>�p�wŘ��q�?@
�������E���!䄬���_��f�`(̾/V�&^�>�a5�e�������
���]�P�q��,vC#���w�!���˿�0�PU[�~-E��;��KD_��m�C��Ape�O��:�ɠVAiͬY�ߍŌ>H�g��#�C`�` ���,��s�d8�U^���#��4� G&
�K#%��JwZI�1cA@�瞳���V��K�T)�.�9�<}E�������R��Ps�dƹ��:�u�Djc��ǚb�Ul,j�5���,�_�֛r��̺<���Y�UH�}E(.ӈJ�Vwz�3�ͮ�ǧ�{=&����뮗�7��GT��M����2��f`��X���W;���X4ʨ�;8��\�'7(i����Р��l�ΊE���\샩F���0>�m`]:�q�y;��c"b�k/���}�}����ژ�Dˡ�X�ĸ��V��&�v�J�Z�:c�ѡ@�w�(��U%_q�s��-�E܇�B~� *B���k�e��%/y1&�B��{!+��-[7s3i:�x��K�������ӆ[��wk��zz��SV����1�fb�Cc~�uג���|F�p�������勷|A�q٥$�=��>��}��и^OB���A���� �t���=��9:35M!1|'����879�&�U���*�1�P.��7[�bZ���O�i�d���r�ؼ<��T�Ƃ��rcJN,�zQÖu�>�������{����+�8�p���K��=l��[�.hI;x�]:�A�#$�iŁ�q���Z�<�F��J���S����z@.��Y򒗽R����rx�nR�Q����t;<�n�@;�@|�s����A˾mBc�p�4���őf����/R��1�%ty8v�F;��fy�8��V({�ݭ��U��K����炛0����������t�p��o��_�E֌�L���ZѝҊ��Kn�j�tن���|̱c"f�n�.V[ =����Mq��j�Z�����_���΍ֲ0�Ч��&�� �3.��a2Ya�=6+����{��qԀ�"���WJ}:�"�����c���G�
`d�V�}�x��"鲿+y��%��zO@=g����� ���N9w�9�vfBʏ��7���r�����H6��';Mm��:2���s҉��
�^��դ�2���ANsK  Pɱ�w�wN�|����"D��&�^Ն�7���a챝/7������_&w���t��IUXW�Y�i87ځ�[����<8$WN�&:�FR^��5t�y�'��8�-���$�B��
�o{[:��<�U{�
�b��$���/�������H_!G��uޥ�t�Պ0�yf�����y�jX$����.��<toB�aeX�d�(����3�a08������̑�Toh ������I�0�pz�a��e�~>�E�Ja�,,A5^�>ßb�n��p���PbD���J�K`��U\��}"u�P֮��cG����c��r2w�8������(�f�Q���N)x���@-w^?��>�ښ¸�x�Gr#v�l1��_���}�wGQf�	�Ϫ����E �Ŋ��@+��x�����=�m�|�^�
j��ч�c[R�dE"���|V�uB�/�2-kU���U��Ӿ���ǉ\ːp 
uO�}�ů �!��&d �1A�?6� ��!��swN87��y�*`4����^o%JME����XU�3Al���Y�6�����E����"P��rpR��\^��'����-y�5ϒ�Π�}�!7��ޖ�O�8�x�CM��ě�ɆI����&*�����ӽ�k��񣌈���A	_?x(��DsҬ�I�V�0,�A�4x�_C�ĉ����, �i�zM���.����ۿ�^@]x�̡��C�E�ׁV���liu�'0���������?��?˛��R�S�t@��G<��@��}��v	,�Iwa�ސW���ٷ��H	�_ђ�	m�s���� ��Ł 3��ܔ�rLg|	hc�\g���t��2t}�k^/>�Kn|Û������⽆�39Y�RU��k6����k�G;XE6�bq�ŀ�֧>��hh����7��7LZ�{�X�	E�w�]�;5Qg��8�hT�Oc�������'�����^Ine�!-�R��c��йr3�XOM���w?A",lG<`H�S��@��r�5yƙ��oN�g��'����� 9��V�A���K~W����#�m�zy�K���� ?�����������=��lȵgw�lXX�ilw�]-d��D5���a�2�>��:��lIMIa�$?z찛8hy�&,XY�^*�N�1%����4
pC����������b� "�.@�9�@6�T��v���N~?�7�ϰ{�ټi+?n�s��ܼ);2KX\�g����܉<�h�8p�^���1]��u0o}ˏ��	�n|������{��gznk�n�Ĕw;L�\��h�a�����{�".��\��a�06����<�Rovp�Yv�]��}'��AZ ;S��g��l���	T�Ю�����ss�c�q���I�y�__9쐅��;w���ܙ�m]{�Ke���=z��y=W�:�k�ot(o�tF�ȱ9)7��)e��a��b'�vp����[6.�]M��8*n��3N��)�{+U��nG��W��r��ϐ'�<�\���u.��Ψ-��G�m�9[�sײ(���M16j,F�PJ���щ��rB0�@R�u:Jb_���xt�j`�C3OH܃/�u�6.t(�� ba!~��{#�c�_-�ġܼ�[���w� "_�ѷ�y�|��JA�O�ӌU`�{6mR�΋�{�<��.yӛ�D��-7�ȦRW�����4���\�����K�7�uF�կyӲ0(�xÍ��0�	�
2i35������.�k!�d�����oY�3pX*F��̣�ؔ��ؗ�1ӳ����wk�ϱ,��Χ�!��{�1�d� `]v׆�OB:{�Ĭ�k#���ܿ}��nn79�`�p.�=w�c�������JL���U�������&�K�J�Ǧnt�!	95WMJ��P%��g��#��N��4�P���6"�17��X�P���:h��"����yϺT��w�x�Bך�� �M2ܪn,.��0�4��c����
ñ��៓�X4D�3?[+=���2<�y��L3�J�>ȦW]t1?�q�e9��:$xp�3] Ō�zj�^���Ym����&�]߽��=��>�Z��"�g��Ppy�_(��������m?!k�n��O�$Նj�b�c��� �/��84Qd��'\���8���/�����O��흿|#؟���]A-?ЅlbS f�@�.-ˋ_�b�(v�ߍ��q c�Z��#�z�����s��BC�0��LC��R�q�Y�Q���q|���꛶kjz��)e���I)��C�'�	p-_��K,�����losk./rs���jf\��v�w���������^��C�NL�d>�驚����k.q�]�����C�B�Z�ŪG�lv�������GtaP���To|b\Ʀg���\v�5Rs�����k-�����
i)��n���������>������2&�y��x2ê��]iN�oXK�Z�@P&w�dC��w�UW:c�q�����|X�ؙt�n�&;&-؞�l�����@&@X ����y�=K�*�;��w�eJ��7��y��[�h^y�k�c��� b�`�b���Ja��g>�P�{���$7�n���D��-yӏ�š�/��*w��+�)�W����E�V2�"@v ��t|?�,����Ÿ"^�����ַ��9p�0]���r��48-��,_��cQ�Y�Z:Z������H�7���qu�œ���!��m�Hgޭ½G�E���{1>��Z�����7���.��k�T����l=g��;|T�:xX�n�&GO,RN��M��V�D@y��x
6�-Jԏ���P�^�ˋF�ІN`h��	��eP��$T�j���P�j�%��G����g^,^r�u�ؑC,&�8K�ue���M��X���c!�ر�<�d�W"��kyNvÇ��E*��'�:7f��|�	fi��@����}��t2 �lf֪����@�Qp��3�8�W`�0�w�8�����{�5)��Vn@a�:���y�q��n&�		��v�..��_��_8c��i�Z��a�1�0���'Y���1�ѡ���^�Ͱ��E����w�E�������a�'�xXE1\;�������<�>�ws4=�_&�`���l�5d7D���u ݏG���׫�Qx���?�$O�O�����f�"��w��1A�$�~/���#]�!Z��n�@��Б9g�����(�j�mMY�S���)m�����S�b�)�3�P<�����@%�i���gD�D�5tj� �i�x�S���<�p�i�������#��v�r�%��M~r�#��v���	���7-�AJL,L t���lհ��"�f ��V��iDQ� ��\a��4.f:�	R?��?���~��r�o$��}��3���k�Z4�jy�,��q�Ț`�A���ݩ]�Ua#��C����m޼���{8�����]�1��,ȎE ���q��ȴYGH|�E�_ [7o�"B�9g�6�U5����.,/iZ�����#�:rd����ew$+�˫{�Ѐ�p��A�x��ȭ_��LQT㒴���S��u7��CS�""���	7Y��:A,�}�u�� E�R9O��18C�nɹ�`A����?g2�P(>�}vn^;�7A�o�~�,.-��_e�%���}^�(7l=G&�7���(��M��D��~����h�8$F�g`%Zٷ��,�̍��5(�j�6	���x��&�(�q�C�>R�y�+��ѭ�d�ב��-oy�r����|��_�O~�c����c$X�)���XNX���:
��$3MZ;��g�w2�b�#G���W_I�ӗoES�e*�5a�����J�J��s�>=3�k�X��T��gU�V�����5 � ���*���R����������{߻�1��/~�\r�4S��s'�;�.�B��!�zM	z��E�Jݢn�Y��+����AĽ	���_4U��	��Ї>Ĵ4Е����k����KC��ޭ�����C2z�Kx_%g5��%n?�"�q6����N��җǎ�u����q ��M�Q���g]�H[etc�.}�\��H�d��RB�,��H&֬�[Α�O:�Y�Az�g�,�O��4Ns�R�f
��e{>��'w'��P��6O(�c���A�ȋY��;�S\ZY�9*�z˗dqy��V�����m-J�[JV� ����N`"������|^�+!Ya$�Z��^�@�	&j����
pԸ!���gi �&gT���Nym�b�ݤD=
86��װ�vMws���nG<vbV�Z���n�{��~����߸q3�G��o���$:�6|�r]����䝜^C�~�L.���53��A�瑇�f)Љ��u���6r%~!N��|N~�g�3Il�n�&;�9W��!�Uc
'��cDC ��;��.���]t��]Z(|6h��sd�b��W�U"ψ�J�&�C�}�D�1ƞ��O��Y#0
n�c�kX�'0̈�4��B�ubz��p���aK��= gͺ�,z��Ot�!�G����}��a�9;����=p�q�Z't��5R�-/�΄���CW�Ґ��yfJ�,O���a��bČ8�(�����Bʶ�
������D�xԧ��ާ��m�G�m����92!����v�
'�cLY�!q���\w�a�G�&����<�`��#G�c�c��1�AA�;- ;	���F��'z�^����XT��8���� ��3^�jk�[�� -��1X/{�K��G������=z�׍�0
�}����*C4�·�n ,4\����DX�"㡽����@Dl���A���}!�%�{�����+��.�!��P��
 9����h ʖ�E����}�B��Ҕ���c\��K";����j�3��a�X`�aT�����Б��%��9�Y��X���Jܹ�?2ݨ���;���9�[�ĝ�ؤ�-����IVG�I,7+)�>Xv����?�dr����L��{QxZ��w�a���H��ا@/Y�@1$��n����ǝ_�n���~������G��S{�<5�]����zc� k�M�k��� ���[��#2Cu�c��fwh-7妛>�Łx	v,Lx<��	�Ei�cn�/�B���b����ahqPG��{�S��X`(H��oqg��������ɛ�|#	G�v��rW�H���*���{iǄ�d�X<0p'��ޝ�&`��=��������ŏ����z�A���A��U���0(��oϞ����7�`���`��sK��ރ���;��[���~����ߟ�dE�BS�$�ե�/���W�^�*c܎�C����%�s��c��c��}>rT[ӢTuE�>�8v�-n���C[�"Twn�6o������?%i�&5���/���yn���:�X�;�$ſE�,,1<o3Ɇで�XϨA��e�P���g��,��J�OSԱ6O���A>��8�ZC%���;�?$�k��ogV��`?&�N@�
;���`�b �b��͂������C�]r3�J*��ZV�h���QJ�q�Ȧ�~��⚎;BI���y��/�}�{�v��3P����v�X�������=ڱ��Ⱥ8h^�6&�ׁ1yʆ[� �aR��@���Qcet}����!���E�Ae܏���ފ�4��D@��q�np>*����h��#Ӄ���$A���1�
f���;�pj�1f��(�_�T �s���v�@c�SFc�Zn���iC����<	�����?�"�Y�Qyb�,,9���6����˕:��e��5ë��@&\���թ�����=@��C�3y$�����}bo�L��ќN�#�rI��'�����o�)Sc%�����]R���J9��{1i,=���<'	v`�� �u�.^����Ӣ���o��\p�y�kDv�<���P���� ���'���q<��#����`B�P�����11
��T�u�{�1�����qF�9t���9���}�ϊ�&t��&��ZR��ڇ�q����H����lP���d��ݥf��h�+�'&-��A�,p���p�W�Ő�z׻����X*}ǎLA#s�)lp0�A�#žVf�1J
ׇ(DT�?7Jm���Ø���~`��A���B�r'��Pι� c��ظyƘũ�}l���
�;��5g��9drԍ�S��ƺ��ꁘc�檃��V��Dl���L���s"�&W�S��lug�eYθA��&Ym��V9z���qtF����1Y3��z7�a�,D��ߚ���K��5���n�g2렯N�8���e�G�q¹F��݀�v8TͲգ�H�p�V3$����D�-�?���������g�K^rkR�wn����a`�^���p�oLS�O�3U)�^3��S�a�а�_z�3凟�<N~��>�����s`���̬�O|�&N|�+ј�JR�u�A*�U�`��/�z+��ο���`�0��ۼ�54��yAh�e��� 7 �j*�e�05���y�L�\��Oo�E^�җ�~wMB�g�\ý���j?��8s�}�Q��"�=��ۜf\̪vW��"L!�Q�i\b���y���nl�!O9����/�e~���EqY"(�}���f��>C�>&O<,c��XI�W��4��]/5�EZ=��G�oԘ&J�c/�j�҃Dr����6n�U}��`�Q����l/���j�(C��r��0:�J;��1���v�Ru�Y^ G@��2����.<���5w�a�}cLe����+�괵�!A���4�-�����K��䎧~���$.i�T�X��q�j��Z���9��Đ���v��"�x�|�_�Ā`���8v�� i�]��Mƍ����SO�eViSTX���$|&�Q����ֲs'�ܮw�K_&���I���+/�����?�W���e���| @��x���ƣ�l�<�cR�Tσ�g�P��k���Ε����PK���[ �,%�_�2F�҈X�� ��!�����9�~��Nt!��P�����Y�n�3Z�4&0"0���S��5��Ūr�����x�#���ΘT}�������#R�	���NT��Tk�:t�C����Z���G��S���A��\wЦ�3�+�`lB���u2�?���d��e����C'�W��R�mf"�P;!��Kn���W#���M�`��>=#8Z)��@�סN�ljvmH��e��5�%e*���g�����V?8j�56�u4��$AOة��4��R�+U6g:|��n8x����#����du2����Fِ�UÄ��; % 3\�k��\�|�k2�?U�8epTd%�2`?�e����r����/��`��O.Pjo�B �t٥��֭�p�=�ݘ�^^���$���rY,��{�|��o�ڙ�O>��3E�k��a����`���W�"LUf�J(yp���Uc�� �&����ԧH�ꂡ��l��|}�3���X���'�L�jz񀫜�	<N��!�)�=��Or�G4Q��8�s-�Â(ӌT�K���BZ�4ji�IX���#�R�%�k��E �����0�kc5}� �)�&>ߍ�Ը3ֈ�8cTv�grfəM����RRwV�� i�&F���E�����V��8q���5(��2"��ri_�}3;��j�A3`�	�f�����i�<���G�Mk��+�v;��w�]Rrb�Q�e�"�(0Q�4{����^��v^�ĥ{�P`��RX���hC��*d)�-��4u�lX\J�����=����e�r��M�.�j�q�����v�C+���k�YB�_���`����?���/��4�{�2�΅�x�K/��[��7�t&č���-@�gP���R�0L�,��9�%���0��e� ��LafY�H�g��',N�m�Ey�% ���^^�g�r���e�&�q��A�:��trC%;��KZc��s�����ʉc�t�p�`���C^m����:h{n��b�\��[Y䇎 �MN�!�M�K%t�G����F�}�_Q0:�<�~{��y+��q\-�p�l�jW��\r����9��^���՚5�4>{�>.;����_�j��w���A'��kJl *����D�lw4{��#�X��[��՝�e)��i�\�X$��y=n⚖&(|�;�P��¢��8@ښY���dU�.L�Z��.�c�:������%Nx&0s𳸠Fˮh=g�����ݙ���UF�=� �d�,H[P��'� 0^'���;׈8(��Q�} An �?�-SB�h-�n��m���G'wO�f�g$}|�c����@\�x8d���o"7�`��9�Ν�F �4	7U�P�������v�Μ{ׄ雝�L�Y/;�m��������?r�Es�M69�8��t��Q	��ſ��='C�rZ��3˔�4q7�:Kl�����|aT|�&�&��p,%j��������.V�{�v�� VW]��M��gn�[F����������|�|�1�la$���kD�5��e�a!`�#m����i��}u��]8���E�@�O;��m�"v������V%==����? �=g<����q³w�wy��\jIk�G�:�|`A�aA��n1L�a�|��``�G�½+oQ���R����'Έ|����׼�U���z�������|�~���a�K8�D��,G����oI��A�UC�\^�{a ֐���a(�Ȉ�!.j>�)����D6C:�.�iw�!��-�,�.�%5�=�`�*Zh�Z�JI+݁l��yġ\D�ސ��+3���{�R[�>>�@0&��|	��c�#���x��hg����v�$Q���i��H
X���Ov4�V��3ҝ�n��S���O,ud��m��[�"ǎ��d���]�:v�3��H�L`l2`�br`b�.Pv`�"�*���O(��'���
����7�bX�-�V�j��:'L�$�Rqh3�b�QC-#��T/_�Љ�Yy�[�B$�k��	�ōkA �;d�P<I ��R^Xi��|�F�����*b�F�������	�s���.	{����ycl�V�.-�-s#ޙۄZ��X�$ޏr���A�Rğ(��B�4'��!���	j�..�~�p��u����5��Y&���y�olhp����^�P�E�f�y���e��CR���C/Gf�I�@�,�Ӑy�Q�A���.��)��[��<�3���2gN���|���p(V�6?`%$��g���1a݈�)*�����o/�9x;-���o~[�M���[�W\%��܉�nQz��oW��b#�����:��RX<��V�V�j�*�f�.C��eJ�L+SN�ְs�al��Y��S�t���L&�q@���ˈX��m����{�o��;�7���~��\x������K��/&��H@)��1#�q�l�rcb�˸p}` �#f�%���}z�A,^��m_�uJ�L���Yx�e���fpa����n3�d��&_��i�@��I�4(����};_d���q�����m�1kT�|ZV��?~�,fd�P2��w?+���5X��vȊn���9�X9�~�m�*W]�<�O��C��}��KR��Rm�ŀ���y�j.��)9�h�0/l�o+7��k��d��X�g֠�Ŗ#���䚲F �cz��Ǩ�4�slC� 3UŖS��)����lO	�@�-��R"����O�FO8���?Y�M-Ӓ��՘���}�1)�
L�������mwT�@����!d���Շ�(�T��X�t��Y��a3��m�MRmk�"�W�p���y]�5�xx-tX�� q����-c 0(02�.@�T��93��5~��G�G���~7ٸ��,--���3�`a1�/,�����<�=�T��f�� ΂{b��c|q_,�l�85\��=�1�l1$���}���s�{�ř����c��Q��W��⋂Q��Ĺ�z>>�< �]�6��q���������R����\��V�Ǌ��P��"�S��U�a�6������=�icgPҡ��xJܹ����C�/��;��	4����}��l�V��f���a�U׺*M�����q�v�fHh�Z�Ƀ�8��γ:)ݎ�(n��	���"�N�m����6��  ժ҈*��T�># ������X� zZvF��6<�!�'1�B���cc�B��dfE`1�� ��°�����A,�
>�13���-�_�%7����������|?ꏰ�[��l, Z�����>;��6��q�4D�]c#�������-y^T\�s1$�/<�w������� y��������i����Q!U>E�����ug�N��%�y��f8��Po�{��k��˞u��=p�!�G��Mo��3�6���ϰ�����6yΛ��d���y���.���ٯ�W�&�����^�ל�}d�Ӡ�PK)ʍN&ʅ!�5�
8&-���띸�&d�b8Ȃ��T螶;uF�'��2�������pz"��u���49-�7B�o
|o�����~�9Ґb2��%k���b��p ��g# l����k�q+O��<��69�0��7�a$e�C}*���:���=`���:�ZPBp2)z�.l�ݩ�w K�Jv�<���a�����zh�4$���9��c�V;�h�-fTm;:��������J=��ͷ��
��{xXv?u@��/Keܝ�߾@�z8ֶ��؏8��^#��*K2�1NzhD�e}}�
�xD{�R9�����kێ3�C�x���QQ�xm��4�p6�d\s�������$e�cu���N��<�^Tfaa��Ky����%�.�Iߡ�jR%=;�ܑ�{܎TIkD3V̷�Z��������i��Ƴ���k�����q���Xw�	���`
�kD��:*\�����,�o=Z���;446��6����F���N��g��5�~��4*��n��]�(��O}����� �}�� {�t�s�t7B[��{@���{+���:�u�CӬ��q�*>tP�>�$co��"����M�߁��!���[��������$A'E�k3���Q1���#�1��v=��\��@��\p"!�lko����>"��#|�9�ٚ	m��a�k�g�4��s�ܳZ�q�Jf~�����z��|}�g�7����C�<ߩ��2�۽���Њ6Щ��z��v�����.w�4m�.�b'�:��JX|�x�X ��~� ��^���>+ʫV�hT��e�p�����Q[HT�ߣ��1W���2S���i� �#��r'+u8��S���H��)*�lEjD4+��k	�]QH2G��i�ݹ����5q�Kw��Q"4=3��uA4�X�;��f�b2�>�0�k}��%%����z�R�1'��yF��h���"��mI�<��9C!u�R�>���}����è���iLA	���|�b�=(תg?�ë�%�Sz~Qn�e��l��� ���9!bn]jG�9K���x�L�l_b�J��Ѻ-�W"��Z+%7��G��Zt�D��P��2؍8�r:y�Ǫ����	;�A��Hs�b��Ё�e��;,������T�u�zc���_[����o@r.D��@v�F��@s�4~���sxlq��z7l�Ti/�7���>�>+��E������RT!�H�����u�����9o��g�5+�Uk�*!
4�* ӶeC/T�R�(�:�j�n��{%)sZ���@���r�^�ѽI�&]"Ժ!]�ش��IE)�)~�K1#�?N�7�'0.JI�s ���(N��,e��jm+����).z�����R�#M��уx-�H,X�П�"��M��U������@���@c��ݷ~�������h� ��m��
��� ;�y9�b���dJi�����dA^[�ER#������h���a0�n�	��lϫ�T�TP�O6�ߣҕq3���#�ㄝe(���J]?�+)��ΖT�	cʪ���[ח��y��><��Ky,��	���%�@Z?fZ�BQ���CMB=�L�K�{qG>��0tL�5����C6h_�|g�#�M�!�hE |x=�ʰ��[MX1�9��s]S���n�@C��z��@y�0ȅ�"@,'�j�k��{���X
�/Tv�?}�����-ݶ,,7�W�d1�qgh�0��>;(�;D�$ڎjq3<����[\|]Ywy���������8�T�Z�*(���,�����1�Vi���^G�ئxN��1k� 
���h�h�9-�e��+,z�K��o�Y�d@Z����}餧�(����P4��b��ί��l1��Ǽ89�����8V�`5VfHm���3^��(�xe�J�����#���ɟ��j0�(�=έ�:�RssJ=��k��sR	��Y��G���f�W5�q�Ţqlgm7*���oE��m|Օ��P���\���/�F,�-xܸ8�|�	���(<�S���wZYEBS�i:ymW�c�"fD�[=�@��:�)eo@�܌�}_�\b� �L�R��2�3@$��+����Z��V���`h�f���RM���U�X�V)�%���v^�t�^�>qo�>c+�0b��]�kh��c��X[�=��ƣ����;�4e������x��{r��� �ÿ� D�U�����"bK����A����bo����2	�zl���y�4\4ʂ�RF�9V]c��w�!��*|��NT�����D*�kw5�����S.0%��oH7�j�i\<FC��GԡAs�g�>�z39���4��E]�X%:��'����$1j�jZH�a�̟�(��,b�pNs?N��0�Єp�h�C#�A��7�2�T�S��bO�~�����?��T��z%nG(�K��~o�����K.�D��MJw	|��8Xem)�pe=�߰��Kzs�Go[�&��Ac.2A1Q���A�'Ӆ�xݳ,��*��E`��Cs�6p����Q�qdDZ�N��֣�S<�ŉ*\����]b�j�� �{�S��(��b�ad7%�z���XI�%|_/S���e�Y32���
Y�v�ͪm(�����@R�V�S�Ph �?�>�ny{VrZLC�1^��'0�%�������Z�*�� ^�̌��[�y%p{�n)�l`�MU.�ӺZ)�/����5jwRd##�.~��fXS�"�4�|�P	�[��M�j 9J
�/M���`1%^*�sJp曥#��3/�N��a�<�0+Q#�Ͱ�q��m,���'������G�=�����T���#Ls�.V��x��2zŊ���=��q;
�M]���^]��d��MD?�J@E�߁�S�r���ym]sK�%_�VO5/�4�\�I-��R@����m[��L�FC��I��+@I���6��d:֪���0�@uT��ҫ�p�c8���r��RÁ�~�v�@J&2������
Dd�l$g)+6.�]��|$>��(�9�HS�g�Jp�"w��hl:Q��A����s�#��E�����8E��(�`s��gk U�%�5c��֪t��b.K�����_��9�;aa/c�EZ�7��<���_�G�3�}�JI���+40�,(0I�?�#��L|Q�a�%����u��sJ�a�#h��lC�`-U��������_������MA;0Xa �޽�u'-���#5�q慑��W�����Ʒ��q1��� M�^���m'T��nw
_�d��|��
C�o2��6l.(	��c���7�{d�P�b� v�A#7u3a�$�O��CG�iIm\SE'��D��f^=��Vɏ�ݧ�˶&> ���.�B�i����w,��b4�(~ч��M���y�yg�?c��������)�(���t�\>�,B�3H���������H�5�>�9��Wf�B� 'Fl
pQ�V����ւL�Y���%L��]��Ƅ,X�=E�p���v���Ϭt�M�RC��n_�4�+�fS3�r	�@�ܸ��rS=?�H���r��6�󧲁�K��1c �r�M��� �fX
bX�7�����
b�����p�ϼ"��e�m?J�ߌ�����2`�d����_�u{r6�	Z�����M�-	������d:��&8)�أY\3�&n��R�ш=�M}�z㙱�r41��	���Y��QQk:0��Y;��_�Ĕs��dA�S�+�L˕��e�\K����Y�r7ht\'dˎ:F]�����!�pb�D�R��y;�`��s#Jꦈئh\e�i��{l�?�-�*�B!��c���LiW�#&��q�V�y��b�btI��D�y�+b2�)�_(���X�ל�+�x�� ���㏱�
h.C����$P{7T�s�(٘�O��&�35��`���q�Ջ������a(òAF��#h�枡�(��M/0m��oՌ��AA��#��1��5l�`Q[7H��_��}�n�����d%>����tSu�F�&��燓&$m%@�<�(���6w��c�㓩Gə�9�}�°X��py�޻m3I҉Z��.5z=р����b�^j�[�b�����$^ih�̑;5��g��0.�`qS50S�['�F���XCk��}R�K�\}f��[���9{�DA�ߙbF�������Βs��(D#Qq�[K��ַ��1��\��m�0}Z` ,��7���O�AWD���E��*�'&&���-U�=����;~��x��k�08���P��������b�>���`�5�
i���9ّ��2�(�mG��].%��N$�V(Ѱ��j 7-�5�:;�E�&�O����OJ�$�D	��K��� �C�7��&}0����dy�1*u�hpUb?o<��q�,��؇b��8��rqWZ���1�6S��Gd=d1H*Z�jJ�p�vGB�\����m�,������D?Pj | 3R�ַ$D3��h� -�7�̘�ap��l�We��X]�D��#4;��[�2]��,q��E�Y"�0*�_��q4��sI���t�a<���s��D�}���wR��H�E2��k�rYe@5G,B{	k#�zm�Aae����jcm���Y[К�x"Y<dP�5�!(r,E�<M��gc"�8gT:��B�"yڽ��d�VC)+]����Kϲ��
�]�)�/�#ՌM*'��4sAe�Lb(��Р���QY�+b��&�<7��*+cqM���j����6oo�������$��Rn�y(����*)�O�C�qfJ�pgXq�i����_%M|l 忹��C�<0l���-m�o@Ɖ����p�Z�,�&��Hs�D)���c�#�*�8`��gm����S�@�mb!�>/�ǥn���T��R�F-p5X��w��X\�q𐓗�S�o��A\Nv���.%ۿ�� �bɢ�Y�x'xD���O�i�x�퀯��Ex�e�L%�^g=�C�`��l�A��Ҡ�<Q)��2RP<C
��[c,ް����zeງ��j�mNf��~6㺈nNpoB�~�����noB}�.Ql����@l(RR[��}��E�@�-K-Hjj���5lB����L2���mG��p����g��K̥�7D�/��l�_��ŧVL�3-_�APV>pʩ��#�N� U�P��6�.H:�űyf r��Ge���eb���(�8&K��X��PT�����ԑY,����!v���|ΐ�.W��u� ��u	�9�UAr��%��%���+�}��$�5�5Z��{0�q����ܧ+B1�֠LA�"��˔���<x����6�&�c)�E�Þ��@�o:H�7gq��/��}��2ă�;c� ����X%���y��I����@���sg�mK$�B�q�5o<�>P�i�}�hpJzhHOm�27�bQ�G\���Zu�O�h&�b�]�=���d1��b�D�uP�4�*Ag�7V#\�H�Wd��t���7�1���y�=��a��D~��������c�/E�����{����6N�@�`�V �, �料G�c(y�d�3�F����Dc'"�1��(��@�a���
� ^��I��g�f�jR�>�!x�\����,��Ü:y��b�y�������~zm��+��������I�4Ү�nB7�UQ�I��(�@u?E��W�Z��0&���������@��*��X��xQ� ��B0�G�k����8��qwϰTX$h��Q��j���5
���,o`�VG:0��-5{�׌���z9�w�=߂�,9�[�KRi�2����g~�dHnJ���8��]*{�G�a��mJEP5.��tC$_;�9�<#Yp5��y� ��1�M����,��8�i�3�z�G*At�$ݲy�4��	ݴ����+���_�7q�]
�w)�[ˉu`t�PH�ϔ40A� o������D<�?#/����te�4�.L�>sF�$u@ˀ���U�n�-K�ݔ~�)�~��)T�j�bws�e�M/G���Rlw �#b(�S��ǖ�*v�\�9)�s�������9�AL®�2E��i�hZX�䢨0Va�we�m� xÍfTŲj��4�c�ı���C,�Ȥ�Q���c�,�H'6-�èO9���!} +����y�<���|��K�ЧN�b�ȘF�����K[#a�8��P섴m�d"��[�����饧GD9�Y�.2D��ofٌ�X}���I�ˈ�(��(E�������@��Q}�7��m�F�1���H'{�w#Z�T����}�P#�J��&��EO� pBh��x���W�٥H]Nr��`�k9��\�V����G�2����]}/��E�˿�V�2�Z.��>ߤ��*
C��~7�Ú_�煙������q0`R���0��%�s`!ω�`����(IL�8&�ο��E@��TS7���EP�KU�\H�B�\������d��°�h�Ӻ�Eq���G����&G�Q�ǿx�܏,�">f�{{��m6�F9F�<��-�?����N��V�G����3�����O�)n:��=��(�SFm� ���=���s3,zhp�1�H�;����(dH2) ��P�`�1s�x~���i N�X,是)��#㍗������D0<��T�k�w����$��Yn�K��x)�d���j���t�;*
��N�-Z,Jס�@���
ur������5�Z��Qom��AF�ktGp�&��;oC2\aP�˨�
]&S�7�i�b��K����d��]j�����
c2==�|���4Ӟt��Gj�� ��q������X� �t��9d�҆�S�`�/�_��faC��G�Ѐ!ġ�Scb��
A�$��д'_�%*�g1�6�{>�-�󩨾�����&tԪx�B����<CϿ�[j�"�U<�$6�.Һ
�s���I'��%�%h���]�_����L=�XTv�v.���7��V�D���ow0�_s��T�k�R��ȱ���Mj�Qg���^�<o��-�6D��dČ���̄�ݚaWG�re�d�o��^o���+R��G3ֳ(������ï�2�����y��i��\p��?� ��)��M�B�/s�=�_�򾗀L��W�;G���X�*	�6b_����!��V0Xel�J}��H��X"=�?Іc��i��X���ş��Y����d�r��?c�}i�{���X�o��24ʲ�X�^1hP�}�	�@f`B}G�w�f6��&����0S�1eΚ}I��Y���~�y�L_�i�)��t�]+�'���w�W7�ZL�i�zI�7o��c�5T��#��H�g��b<��Idq�B�05�h���O�8G������c�q1
��<��� �B'�nM�I�xN��#�w����MzG.��y	�׿���YWɿ|�f�[hʖ�9�\����
@;}jW*H�OI���Z}	Ҡ}��{�t���Iy�LNOQ��_�"A*�y)I�r��85g��x1���B���֯������(���`|����{�iؓ3Nl�ɜj������!2�?�Ó�Q��j��(�����}��Y���6v���{�殺�����T�!�ұW���_�~�h����c�h$� $5��s�)��u�ڥ*3 �2�hR�H�D�6�҉j�i��+Ɇ���yx��}�qپ�|�z]���|J��ؼ1�G�pI.{u7��6	�}By����o#�v7Qc��+�1�E�մB�$23�`��%����j؂����
���2��.��8R�>�������E/t�8z�%���ל�h����!�K���	�J���J�5Bj���:w���^_��5[lA~L}b\J��v��;���	$`�	�3�>(Y��Rĺ����`�ØS>>CF}�PRב�F����ӡؔ'Y���g���Վ3[�SN��v�r�-�N�ib�z�&��_{"Q=�rB���(��a�;R=S.S��)���zz�q�r��0�_pIG,G*�P>���M�j�v��¸)��@h��@�ԟ����,�H����
�� ��oh$V����FQ���I	2�Nʖ�Q�VQ�Ly
�U��v�X�,,�te\N,�ʹ��_�����Q����or�w�6��켔��Fl^�����5E�v��5P��:@g��n��%� 2���# k��hO�.�k�R���i�APL�n�8��P���v���x B�~F����������D�)�#)��q?����N��!��ZR��ճ͔�}��j�8:('f�iP�]3\���y�[~\^��3���tZ]�CA͹7ǎ�-�i��snf=�ݽiC����%j6s��yl����	�OOKԀ�ac�vh���3�ayC��~����������h8R$7\C;D���aqn���n�۔N��(��9�,�	Iܧ�U��?m���N�,��`l�;d���fh0�9�_��.�"��M ѽ�7>�5u��ı��4h*}�(����\��̼ް`'��?o�,2yJEj:����r�0ӈ*�hAg@�<.���|���2�6�w��-7y��]Q�esmh����\��Y�fF6���s��#�>!H��Iyb�>�/.H���g��Ή�}6//U�ql�ȍ��H�k�����(IչX���[�`#ñ��k��3f|��9cWRJ4T�i��9T��b팈�B��Gw��	0h5iv;�-0����el�E����fG� ��>�
0���v�299&Ks'$rs���cl���+��R^��9۶��8���s����3�'d��)�6l ��Ք���G�����Ԝ�Sw�i{n�(�젙���j�)�ǝ1w�\�h��E�N{�;�f,���A���2tu��pM���x�G���؈1�!�9[=����3jPJI�w;�WɄ��^���V�Jz��h��v]�.-����I�q���4 7�NΝ��H��cu��m��Qp�\�I��a�d��\�Ǒ)J�>�w�b�y�b9�B��g�H��u)�����*]����ӫ;����&)�S�Ey��M�k�yʹ��)�E�=��h���VY�v���!��Y�c�d���\���G���2^��&����L�g&�D�L�\wK�W�V��� ��h�<]�)��5��E�"v��+�U�	Y�(.��N��� x?C!d=��?%�T���6*|-�yjD��֢�M4���O�����E��J�����yԔs���k������g]-^��95����ƾq�))6)���9�Z���gš������ƖC.I�ί�/��jl���yH�*�Ǥ11I����Wd�t��<3f�b��ʟ�����pF(<��l�ꪦ���m"�z�ig8��8�\�2��R�y�E��+���8X�m.:�6(�Q7��O�A]��w��Z^�e,�6�:6�&t$m����&J��T��q"���r��4S����>��FQ�V�r*yp�䮤�`�57JF�ꋲn���^d�Í���-&�dV�$?�k��شCU_0W+��,=,{��wK�VRj�[��[��,�� �r�)2�Vd��Z��̽�]e�>��O�ezf�+!=B/R�"Q�������c�����ZP/"
,A�&=��Fz2��zz��[k�{�9�Ѐ��7�̙sv}��>k�g=�5�$�p�Y"���S.#����q��hT�eꢝe�y�9B),�M�aY��aj��+w��v8	��,������|�;��T�
J�T�՜�&Ǥ�s܍��x\I�Q�М�����!&��~nY�Y(���ʤ��K�~�&x�d�8�'��=����'?���j�츸N�۴Z�R�)j�zi�".�!������(��d4N���"��d<��0��K%�-e�+����dH�ᐬ��Ā8Ը���j�YI�A�q4��l��]�Q|m0���q���Y��k�vHu_Ԭ��>*�jY1�7�8���새X3j��V�7Ȅ4DйJ�P�V$�K�#�)���N�pG9W02�\2�,��{}A_$r���Qs%C�*��,Ƭ[����p�IHpա��f����5�c�Uul������@aWp�F&Ԕę'.���l`y��:�b��é�/Ĝ鋑�ɽz�Z9��PǞ�~QB�����IQ����}��=H�!��T��P-j؛̣�~�T����)�IS&�J�#x_@�&C�P�A���Y<�������P��BpmF^�."�M�������ؖ�ӫ%1$���mխ0��dwF�}d$�FEe�t�ī���\:!)���Td��l���KE&k����G(�@����	�X3<zO9G:��|��L�G��s�ı$7FGS(�bPB2�z�]�xn�+��3+i�
��#���E��ۑ�U՞h�Y�~���d��헞�B�-�kd�%�R����n��je�c|���>[�r`���|�g5��F��_�+y��N���T���A��,iVi}aB�6�z�� V�Dô��!��4Y�F6[,��V�C[�J~�ۣ�m
���}��	�f�ݡ��$�oزh ��N4NŚ'� i0��.�7�5-�kSV⊝۷PH=7A�S��}{ˈE6��g�>:�
��Ŧ�sV��6�O��a�:�ձ��#cz�g�[��0��ʽ�o�2U����ܸ��Qf�e�[�I��HarY��T%Hή�7@F�&�-�z�V�*���
�2��d<#��Z��A�8��݃��]�!8��`�޽�V�%���gv(Czu	M䫖��騉q��?lLC�ϐ +�=�98s��{ɐ����N��FJ�i�yPf��B"N���g#U��yӏn�.�ڦ����?����5)�a��P�KZ��t3i�&7�
��V��iT��&7G�AhjGS�8%��P�{����_�gQJ�𗡓as����e�XJE!*�뱤�uuƌ�b0��# �+��aa�T���Ь����~~��X%�<w�Lv�2&V��i�/��E(e�n=�whJ��&{�P��h�G�ˡp�F��V��ڽq]��?y������ӏ�	O��<mʔ���?�g�S�?𷆇�����=���'t��
���F��	9��__�]C�=���~�@�ץ��Q�'��1QLsL�Ϭ��aQa�D���׀�,'(M޳�{�C^��j�*��'D�:V@[<4I5�5,�I�`΃߰�a���p&�G�ɉtŉ�ɀi�T@�Ig	T���܄�mp=�Q/��$t�hm��.�X���X�v-2EBAr��Y���hVlH�׳��m'��r�)M^6����4�"@H���sjmjE�[�ޝ�%t����i�LF�@�Jנ�`��p)C��:�� RW,�r!� M�l#}�uAO�����-��a�R#N\a�3!16�`���*䪸�w	p���b�Pe.��l����t�AN�	��|��P�IFm�C�ň��ֳ��Y��j�2����x$c.ԁ?�/�V�[AN~L�\���b�&�o:���SuERfU!��A!ו֦��m�_|�sN�����b݉�g�o�ց�}|GW�����7���?<�7�s��R��]	M5]���I�Q�<Rf�3�0�r�q䪪�"�4i��P�MΫ]۸G��6��cg��\��
d��I�=�l�V��o�z #�]4��hj����Z���r%������!28I9F����O����TȽHf����H�9d�9���?.o��\%��
���	h��5���W��f�R��D�b� cr�g?�s.���b��/~�V��f=��$��z%,UQ��)88+h��^B(��Ɂ.ҁ��!�#�3��	3p���LJ�h^k:wn#��������۲�;�_A�c��F�hB���b�Yơ�s�]I8l|u��4�}��'4�C���~����_�<��ڬ�N�����\�_�Ώ�PF���zP,2�DB%�B��!�ȥ2d�	Js��bҨ+�mEt��I8;<V���?{�ڋ�Z���g�G�&�K�l�T���٨�$��5T܏@��t�7��u�Ơ���T��8E>Hp�4�Ds,R��ܹΣ�����?{�/y��_����u�}�rx��k?����k��������Q��Np��R�W6������&)����Qk�d�;f����R)Zu؁�1o������U[d��7ϖ�Y�D�ݏ�����G>�E�I�c��d9��w�$C_��-hI��q~Ơ��is�7r��PSL�N��PI���
e��<	E*��Ak, m���ס�)��&aBb��Yd��ع}�p5[��N�j�q4�x�x���ەC(���%w��[6�N	/��+�Є!����}
�l�>���zi�pC�&I't�I���G��z�/O��/4N�c$OˏA��]�d5<��e�������߇�c����pr�ϩ�ʲ��Jo�^�i��;% @�!ϓ�D��L����R�Jz�V;>wr)i8��%��i2(9qϪ����8����·�U��֜�����E������U`�wNl�k�VI���UL��4�����k�Z̦.��F�՜J7E���u4<���~�X0�X9�\Ƞ����vD=�>v͕����S��+Ǻ�g7���}�{~_��pه��B��~)�u�Jp�	u�i��^�	I�԰�0�5~�/ZA*A�54hG��n����UǳK��6�i��/���׼�(���k��o}��,�(!.{��A�h���~��X<�F!�Gz���.�r����-�+�ǵ��	��ZYGn7�ihn�]ʎ"�s`h�f�����ܓ��?��x�b�y244����	<���p�}a҂aD�f � ���V���'�P���Y���F�&z��"���o�!r��5�6#�3]�Bè%�� u�����~�]h�K�,�̙312�����տ�,�D��c2�ْ���a�>���i��O�G��r~�R�R���&7��IS&��BvN2�>:g2V)2ʡ?F����HFd�A��%+sw�-h�@ƧTc�����B�5ľߵ]�$��c�xV�zo,b��l��<�S�VK�HwN�e��!�y�% 9oC�٢�3��T�J�W�,#��x����՗]�/{���|j�����O=�n�G594���9�va�'S�֒�X�>}ͪr>t0{_:�VgTl#d��̱�];x�(�.	���JC9^=��k��ɺ����94F�ض};:{pz�D�鿋.:w��7��K��4�v[�CT�H�WS��<�F�&m�PI�X9�8���2��;���۾�ӗ/QU:;6j����nCC���"�s����ȳ�E�z0�%dN GR��xlFэ�泤	15�6Jꖇ�����7!�2���~�0��hz2�;f9�ﶟ��sO@kt"�L��k���?��4��N/9}%�C!h���Y��'�.JF&�E�Nŷ��c��;2(%��}.�IBoyzN�H�N���w��N3�*������w �SZE�v���Hb��r	��nP���Xyn�^)K�\���2������C��̺ɿ�g��Tۘ��ؘ�#��}o����1WLڢ[��5w���{b(���h���e�p��5�ٞ����������q$���o�^r��+���9!1��ȦRQ=�P�+�T{�#U5�҅C �<��Ŧ���4�tr}y����Q�}���-��
�����\8��g0���!�iOo?��m�C-(����ř�i�d|����wbbC���.���;��H���")���C�G��Р�Ѥ(�p�Iu[׬�m7g���LV��5�ӛ/�l�tE��=r�k_�>�%�ٱ��و�#H�V�^i��h����z����E3hb�.���H�hK$0JGɐ�	�1�;H�zg���߿K��&Y�͙AnK�ƏS��KK���%qh�
��,� ]Gǌ9p�(� �c��� ص��cp��ᄓ�G(��J�	�^ݍo���9��?��`ȉ��z;w#�J
��!	7&P���)� �jm�����w<�����*�B�L�����#j�sU-U��εQQU3]���R����#��K�ٖ� E��r�j�#�^��<����w����{p��k�wզo~���r��E�P[�T**�®��e��c���,�٘�Y:��U�O1��X'�h������@.͜y������O���Gw4�N���=>7��4�bq�����W��7?{��ON$���#d3F`<�Uw�k��j�	&l�\��<X��_�aB��s�ۀ�܂�p��w��4-����=�ajG�|�����p�%W�m���#�n���	X��'�hn��}��<G�����oۄx,���nF&�A6W$�#7� ���}�{0�c*�Q�@��cZLd�X>!"�ǋW�Gn!��G�?F,�������� ��;���$ ͏�����)��׿�=�?B�%ٚ�gMG�`J\���nd�)U5N��64 �#T��,�@qg5����j��'��lppPn��6۠���QgH�y�$��-�-0է#���f�jS�!@�yR��i�b&�;�uo9���K�je�ۇ/=���K>�|�H��l.��ODd �&� ��0��J���y���k��K�$�(Tw[UJ�<h��>���� S����4�^�Gu��q����J^�_�D���}���+ޅ)�QU�/�_�u*R� �v._�9U��~�/D0=��W��;��	�Mu��ݗ�{��vt߃W�\r/�X�/}�8~�"a�Ιف�d {��i͐T.���6lIL���r�kN4�uW�	8S��L�h��$�^7B���`j[�Haz�)F��"�3rl*�r��E$ˈ�!�pti�^,&�J���k�ft�����?�s�z:�5�Y��S�Fޏ���{߃��5��)s��>�|��a�ܻWbj��Dw���!q����A�z0]JF,���<���8ж��A��q|;�<�y`v��@ռy�c(��KIX-˓��r�ZmM�7.;��~���q�.�������Zf4p`�V�0�����~�A1�[�o�k^��maZX��[]��,M��.���#al��_�I.��#��t�
�1*.��CA��p�6�}��E� 'W�Z�\���q�͆���͓�!���L��& ����?�}IL]��PBb�f��݋����r�"!��Ac"�dN���6Y��"��*57<L=�z��7⣉}�g�ɗ��{]�/&���R�Ħ�g�m��p�y�"Lc�{�R�&g~�bU&4���ӹ>�������n�ނ>u�;�L W�,G�9�X���{?^Z�
v�>=� "�6�
6m߆I& �`ݺ��bq'H��̀mhB��S�LQ��ș����b�ؿz�k'�!8�����n�����kд�|~l�[+�UcW��V�X���#�Pt�P��Ս�E7���O������K۴��mV��Rscca���	G��8���rӴ����T;��6KQZ!���/m5�K���Qk���ͦ��VS�"�eY˔��?w�%0��g�:y*�!��4�a/8ɹb���˟D��XG����7�Z��b(�t����;tm~� ��!��q̘1��Q���������Pu���=��ڊ|jg�u6^ݲM>�bO��X��w ؄|�[�D1�Uw=��q@ύ=�}Ȥ�༳��ߟy	��˓h�4,:X� rU��+񶳖�_��d�LBYé,��D�*R�D��+����,>Mn5�I���
>����w�N����14�t+~��{	m�pԜ��1	�Ã���������������Z&^q7}��c1����i�*���'�����m�1����P|��}���M����^���Y}��B�̿�1Z5���ȕp@��Z4�EN��RK,<�7x��4�M����\9�Pb�V��.J��U�����h	�r@�b�%���U]�u������a	T+֯��1��H6������M>rVBmt�
�"b�M��;��Tm����Rl޲Ϭ|��)"3�~>�<��݂�x�)�s�V����7�� [��T]���8T�n.��՗s4
��f�锔�S���ٹ���vP�N�4� ��B&	/OL�\!O��)���I�)�(.2,��*��>V���;���	�Z�2�za�?k�dUn���p첣���W�z�K�	�0��q����y�#4�r�.�����LA����i L�'D�	f�j�L9�
��{�!�;��"��1���w����:r���U)�Z�y��1|��Gb�l*N4���|~�*CW�ת}���z���/Q��d߉o�P�m[�Y������m��'��J�̓����[	@9����w�QY�)���>���C^�uyx�����rjB+�f�����1�T�Y�4�ThD��P���+��m�AY,ʊ�cV�栢C	Y��>c�Z�&��-���7Z6a�[�F
\7��V�ĳ�/<s9�(��?�·o�Ͻ���(M.rٴN:�4���!��D0��+;��3/�i�>�v��,[�ATF����|�ܛ8!��LB&tI%3����-8��ch_+ɝp�J������M���\"�.u�ND"!h}Y�_y��sB�5+�N�J56���W��L2�-��׾��?���mx4\�pե���b�D���U�9�_݇�LmM^��;�ZJ���7dhY���	)yP*��#7)���P���7�y:��f�̼QT<6DV���B���r
��Fp3��)��>L�U�7����voikA?�H��`��߳"�5��'�b�8�X}���F����f���p$��;�~������k�F<��I����&�٭3*0�ȁ�2:M]U,;T;Q�	�k�c���E���9��nJ\
�-O��(r|�l���q��˥v�KH�_�ˠ�+�҄��?��pF�k��y�yZ���r!�LҾ\R��n���4,cXA%M�°[:���n9�h 7}��(�ĩX.4�V��B3������
Gpu�x6�p�������1�V�<��2!�<�P-X�e>}��p�OD.n��4zK;�'�z��M?�5���F�Zt*�e�\�� .� ɊeVrc�M��EC�Gc����H��f3�Զ�����y��*i��i������U;�N�Kt��q7��"CPO��Ԫ�#z<1����i`�띌G,�8G�1�?U-da�xc-[��槍�D�K�m�T�)8d���\��{�`]W�\�x<�`(��P�l� �T܎��4���3s���%�����B��2Mc���Hvvw��?7��V1��G�w(ގ��6���	���cҤ�@<vE]�K��	�����n����>�yK�GϞ=��J��!q=T�k%��
m%'��Cҡ�'a �k�r+i�ݨMh�{Л�|V�Ǒp�.�].W(�2t���[�_)����ʊ�xܴi-���]p����/�)�����E,D�&/��y�5�姿�I��k�H�*\�%�H�}�U�2�g� �}=��_���ȧD�J�$�h�N]�w�IQ�U�Jvt�}^���s�9(�N�1J��0^IUeD�8�a���?��s35�A��B^��$������'�	�Z���Hk�t*���yi�{M7Y7[	]�	ĨXmv�;ƺ��j�{�U˅�	�pZR��)�u}�
��6K,�`}�Vi��띮Vp�ac�1'����-M�/��",[�3&�$ �)�|9Z��������?Vn�ғ/!�@�2��l��&Th�w؂�tM\'�r*�R(��@��&�ƍ;�|v#�2�^7�GLDb�ds8�V_G�@���V��FS����c�!��}���^���P��E����}���~����7��w�q;&N��榩d,	M��3�.`���X���6�=OמS(Fh�� ��k�j�������m��P������p�e�Ĕi3��{�����
����q��y��Fj4M�,���0�tͻ������hR�U�zH�s��UMiX�Z������iTjC�0���t.5�m�{�(V�Ŵ�v�@��~��
��.M>S���,�S��l�VC�ix4=}�i����oжcwWXs����|.�*X������5`ج���K�+�V�\ �RJW��U��*Q������S����u�B<43tV��"�>'�z�)<����+��b���=�R�ݽ�8��)b����G�(�d߬���lZEjR?ň+_$�tZB������A�t�w���߈�c��Q�1��tɚx8p��r',4��ʄȺ�U�^����z���`�w�
,2	IQ�%b�&]���eK��������C��Oz��o�k�/���yp���ї͡�2�\�̈���K8�r}��^��T�}���`b�g�x��W��K/�ob�\y���X_p�����A�Z���#��!�e~�����w4M�� k��x`����M��ai���dۿ;~�Ɖ
0+��oJ ״Q���d���<��Y����2!X�-���ѣ�66���lk{{?�Νs�S��K��m��
X�HB�"G��;�⁈�������kԒV��U�����%V�#�Jm�t(�U�: =܉Y�ø��D��_��.|���<�8.{��p͵�B8�*�^�]��{������0u�R�u��Q�յV�\Rm\5hFpʘc6��4��Y3�9ڍukW�}0u'�,;.2j�7n@W�Vx�t��`"!�;����2S�B��3Q���)�T5D}N�p�9M%�ȁQ�ɹ���)DVѥ"���W��*\��˰eW7�|�%�����Ɗ�>t̜��x��*���|�0"�ͩ�
p�
�xe9��(J#I2�.�	Q�`>N?�$r�*��{��Hn_	.�DcSD�������rU�<:���w�z��c�#�u}�0�l�Z,�nɑ��H���}cA���WŴ�c̠�U�<�mi��,�a%N5ͺ���n�8�������lj�dP6��������|��F���U��MN��0�I&��V1#7]*Ҁ������5iiZ��;i��F�r{v	�l��Z��_Q����Ws�g�&�z׭X�h�|�G�F���D���W\��|�Ģ�v�0m����a��W)����
g,h�p�%��R��	-���u+�5F_ل��[��N1��V�Ó+Wb��iX��0�u��༷b��s�`ŋ���s+��|f�rKS�[��}1U���$K�N�>7Mx��/�ß���?�J���Z%]��O�죧�+/��W������s+7�&I�e"&N�BnI��KV�� <,#I�$5�/��h0HH,%|��~�H1p6����[��)�14�"c������ �~�e$�,\8s�ÄV�~/t2L��Qx"QZX
c(�PM�8`/Q#���I�7`���(Wi�rF ��fyL!��U���W�E��𰆬�?�+^>���T�Ҷ���<�/l�y�OJg*G�� pT���Q�����}PҜn�9���̣\`
6׏Tѐh��Y���j�a�vE����ڪ��lvq�è���Jl|���?���M�3e"Ϟ,��d�%���V!H߹��ϩ]����;S��]��x����
�3�L�1� V���3��R@��G������:�s����o��H�'��}#/�`1M����i4�|�Q��I'��q��!I�G�{3�=E*t�fQbLRH)yŪd�X��4\��wx0�����k�'��f�.,'q�9��ų�>	�M����N���݀��,}v�0xvl��?,��n�;+��1!I�Յ<!�Ed�Fz�iO�=���6K`6F.۫���˖�Fl���;7���|��7`>&r&-Y�!i�Q)g�7]R��i)��c�^�3W������������ԕQ}wl����ͬ��KJ�Cey*r߫Z��&�q�S��8_o�����Opb���3�z����#GԠ<��K������ʹWhB����c��Xu;,����;	"dh%�+�-Y�٠�^"����c�ڇhC�|��|It9��ęE��Tm9k�[�+d��ѭ�ld��e:ւEs�J$֭ڀ�y	����9�m�~2|\�Z��|��غ���/`r{�Lk�1��^E��]:�:�dH��r�}^���(�O��1�M��������#����~!�уC=8��kjƄ��{��1a�$C���b�~ϟa�G��T	RSmӊ}fz<r˺�|f-@�e"�ߋ7����~S��8jF�\��x��o%��1�Bhb ;N¥������=x�����x-VE� �J�s2���2�/��uEB�ZW�'��4������D�PńI�bL�8r��2�2w���3a���Bp�JIR�.�Z�Oe;�o����^6����q�y-�c�O�+{���vg��Ѵ1�R��'�p����PJ�G� �!˛QdU,�|	��3`�=��'���}q�ʳ��y$����0�g�_�7RXXҜq��N�O��ʢ��K�	zq��L�2En���A�Q�Ҷ�C�>J+m^�K� �}x��/鏪��V�?{��`a�HX*m�Y%������T�M��{�&T�):.ǁ��8h؟�o~�g���0wƣ���'Jb�M�eW�Ce�S�����,���2��b۷n��i��fВ��5.1���]���"L~ՄX��tH�+���?�m7��|�}f�Gp�����;�0i6�YF_�E��R��Uae�a �c�Je�{�#c��<!Z���l�����ǘ?w:�8�\�K1g�|��3ݿ9�@a���ݣ���128@H�+����tr�^X��V�����Y2�����CaT�D_t����oǮ�r���H��K�,,��>Ħ�WVgs��X#�Y�^wh�4*�ǈ�NP�@�ھ�u�~�������K��g��T���%�nkRkj��_|�<�#̔u�.�nJ@���� �/2�)zja_pJ�P�i����{���W�8c���bL�[�����[�R�	U��:�\�aA���e��k.Tr�� /�k�L<��V(}&�I ��bxt>��8�
@^��u��sU`�c�럌i�C2P5%�����m%Y�H<"bԌ�����	��)˗�q�$�^|�e2�	x��x��������`<�?M�g���&��|�(AV��-���4���Ӊ ��bn'/[��Ɛ�(Y���U�s)\|�y��a� ���x���ѹc3^ye=�;�4�L�����c��(ЮD�u�Q3�B��1��x��?�u9N��!�o��b�֭�܍�Q\w�q�q��1c�L�9(U�=��d����=�H��"t��T�'�e!�BAz���ۍ3����4�/n؍�)�H�C��mw����������E��z<�&��X$���!	t+&��|(�Dz���ڔ�C��qO^Zy�)�דAr�G����A��<T=�79�bƥq�A��/�h�L����F�,K9[қ�-���z/�����s�]�l�ιMM��s�'V��>��YO=��=��o�S�eݥy�
�V�F����&E�$�zaـBv�t�Y2��(=b
���@(,p�q{�R:)���B��d���&��5��O���5a�ⳣ�W������������wX�3�1p���(!FGU3�2�<A2���(���A�9^�I���hm�0�}Ȣzi��#=ҍ)�E�[gո���s��p���V*�N�0q�\qm���"�'!�.!��v��+r�t�0��AU&c%�D�Υ��Iڋ��.�Cn,[�o��58��H[C~��?k���Ŧ-]X�z�� F�24���ܞ)Jψk~8bå��f�[�+���K�A$�����^�^�|��e#t���B��GCC�,�*�Q�f��,�N��N��Ȉ�f�bI͋�n�Qy]s��ƻ7�k�w�ajn���x�E��8�B7*�U���t�C����A�����U������s�7�z|A�<Nf�.ع�'z����앣���#ϭ>u��-����s<��Չͯn����>rF�ށ{���פ��P2&>Za����U��(��qq�O����r�c`��`���G�XZ�FM��I�!=oS)A$Q��f�	�%ˇZ�$����ז����M;0+�Ф�v�U���dN8i	�}�8v�q�<�Q�=�6l�O��&A>x���j������3��;���7�"O�zq��&B<��=R�'�dX�P��ȅb��~r���w�!m1#���[�yQ ��%ԣ��]�R� ]	5�qX�+U�6C�J�:�.�LLC؇mk_F5?���<���%X��h=m2�
��̌�����{�=0�����_��t�B,�|-E1�A��Π������t���2���X�j-6�݊����o9	?��[��M�ǶMk��8Az��C���_��W0m�9����n�g4�{�U�t<�_��«1�&lM��\��x#���W�P�0֛��ic�����/��7�p�/������UI�I�	V�&?n�DC�Q�L��&��J��K���o�޽��M;��]���i/��S)���UJ�����G?{cG2U�S2��}�t�چ3���u /����Hʘ���Vâ
T�V#ne���$�B!���(����	����ΐ�� 7o
Q�>��9�ɱ���W\�]���`�0���k��0wϳ�r�`w_O����+��k�M�����$��B:Vm�GQLs�V�����"��t!SF4'� �o��A|K{�|��M�0�p4.�F&%"��o c��	ZF��f4O�c�����"#f������%�s�n]W8$����(�GnB�E��O��eX�e�^p� f%��ݯ|'.m�YV�i<�BdLv�.c{W/v�u�����7m@�K ފ�IH����Y�`��`�&�ϋ�QF�uȯ玄��������{��ҙ����e�g�z<y��xiJ��B�w��d�C`�X�u�	�����8���tApԄ�dӬV���oƶ_�C��1wt���1c2ޭ�e��1��CmG�p�K�:l�^F]7A꼼�d�����'�TK�h�TY:0�3��o���D8��\�R�	ޡ�+�?S,�FS���H2L+H���p��A,#��G�\A�&��V�b�(icN�r��;ױ��&����EV�d7��gv�5��4g).o�lС&K� ���<pL�U��M-bc���h��W�g���}z��U��?���_J�&���2�>`���[n��z�WN;�4�L�#l�1�u�w#1aF�Op��o����� `�<��j��H�HD�F`�I`#^zq-�:c9�]�?��>� �������?�$��f��̙5[b,;���&���WŨZ��J?�.��VK������^���.."y,�gx����-?�/�Z<h�<��y1r�"F��?�2=K076���p;���x��%!CC�3���k���������C�k9"�8\4>���2|�~����uQ�l~�N<�1{�)�=����R�W[����&?�:�Z��CL��	#տ��a�������>��d	]�q��g�I	=��=�v$��95��%��t�^��3T���6+v���ޅ��R�ʨpRY���aZ�{����de�,�:Vҭ.u<�4�K+�;!�K��I�&K�*��*� �S���/��>&.2t<6�+�(�����YA*�b3B>=� �����a�bCf6k���Fxied�TE%�i�6%�ʂN.��<����\�gJ(~�$������{�%� �����0ݶ���剧1w�b��;��+�c­E��!lLbʒ�afKHBI���"�.��!BQܓ����R4�N��rrm֮مshµ���<=.tn?�$�s�#���T����.� o{��ҩp$]Y�p�C��T�*�ŵ5+p)D>�I$�%û}4�(��_����X��UzD�1����Ch�'o.UF�{��#�t��U�Ӳ�B�E	%�#��ㅻR"7��yi=��ND��+����)Y�����u���G,r��iz�k��o��C<��j�&��,���X&�����n54�vЙ��ɼ��]}L�~?F���Pt���f�rH�F���>��澵d6��>�>�;v��vm,-ɰ�����1��q9MF�9Z�HN���%�a��eM�LlTkRq���pg6��!��G�D�K�i劺���hlE�{�d�<4���	=T4��lI䚶b�BG��n��[���9Ž�1����!�~I4��\��LR����1-k����ӢH�ĝ~����"�z�RLQ�rk�I SQ�9}�z���a���o�{�E$"!A=d ^Y��9eF�q�oC��5揼�b-��]�d,�dآR��K&��պ�5;����&�W2L�b�6�ٲ��'����y�1�6�M�1�ؓ�/��=�'L@�Ν�{�|9}$�ڙC�h	�gNB�ꔴ��[��{��4`��
m�M&b����7����E,ބY�N$�C�
݇L.�
]��Pa.EH��T�Xr�OƤLnM�]N�%�O��=@ϣ�K#5ԏ���0��e,<�L���OO�«�~�fN��O�,�zs�<�tva����ڧ΅�a� -l��)QPn�!�T�$�5Uk��C�j������/b8���,����e��;���z!���;��4���M���}gc�ϕ�����>y;�L���yfo	Y�K��i�a�x�UejH���.�P�y ��$�a��@�j�l��ݟ��:�*
�:3��i�ɬj5��&:/,�ǫ9�=��y%��{122/���A�P��á2L�?lj�V?e�+�U@�W��d��D�L��W;;QJnG��G!�ͨf��?K�%t�a���*�Z�"�Ҋ������a�(�"F���9h)��_�G躘���6m6B���{�࿿��)����D3����H��'̘A�N+
Y�XE�0,|>?g�	Ug �l��Wb>�"��;�K�qqt4���	���F�&�KOD����Ǜ�ȑ�.��yWp�>�E�����Z'��|dp���#7��}�	Y�����ez1ԝ�Q��c`�@$6�MCOo��wѳZ'��|�@��G�9�p��:�;�"�YB��Ù4�_	�D��}�ܖ���`
8,f��Q�?�v(y�C����
���������Z9C����|�
]S��}Xy�����f�(���BO����f� ê��S�*�a�d�.yE��
�ְ�5!$9����Z�i����f�2+�K(�+���˪�T2�Z�N��B�� ���ZeE���M�XYDK���2 �,���yt���ukXOU�����'�/$��*�rY�&�������M.�RY+�E²J:�~Di�v�5�Қ�B�w���3��^g�����
!��G�U��p��ţaL>�t	5l�&�����p#}�D�F�P���j�a�t��is�-��F�ý�4�b1euKhIM>���Z���vlށ�r��s�6�o*�ɂ�V���t�|�84�vVӫ
�5����+R"1�׃<���PT�IKk��"� R9I��Z&��r�"�5�3t� 1�X���4���s�A���TȽfd'=���U��2�5������Ú��>��@歞I˨ܨ�zKuš�{dy(dLh�h�5"��e�.(�&�)̃����n*mW`����\�����_^�C�gXH��{��w���MU� �M��djȭ�uz�f��X�}`��Њ����v�C�7�����@X6g?*R��2#�9v�����Z1���n����@\%Zh_>�^v]�L�co�\�Y�ЊO�.�&c�1BE2��/vq؈鴚�	q���eF�:��~_P��z��2i_Ä�-�"��݋87MόHCv���`w'��F1�摆�і6d�9TL	X
%�r*r_�O�Vt���	��k2��
�drE2^4�}�92�%Z����$C� �����h�@�M�RA��y.EƤ���(ݏ�Rh"D�g�?B�H�h(N�ˢ�L$�C�~
,E0�%U�UA�&8B(�cf�^|g|�n��oM���
9kJ�J�e���0�;�g���޵S�Z������x�.����G4([򆦽��'oR��U�?O4����Q$�ݱ]��"٨B-]I%Ȫ�P6�F"�.�wr��Q��PƉ��Y���G��IJ�˴�'��arq�	F �r�@+�^M'`p�.��Σ���Dt���NY�˼���&��dt<naɥ�n��p�Fa�D��&�0Bd(��n�*����lm1�c�kJ��$Z����B��rA�j�jdT�ڳ�ZT�)B&��8���C\8N�29̚>i?!��.Ljo�ը W��)����UޣZy�̐
46
?�LnO*ݩ$'Mۥc��j���{aB=;v�4؃ }���~Z4�/��o`��Qu��4�&�ʢ��g����UV#W�e��k/g(]�a���2B�J��
��!E�R����� ǚ^�Xg��䮵�&�-��~ѽ'$�k�{ȨW#t�U�.}�_���cV�h���Gׯ��#��6P��B�c0:䶴�`(��y�G���.*��0��Ӊ<ok:�"m�K�՛BW{���i��aZÔ���V�y`�=އ��ִ�7���C� [欁��H�༎��M�"���ZA��p,dYdpA+(�����$�
�� +�s]#+2',����k���\�'��r��8R��i����d0�p��r�L���"���؂��C��'	�o޽^2P��>d5r�b�ҳ�D�`IcU6r��.�8�A��Ap�ǫ��N��2d�dH�r-� J���j�fN��0O��sfbæ���7���(���D��U���u��k�ɨ\ ��5�-�e�&q__7���E�uD>4��d'�K�X`� ��N����+����Q��'w% �Ƹ�B�?��O<E�'���1i�$r[	�U2�_�j%��B��T��ہbr��Jl-�I&1�І�3�x���Oρ�9�S����/Y�����^���Ƨl��1Y�� 6>�c���?dp� খQr(5j^��P���q��Ñ[<�1u^��C݅�f�;��Q�	���ap�,�Q���9��J��X ��:H��&�X��u���xj��\���V9������?�U��A��4aT|�2!��R�'#�D�"\V�EB49�7wg�'��?���9��n�R���';O:�NW��� "�ߍ�hk�c��V��Ed�#X��E1P�q��`��%ˎE�!�ph�L�͝�u!��]	Z�y�t���
"7+�چ���{�"�kJ�{�c������#�E��=ݻ#�ؽ%!~3�T�2k.��6-�Q����P��=;^E�i�&4�j^	DN��RS�,� ոo��0!B�����tO�������^.͜!B}S�kr#�tK5�!�'�|2��𨰜Y֒����
F���P\17՘�\XB[fi-~SĖZ=���+��T��TXG��B3��=Hq31Bp���1q�)2�Ө���J�@��u�����H���d�Tp��CF��(B���H�cT��N���~�P���"��N�M��kV���bk�X�Fo�].S��/�
��ͥ-��2캭��e�}tC��+��\SR��+��1GӴ*�!c���ps���w��ф��Ɏ��
I(���\��ȩ�
�T��Rȃ���#�S�B�ko���P4��ӏ?,}g.�8z�<�Q���׮�]w�%}{�y���1�VP/�n�I�r���ii(�q���o�]..��+On�VFT� �,�~<��3�1���'q�qK麼b��m܆���c�Ο��u�;ߍ9��~�t�#���uH��Qa]�Vf)�5~2�&���N�*y2&&�>�x��h��g��9��׾�&uH6����]�����?�N;�B�=dK�:�ENg�Qa�[.#� .�l�Ќ*��L�J',��+��>OHQM�ch�frI7�S����K�G?�L������G�ގ�&�  ,�IDAT�{���{	��è�U%c���Gb|�V�䣝��Lr���S�)�;#2~�.�_ȸ����G�"�b�u5=�i�r*W���j�0,ڑ����'vTjF���EF�hV���(�2K��͌ĻQ�ş�>(�}�5���HDj����� ����I�[z��d�Y4q8{�X*CP��Jр����}4��n��5�x��\�^�%a���v���n��8�Q%�����	q�>k�p��Va�҅���(�-Bӯ*9{��x�r���7�oyo��LmoA�H�v�B�1BnV�����0���@�Jf�@��A+��O�1�cV{�ӽ�����ޫ.'Wg
J��;I$$��p�B��ŋ��/������ko�h:�$�!Z���HI;N]���X�҃���m� z��Nĺ�/b�9��?'��� �ë!8k�4:����{��/~���g����alٱ	WT�U鞅��t2 ��t�iR��>�Q�*#��$1s:�@���l\������x�E硱�����h"����`����W����K�����(����):��?�}�Ȉb�>; ��)<`�E*�W�������a��k��]~��Z11��¼G�s`��Th�3��e6����m��E~bc"h�E4�ڃ�!�D�/W�^�abL�f,�l�^�ñ� ��1���|�1C.��"!+'���K�!&WeG3��i���H�jl�Z�C��W0:8$������ %��LWznhU-��D��L#��W̟7�&�g�E��Y0��Y�s��ŬSp�?õW����78�?ލxԇ��=�43!�nZY��L@�� �Pt��D�:-MQ�Bvo�����ߏ��fr��:UK	�xIhlj�UW_�����O=�O>�\�tm�E��]���͙�����u,�u�&T6c�D�y��G�p�w��H4���>;��_�^^w�Uرk|�	�������~�*r1G��6�X!<]�?N_@X��b� ��Dv���,��2>pͻp�՗�A�h�B�s����YAL�h�o���[�MM�M#��)0\��X��d�hV�G;2%<o�19ֲܽ���mv���,�J�;����,i�Պ��3j�9 i�R��c�����1�u�S�	n3[��|f��j}F�g� ^�,@U�֢k��C��3��N.O��P<nh?�����*��d%��#�H�>��{B�X� ���X�KpK��RWlKn����rgV`bG��ǯ'c�J�)<tY��9���ؠt��/}�s���@�#b��0�=���,�+�Q5*�1���s�kt���k�zl&w�܌��FT�#zp�}ֿp{U����7܀K.��n܀93f��W�`td��)sȓ����:؀q���p/*#=HL����nl���~�O�1��ܾ�h�JeKB��-�
�������� � ��Ư~��"2#��<s!tB�\ǣӳ0K�4VH�cC|�Kf��1�;���� _�V\x�[�k��˥^�X᫔~����D8��p��b�������/l�-L���&��3�r�p�J��f��uSh��'��ic(*-nzݞ\�zS���T�բ!���_R_�hS��VQ�1?P�6k�FR����b�s��6"����G�N1<���לѱ��y<��s/$�(2�ڱ-�:�{���OF���j&ȧ\�/�$H]�����@+�b��p�-7c���ʬHVC	S�R�hTˊ�OFn!���+n����캏�я~�g���*\*�`5ݚP�ܲ�F����IXBn�C�܉����s�\)p��r��"�o^�]˂1y��k�y}�Ə~�3�y�[��S/c�ࠔR��T����t����E!���Y��ɏ^O?��%K���t��[�pobP��v��oQ[[�����߸	W_��\�*��{�J�E�9EFU:�tr3��&�3��'t�Y���Y\{�yhii@1���c=��� X-�6�
ޫ�%��/�m�����	�1X��AF2/\"���5�8^'�1�|�����H��-�0t6����_o0U�x�\TO)���zGt�.=�vD���,�f�,(�b� V�3T����DQT�X�-
����L�D}��ڰ�'EtS�E��e�96��1$s��Kh��b��r}��ه�knB�&^��K��i�rV�[q0G��;��e4���x�XS�A8�C�2m��ܸ��YфK�I��X�7+-]�/�S�/G+�^�p�bpƂ"٠:�&a��*r�qtܲ�x�Eg�?��9�E�Q+-����.���}��\�֖��W������{'��<���4!��0ls\�lpc07*Y��9�-����6g�}Ml���}.>9�r��t���F��n,?�8L현w��l�rۯ�~π����"�6,����,�ғ�����]�܉��&,[�Hz{��V���.%�p�o��&���o;�<|��C��JeJX�"�㲢�:M2(������i�ш�@FM���i��Ra���Y��p�Jn�w�߈7��B'c����z5-�%w'�v��v�6��2+R�c���H0j�1,���Z�7c�c,^Ro(ff�����(1�bҜQ�cI|��&3�Z��1��{��G� ��. ��F��x{� ���vˠ�e,V%ůMW�j�AF�>3���];���W�euAܼ�O��&���ED^뢕�!�!���<������s����t�Kt\�x��#�t�R)�]�زy�̞!�S�Y$��jFF7��R��T�st+9��H�~�#��x�v��\���aJ�Kƨ���lJZ\lټk׬��͛�4z�T3�P�t�W��U��l���E[ �+(�&���UP�a��:�V�4�0g���-ւ�h3�,fO�M�P���Il*�U�l��Z27�Թ�^L�8�#�� �璬�aq�a���f�,C��E��c���^����k���kǭ���O��ԓ��&#����r8F	�v�%]Z,\ǓDS�C��h���4k�Q�ֈP����1(g��V����5�e�Y�πV��H�MUYy����Lu��(�LeD�X34�z;�"؜=���̑ad�U�n�%��/��Ti���9�2Y|�a�h)$bB���8x�a�P�#�U)����|�AZ��X��;vw�f�"�̣ '��	��L&�F��A?��
�tk��y��1g�'�D�����U�MF�'����?��47��"��� ��nf��R-ҋd�ax�at��B�a���ظa-��t��n���w9{ �<lq��R����c�b4���5}d|L��:7'=��	�t��L^��n݋�;����׵���&��h%a�1��nV�� 4�utO{ɠ�
���w!�/��k�J�����{�WW��mB"���!.��LDVA����9
����G7�
�&�2LQ�������Kz�Z������1Aϙ��󺫫�-�������u��d`�`A�voI�CU����BxW��^!�X�_*EļG�f�s��Z�"-	�R�I9��y%'���*P2|��G���VT�{�i�j"��pW�F��P���Qj765��8�rQQ$Z�L��H|�l��Fы<�顽8�ol�P;��~�ǬO'b��rR�CK�rs�T�S*	�.�Ɂ�x��4��������ۦ=�kᨳ�	�:���?������h�B�M蜮��$ąг�9�����ȷ]�ux�gt�ٗ��� �{#�SHT�h��x~5\u�RI�z���g9�"%Ӹ�q^��C�
��f@���7�W��q�Ip�u7� jL��fhmo��Y�c�	�u y ��V������_��~�ظ�Y����Q���1M�Q6?�~��f��R��e߹��.���Kax܃d�M�<.z�2�4`rQ��ZO���b��;�aǖ���o_�_s%��eт�0���3.7oN��UO�%�+.��G,|,[��NlgS��d#1�����ȉC5��Ty�<��hĻҜ_�!�xh�O�5��j�]�#���Mʣ��Rv�@��i�t���v)$P}U[>v2��}�ю�[w����\6�WZ����[�G�F%����yU)��h�RUJHRR],5=*Fl�F����0�3��JB]���1a�ƪ�>Z!	����x4��m���X4;�(��I���S���������b�Z�gs���Ȗ�~�l�K��xr%\s����]�D@�-P�Z�5D���q.���U?����G-�5�<n��t�pv�(D�2�<��%(tt�����ǟ����Jm�p�ŗ��_|1~g��y���	*����7��M8��|k,�y��Tk�ݻ���W�RTO�5%J�o�Ϯ]�Ё��<};���_�N?Ł�THܩ,�0!�:;�|���d���^ϭ����q /P(r��	C�� ͆ pj`��x�}����n��.���? �!0�Zbf�j����\�ëQ3�ള�7�g^xa;��MP"G3���~X1�o�2H[�8��E�D6��yW��Hv�c�)!/g9��ߌ9���ϳ����u&
�eJr��	�2�ȱ�~$�����WJ��)��n�w��?<���ϟ�������^�(��w�}_����Z�Sl����Hs&��
��>�$R|;a�8s4�؝� ͤE�y湩�C��x�[?~�v�h��F�K�ΔN��S!TigrT�#������ ��lr��t�f�Wh���P���M0o�>�`�"X����|��E�"��V͕\�� ��K��l��KN�ǟ~FKU�<$���4 ��w�J��m'��
�P���"tw·�)���Ї/:
�<kl6%�c�p�����+�w�����Aȷ L `Ren	5O�'G��k4=�4*t̅�k��/{>x���w-�
��= ��.h*�@:���c[�^��~�{�^8����^�6�*�@��Z��F�8w��~K.k)�q1��e�LBM����p��@siN~�	0gN7'j��I[�ÕW~�s���/\Ś��k��w�&'�j�\^�1��_,�I?��?��d��<0�� �|��DFҥs�M��Q�>)l��j`S.��%�c���u�Ǳ�]��� ��cZ�ysf��������~�����ً�_9W���� �f�_9���_��S��Vf����E��y�rY�;C&C�j&�!Q�iG�iVM��X����u��`Ğ�H�����^�H�x]�K��dlH-n���P����E��&H����y��6M99)�B�n@�G��ekyj5,<�Mp�����r�x�I8��O����h]��
�[�	n��6����q'��X�v}+�δ�F��u�r&S�����$�^u�hB�r����Qطs,>�L��}��e��>��sa����%�����V>�N=�l���`��Cw�45�͡J5T�\N��C���)���T�<﵇�%_�V=}�n�.�؇N��s����X�d	�����Վ�:˗/��������"˰q�v�(�J7�T�r[���L�QC�xB��4��aV�A0����3P+�~{�������=�T֊aŊ��ƛaͩO~�"H5wB��m���ҭ������`:�h���^��,o�뎌���:�39�`Fd�Nl����kbM��H��TO�0�Sh�P��7�*�`y�t��lY�5Ty��c���sz�^r����B㒓滿}���m��}8;H��Q�=޽��*�PR��@=7"�v���bʈ~k��"(Ԑ��Q �<�K�i�mF�)YUwN3����·2�S�d����a���nj�[7#0���'��a΃ŧ} zV<?��mp9�6�vp�)��0�o=�4(;9�E�~� P�a>��p��uO�cX�g(0Ր��=��9зi=�Z�Ao̝���è	����!�M��8�����(Z�a��ax��?�6��01�&��۠X������q\ӜPw���>s�>4]~v�Q�p��;�&>Ԥ�[z��kYC�V�|\��H8���Q��}�;XBM*��ZJ*�h&����L����8�6�8^Eͩv�B5�{|�i��[�;V<�����B���3�ܼ��w�ʞ5PB�in��
 ��2.�����B+��%����e���Y����36�	ևg���_E��w��ףl:#�qN�Նky-M9��
�m�ѱ�M�R��;/���;�~�f�+�^_X����/[u�}zZ���h��G��E\��U���{���$�Y�U�����ƇeL��2�h3e1��9�`i���I�^�H�(}ނ�L��]@��
�֌�}�P��$�m�m��͈v4qVod6�B�\8��p�lWWj�jO�o�1��/�-C��,���P �V�%�����"q�$��w�N���q�pA5�D3v��Q;�m��ܩ`�A9h��r���m���BK�\��k��ȴB����<��\7K��=r쥹S��s�k_�тG�e�w!�6����9�jv�ɥ�wd.jG�%/i("�Up����ՉXҊ�6� IQ�0t81�o�=n	���x�7S���$4�;��S��3�`֬�𾷝 9|�U��[�o�aԂ�=�,�n��W�M�7J�!�͎� �Ze7:Mm��f��v���q�P���^�15�k܉�f<�9{S��r���ˬv��ו����E⇪z8��uw6sAq����ݿ�э?�o?T�_��k�B�_�y���yr�k7z��j)tH���ȓ�}/���g�$I�D4Q0�7 �+;U۰!��W�X U����ӇM�y���;1�DqF�M�#�W��D�#�4b��ߛ:_��:a���0���F�՜���I��3�y���Ќ�a��M�y�N������J�P���q�0�Z��rV�(g�T�L{7�*E�>Џ���xZi��h��z7p'�j��4���w��YUN��@�P�)V���痌��9%"�4�+ʥ"�h��QU�f�h:tZq���n��Y�iEm��N�}��w�<m�����	u�zqXߴ��&R�Q�[���E.ی@��H�
eԄ�.j-�ŕۉ�R�$k�%���2�Z
%;D��s����J�{J�l�����"��{�:������QxOh@d�q����ʘ��߬�n���gꦺ��+V�n��_e2~_���hj��Φ�z���K?���_)��ث�B���>��w.����������rX~c"�� �Pu�6NGv��Yj=BT�:1H,i����-�N�4�BM����lK*=�[^%�sW���k�|�ٟ������X�>�pP���/��
}�JՃ�}����jpc����Or(��
����C�w�D�"c������I�R`r�ؙG�%���?����2�Ȑ�5�`��0��i�u�`�6\���x�ѐ���-��ܞ'�E"��<nYqD+�(
��P�^SS�J%6�"4/��p$a����[�R�os?��1on���z,�<�|�A�l��s���~J�ݸ�k���h(��(ӕ^#3���Rԟ�RF�7��(��c�*81�y��Ԫ����$�Kh�Ն��MH�꣪T�(y?b�JMT���,��&v;�h>	�X٪�gYɲ��&wf��p�D-��5y�z�l������8&I�#��{\�9��ͫ�|���.9a�9�9���^�v��kYu��K�[���H��yn�%�zx�g�`�&�j�[�(�����f�.4kV�f�5=�}(1��ty���?v��
���&�di�la���g�J�X
|N�6������3@���X����N��$�h� O��N��"�WkPN���Yv�j'Ŷ�"Z�@�܄���)�R=H؈N�
��-�ʸ��Mͼ�j��7��nL ��_& gs1ץ%*E ��6;��.WyS�B�*�ߝ"���$�h�eV��Me�f͝�uM�
��?^�L"�ϗ�6j�B�NM&�$ �����Y"�(��$��P+������W�(���!�+oʹ �𭯤�¯��:�pR�8�}!P�360�5Fd����
�?�[���{��G�u�k}4�OD�)2'>:erc��-�T=p`�(^7�y�(+�"\Ԓ��r
�,j`E��g��7=��q�p�e|�y�ǫ(4>�����?�s��w�_+�����3�͛{Z)q��876�3$�j5.�)l�����É�DQ A5�m#C�g��>�4x�B�w����1�8"��&T�$���}��D�8:eWt��yL=snihO�������;�Jҫ��t�MD���k��*Y�1�U���xG4��rp�Š��@���Z^������ (\Yd��?�Rvs3ĵJ�ȍ�J���q`�'��]��ĥ�%DS�Eө����()�Y�����A����%�y2+��8S5�L}��{�b��MUs�E�V�>Ȁb"��G���o��1c�h�n�A�2ZG��8i#���8[�GD[:#Qӎ*�#��!�5J%_��k�ԡ���/OKd���B������I�jN^ۧ�0Zٹ����j��S�~ϵ_��h΋�WPh|���o��mw����7<��Y]�Z4⥺&��H͘qgbӇ��6v%��aOK�SG�E>!�LP�=��
D���:�V9��P4j���B�F�"I\�������]g�)FK�J8T��M6�=9>rʙ��Q��7�eh���$W���D������.8�zH6�6im�/5���p�8�iG��� 蠊h�S	1Rn�~o͋�ږV<��LZ����Pxrz���MG��n����o��k��$�=�>�,^���&�����{(��$�I��'��.�7:{dH�(�ϣVfC1sIA%;M#at���y�V�n%Rx��4���������9�k�G6A���"$�>�g"�&u>5��k�K��mͥ�2��#����O����/�tg7ƫ
(4NӜm��W�����O>��D�~�_����{�?�s1K�p�:(�w܅��V��W��(��c�t��3�{���v���R�,X��[J�jek3���K����3��j('��P���BpD���0�	�*��^L�!���.n"���IL|�X�Z����-�G�6zf�M;�i��pE:v�2M�A0vL	�pض&ܐ�I �4vͮB�x�*k|�R��
�]�r٧Cf�����3>'%mT�g��=�i���07U3�64��Ik1sy����<���FF"[h�5֐t,r��|#+ �cф��<.�Pdؚ�F.Is�ʋY�fG1K�
�O�ԠY�5��H�?�;�� �f2mBc�7������g�w�;`�WPh�T��7�ӵ=��Om�A���l:1�[���Ԥ���)��I��*gX7Yl3����}(vB��fA���	>�+���TV(�aG�T-�X�c�
C$���Miu0U;�uj"�'"A�MHry+2�	b4��S���H�p���`����� lն��T �(ٮ,��P��k'`��NQe.��;J���6&sGg���k�C�/?��MI�3\�95���	�J�����I#�E�vC�)q��Z ���1Ϛ�-�y����QLpm���� ����lH0���r5�c4
� �!c%�e���Tc71��y�"�`LS���s������cJr]�OFL�n��� �/M�J%�t�����N�v���Ae|s:(���O�{�'����� 
��nE*֊�^y����[6�{�P+�G�l���D[&��9�t�ٍ���q�l��W �//\���hs�h���&��M���FA��
��H�ٟ��NPh_��7*Sf��d*�4�_����$�n-_����x7��0��`SRᩤà�EQ���L���p�ජ��<��U��K�q��5%�)��T������!���i�!�%�rࠕ�1��3�/a7�,%���B���  �\�q2-�蹻l�������ݨ[�gx��(�RM���k-�\��a�I�����^p9,Nnm�C�D_Mk&A
��j�WY�OҐ(ľ����Ӱ���վ,$�����{���M4.Is��~�⦅�P�#~چ��$�������L���b����ĩ��Ϛ=ʘ�����ˤ�`��%���{�G����O���'������W}��?�r4�P�X˔�&
���t���� h�+��\�Zi+���2���@	%|����@�[�p�Jr�\{�H�Nrn�*J�eBe*�P��۴f�Wh5��d������!Uܚ��Y�L�˙�r���h	�A��/~�DJUd4v�c���e ��x��h������JE�|�(�!��#HěА���*�
\�T�[d��45č?$L��<�(�B�"�� �j�)b:y3|?��Qt�@����Q�`穸P�.��,?���Z�����#'�+�u���ME.Q��P�B��$�4w�<=�i��3��j� I�U+�;�8�@R����O[?�	�F�Uxz������3�mfy��p s����F�'eGI33���R�_��zZ3SxhP|z��������n*�³�&�q�	C��"�lv���F|}!�$�u�,P���8�6�bU�Ҿ�U����x��ڒ������>~��?�����Ph�s��/=I5���(w4D�l��;�?��%q��L
�o�!ofjB���PN%"�'����f\�Eǘ��s���r�;U\5�R����ڟ!���h���R%WOqȸd3�$.ry=0�P��ڋ|�&�=�3��a��Gɡ�8�j_�M�?u�21B9�
�7�?�壼�w�փ�R�Q��r�p���?41���{���rj���{j5\��#�ϓϗ�P�J��c&��y�Z���&'p�A<������j)�4�r|�CWӹ�T�5=����A�A`��X��	�;�䡊��J�H���	_�J�å�|�$.[��/z&A���q[%"B��B�K�[u2�`(���������F�wrN��ND��sg�(:(TI�z�o�d����Bp��!/���$�^�>Z$a�J3xcA�5u�o�g0Q�q��#�:���k���S�$�r�Mps
p�a���e&u!?�M&F�`d��+�J�&����u�C ʮ�����qf̌��ͪ�cw��|awA��k�{k���̘�߆R/W�����+��+3�23f���ccPf�̘{l� �̘3c��?R�W/�}    IEND�B`�PK   �KX�����"  �"  /   images/a8d700fc-8f9c-456f-9f71-f71b03bdd111.png�"݉PNG

   IHDR   d   7   ���   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  "pIDATx���y��U��w�{kJ���2UBI !�DA"�Jd��->�x*v�zK]�G���(�����2=��L �		�TU�JU���y�o��w�͗�M���֩���θ��9_L��+5�W��5G4�(����e֬Y���&���RZZj�g̘a����e���2g��:u�����Hy�AY�`�L�8�ʎ;&��s�9GƎ+�x\>l�K�,���+������r��Jn^�h����K�.���l-���2�����;O23�dpp�����om��ӵlP���csg�h4j�w�ޭm2m.�HTzz��^nn�,\�P�G�����7N�ϟo}���[�)S�HQQ�����ظ�=��q�����_i�s�|[��ͺJ�� �	F�1a�1c�Xx�XXɬ�l�S�Z=RQ��Sh�Y0i޼y2~�x�q�+�a,�z�@���@�!MK"��ŋ+���l(�����ٸCq��r��u>�A�H�,[���g�V/-.˗/���?''����͑��?_222$;{��5//W.����-�YY�V�H��u��6��q���0�4wh^�ȟ�|S,� 2k�]��!�h��Ha�X���%S
��92a���˼	ݒ�5$�+�����d��.�Ȯ#AY��-��)]})�ɲ2ڮ��!�m19X�i���ʧ���PC�m�P�e)%ʥ�ڥ�:Kꆲ�3 �guȎC��8r��䳋:ek�rNN�jж�������dDe�y�,�
D�d��9]��4G;V�� �O���7��w�ebn�O��AQ6��Wf��-�y�_(=��_5�i^��7���� �n��͚�I<7�-��5/	) ��7*������D�o0�T��֮���2�5uƴ^@�^������ֵ���j���?bm�,�IMkz�����ֲ�����BY��,�+�g�2AE�����o "5:n��As�m�%J�2��О.i^���K�!�5wiި�� d��r�[���G����$��:�|i�[�Uy^.ӦM��h����`��;Xnb��=���w���#2{�,9�:���z����c2w�\�l�1���*55��6�8ioo���F����ri--&����V˴^CC��1�YiM�Dӆ���Z9k@�2SJj2$�KU�QC�4Յ�E�ޑ#�U�d��)S���E����$Bt�$�W�ieD��r�.S��7��G#c��[��1�d����	F8�yn,�f�k���>��!uuu���ۍu#
��"E�¦(M�켌z�nkkS�5����ߔ�d�e�_6���@�2�eMM���!�������̥������˨G�C�����{ƟX]ce�G?<#��GOOOr<tW���ѣ&j}��-�&� #�7J�%�5Y����VF�CHk֬�ɓ'KGG����UV�Ze� Q ```@e|�TWW�$���.��@HXO^x�!�	�J�-2�����I�&Y�|�)}�0.ϔ1(�� ���\������A" ���!��7s����&�qS�  �{�����ߖ�+W�a\<�����e�]fk���\7j~D����I�OwK`�"��k�O	̍*!> �۹s�Mj0,�Hʜ
��ar��Ƃ $�c2��ȑ#f��t��2�ji�����Y�����7�'��(q�5sչ���ː��/c�y��qP���q*��Oo��:���3S1�ܦM�nEEE���jY�b����R�|�4�^s��F��!P�W�u:���L��
۷o��3eήd8��x�y��7�>�#C5P�@��:~�������p�|�W�Y+�Xc ,F���Ha�!��ӧ�5��HΘ,��Ҏ�"J }:^�X{z��6����+=�u�$ѥ����1ي �'��I��ի�c�b��Ա�y��Ek�_�D����3f���
���?6?�#e�	��C�i�o���}��GM����ʰ>J���/���۸��;�AE�����7��"9����p�O�[�t�\��+�y�����wݩH��}�{�$�.bq ���A~�ؘ������Ųt�4y�߶�u�_&ͪI�n���޸B^���5C}����?m��CG��l_������4�c�{���d���!�Z>K��@��v����Ȗm�r�Wj��2sz��9Y���۴ϕ�g����������{[+����Lfj�Jԉ���?6j$�%�s�=&b ����M,̜9S~������G��&s��G�'D��wݭm��&�QJ�ʯ�_v��u"5�Tt��%tx�������,�}�.,6N����Xd��=*��&���ϕ���R~4OV_|��4E��[6WJFd��OwTT���k��õJ�铤���RV���Jsg@�\8K�VFd����{��4��sR��}Α���[���5Wɡ}��}KYe��_����,+�!b�u��OJ�=v�%��ۏ�裏Ј�;�cJ�ӟ��a��_V�8 /���YF���Ɔz�U t�	n�K�n8�O�K��3S��ʄ��f���~e����}�����O��.��⠽�û����uލ�=���$��=	`"*r�z �y!=H�"��$�cP�"=���Fl��,Dy"���S�����-]�0�"LsLe�Ͽ�zx���G���:a���z	�7|\��immI*g�h�o��v.&�/��GB� �caڟ��C�yb{����3k�-��w�}��)���@�m�f��e �o|�V��q@O���$bS�'��S�k<��To�����C��M
�瞓/}�Kf����@☄^�nD�y���Q=��w1�aEbQ�j3��wl#���N3Y�.���@F����{fـ0��[o���r�k&e�@��{v�R|4)6|�,��yHߵh6��ON���|��&"`�c���φ����7�h����ȸ�~�/��3�! ��'HÄf.�f>�"R"C�B�;v���b���$wn�'i��L楗^2�v�ڵ��� �I���!��#����Sp�#�����r��9�%��O�ؒb�b�*����`����ȑ�!㤫���l~2�""��  Y����(u@\򤓉6'�A_n��;iw*.9U�.�z�	�|�<O�x�(y�q�7ʖ-[N@��Z[Z�M4A���:��T),��|2�7����(0��f������;ԏQ��tu�����7������%Ͼ�S-���7s[�bE@ڎ��!I�S���snIe�p�W�g֍�{6\�8�H��b�' ������N	+'�`ee�Y6tx:�6�������֜�C�u�2$��Y2�S���x������Y1ɻl����͔%�L5����������N����l�}(���l�aY҇��F�wR2�S)1!懄>��C�h��;s$��ݻ��S�?l���g�Z�H}�|[,Y�Rٻ���d�6�ʴ�C*͎��<5i�U��7���y�ޛ�`�&�2��D���@�H��	�aU(n�!�0Q�D\��[��l����w�+W^y���]w�e�qx'��P�٦��xA����ʖw�J���7�"l�|���Y5�ӓ�R�ψʄA����C�y������1\<:W����b�t��[�\����l��C�J���|g<�C-�9�ǽ��+���j�!N"�sVu���Ǩ���=�|O(��UY{�W_s��^u�������;,+�Н��e�ª�ќ3g�\�z�4V&�Iy��/��֓Ň#���y����!��I������APD��r��>����5����o���f`�Hxd�.����c�=&�<�ƫ���@�QW�R�u�� ������G�(�w��Gy��-���o}��ҧ�xB���ԔdKK�E @<2��k�Qjk�l�K�_�{A��X�Es�X�����"X���J��,J�p�ъF�<��~��%A��g,���k��`g#��<g͞=���m.? Jc�@�G-	0ʭ���$�p�"s��0�_� ��hl��Y3gK_o��< ��כܣ�@��nQ�l�Al F���l�ٛ�Қ:�d�x��a�A 2�|
�1X�w$?$�:�ebD�;� -�d�B/�����
"*�S:q�m O�`�'f{�j�q� ����=��s<^��,++I�8�)/�/���V&��cǪl;��K/M�E����6�S4�I&7� /K��l��Om����b�X4 eN��7z�Յ��b��aB��d��1@8�t:��Aux��
s
	d���|�:7���e�$�D����d�V�ѣUI3��VW�Z蜄N*Tj�8X����d��ܴ^������7����[o��a^�r�/_&6�ju�;������3�N�p�U��&�5B0�SI0`�.N|˙� �}�T��$�J����+s&���N�?��(2�Y��e�I"�W���_�w� ۷o�쉾���O����ig�%N��|��f�r���O`7�A[8F֬�cGsR%��C�$c8��C��������Ɔ���$���Mo��"���p���ş��v�|�o8�	����roy�Ώ�U�O�+�/��[p��c�:���t�=�q�ֹ ۴i֗�+_c�u��t=�&��0)��t/��(��S?]����yx���.� r��jY�l������-e�?���vp|���R�|�9���9���w���,��}���[! ?�;�ԁ\)�� yg�|�s��=���w�A�4�L֭��&WVv�8��1*�6�i�k�~J{�{gg�^�[�y��4I���7������:��ks��3��;��9pg�q�<:aTd+¹�x��K��͛7'�x4ł�,���<��}�D��L�l��T��$'�f�d�o�vB9�[�Α���H�����2�x�)�;���'p�w(���c�9�Q"��J=t�h�*F�4�/�d(���r8��d`s?��1 � y��ǒTw�Й&��c�G���N�>������ma���+�P��$Qq�vJ(yp1,
InR;�����c�vGd�Xsd�i�h82h�E� <�n�р=j
`38,Ɯ�����?�`�<|�� ')';C.��Hj��)ڧ�bF���F���a��uE�}���i���T퉠�E2<����pVcS�mK,�ܕ�P����'�|2����;aSz�D�I�&���9Ë&!68���IZ�z�W���k�R���&;'�޸�''�ᦨǲ\�x�NH�|ox�c~ZнW�7my�@��k֬U6�ׅ֞�)�/�~?�����s7�f�IvAzkk�9��p�4_=�u�]$-]�ޛN�ׇa��u1w�+e��.p�CF���ew36j;6H�_����P^8��s(�M*"�L������{v�A�+ s�z���D
[r�v4	J\�r��;�q,Z�0����+7�؉�R�� W8��)�Bq��8��<��.�8^x�tɈ7'KV�?_j�e4����z�'��)w��_������?��IC�"��X'NYpD�#6n��qԁ�	@�N9���Q���S��h#	MS�(5N%uu�I�F?9���5�u�p�D�� ��!� )~P���x�D��� [�.�-o�,8/6
��@wR�?��S�?�)ɞᐃ�w
;��q��h����'���������@� ��������㔢�%��+/�T� 0,�����\;�0<���{2��c1�`��	XZ���hYă��ڜ�FY�>V�,o���'M�'l�~���7���w�5'	������<��AO�cN��ku��w�<qB}��7��htPuG����U)zlR�q�=56wʿ?�S.��̓j9!��9έ�(�a^�Dc Ġ���)���n4J=pF�k�)���ݵk�\q�F�t�����5�\m�.Qx[�l=#�)�Pf͞m~D{{�����x��\���QnzY�1�LN��\�i�X[z��!���ALn�;���� ��p
F'5c ����j�(����Kd����M"䡇2d`��s��eQǘ$�w��i�=��W��&�1
��%8 44DT�u��2��	@���l�u��C�w��a1��@41�v9q��n�l$���W���XuHը8b��2�@�'�Һu��.;rq�%r��!���{F���2}/:g��ٽK�[�%��(CL�TU�*��Y�������"��&I{��ɣ�Wn�Z�C�xh�nG����{�X[��X����ok�-�h_]�6��i1����O�S����p�5:{��g��?��-�@)sWJ:��/���"�1���{���;� i��-v�=��E�{����?�)�o��¡?�@�D��?����K�ͪ�I�wt���XnW1�.1��a�bU1�_��I����nR�q�!fӦM����&ĭXڀ��F�|o��G�\�`!�`�V+{�|b'T�9D��ܹ˨������O�: ]$����Q��7s�-��C� <��g����X��Sb�.��q���+A7����o$�d��#1���o��V�����0�pi�3�''���	����GW	�p�ȯ�s<�& jZ�����͕g�:��񹤧�F�?%B��v,@�'�}h(�Is_�|D�}���ZX��@"J�;(??��=�#����T�`�|��7n�h��������0�&��S�T�2���|��=	 �D�'��]P�AL�Y�s`<8D�!�p�� �."}BC�����{��6��k���g��!?�я��1 ��<|���;����H8�{��N��wؠ ����C�	���loo_�T��t�b@�7ސ@x�!��U�M�v�r PW�(����%�䉿| �a�46u��ͫ�6|"3�Ȣ�)��3[e��n�:<$�^�(��fI��,������_]-7�ܜ-�-xz�����-�o�{���������3�d��VG�to����er��.�Y�Չ�hė���n��6�Ǯ|�~��X�'�0�GM�{':�`g�> �/��5�T����-�
k$ l���u���޶mۓN�By��]��;�j��˃m��m��?����v�0a����N�R���Aff�|�����I�1�m����6$/m|��|����[�hlD�}`����+)���7�R��ȯެ\�f�������]}I1�KB-���C�9�湚�Y�pe��w���I� �.��rS��^{�Ev����N��'f�肛� Āg�t�����17n�`�n��H�\gN��R�!�T�}��_���&ikm��7�r��|RbD�q7�Ζ- CgaX@$lJ���{���믿a��H�K,S7|85ÁA��f ��LD�2��/7
�W�O2q}�w�S��$���<ŷ��~I�fͅ#a.  ��t��������"���I���Y ���=�nx�׌��N �{LZ���C���m|%"8>4(�� �4��-��Q��}��Z��BԀgNUr��q;:��q%��z@
Ҁ�p�K��bg{��PX/D����`�:͉mO�7�e��!�X���apFA<���i�����|�t�Ꙥ�$��&
�6l�`�P���2Bh��X< g�hD%��m0�$��@,�F�S��v?��~B�2 J=?�ȸ����pm���[%�M�Dz&�OK�i�)�!�Q� M��� 0�{Vv�����^�ó�se�v�.#3؛��갽DA4=���������fZ��tE���s����mjb$Q���`���)ត_���Civ�`p��ʘ�#,ħ���Iܔ�b�'M�K;��_����7]���\�!-�
M�ć�-ґ�"P*E��@r�R͗i~-T�u�	!�˦Ș��-c2��`}��� ���.��L+��]j*��R?d���E�T$�`N�1߄�y:����w��<3/N��V������A9gZ�mJ�±�"��i]Rѐ)�pf���Z<�[��f�$E�}K�xj���4D����H�J��dQ��>)��+%U�F ��̊�ɬ��R�e
e9�2�`@ʪ3�:��e�ȸ�9P�mđ@�?h��|#�z���B�@�����%�e��2�d�G�C��=h�
�b���w�xW�e�ǝ-��3h���dN4��Bz�^c����ײ�.��� ^`�O�뗺6��z�(`R��}u��?��`Pv�N���}q�?)�_��)���nv4��U�%����hB��/�ٸ%��\f,.�$^���o������˅�g5�)�� ��H�{;��[%�#���+�C|Hٴ1���Xd��c�x_m �"i�Z�d��Tei��F+�q$7�>-k��my|bQz���ݨ���|s���Ղ�z��/��ޮd�|���̞�;]�\�(+0�tuv$O��QVh�X�x��_�h�-��.I����Ҏ�F����2�^��ʽ�3[�;��Nb�* ʫ[���%���9�DZ�Ȩ��D>�?��M3����/g����PrX;��B^��4r�= KBibY��~V�&|���o"��!\�s�X,�CY�.�@�a�����n�����8��Q�E�B&��_%�9���O-R�a����e ��y��2��_q�Oq� d@����������    IEND�B`�PK   yaX���4�  	�  /   images/be3f368a-d9da-43c0-befe-16a00a90d491.png��cxf��.���6'۶1�m۶mcbMl۶mNt~�}���}���W������ֺ:BANARBD	4��~& ꟶ�?������H�4��������e�E���+��֟a�zS�+Յ�g���M"�@�	�G���:��0�ޯ��8?�P�	8��{��|���b*$�y�0<G�QlG�ϛ�������߫�M/R��ߒlK[�] `��w�]׼n�N�B���R�)�j` *�!j`��0M���0MP:����#u ���(��+��pS �:����o�M�|����_0^� v�taʿߌ����'$�_<&����Ȁ� �`�G�y��?�����nsQ͓Ư��G��͚����������6D����{E��e�&���X4�?¿$�c�ח�G����I�]��{Sza��;�������������7@�/��������n��e%}�8=h���h�o����0h����<t$�R/���|	�ώ�_�x��$��D�H�M˹��KIe� � ��-R�*RwO�K�VS7cV�jV��."�Q�E���H�e��c)jp3�aRFT>�V��3�*��T!������8Q��C�{5B�Y���"���y͇�V3stNt�<���,p)�n�ArdO�DX�
d�ҭO��Ң��[EMV����j��3>{^��΃?`$���/�-Mn@ػo���&�C���[�^�P)�ߡ��p���Ԟx�ط��)f�Ә؅��HоƃP�Ђ����^Q���O�)^$/��R�s|���yw��Vl/�왱܍��|��k�l50~��M���⇮,QF��(R&خ���Ү�ef)��_Sl��Y]G�c�@�.gh	R�<��j��bJ�|x?G��LCM~Sѽ�1��/�L�X
��y53��C$,�������矏َ3�M�khD�M�Uz�ih�����/wv܋�%�|C� /*��v����>�WWW��g"10�v��r�"��g˥˿8/�3p,�{��Ѡ�y+¤bEs|�
0w$�l��W�߳��ƽ;o�=��n���J�7��Úv�Hߞ�C����r'�V�oX��.9*.SVH)J�����������1�G!�ݠ��tG߷<��H�@0tHX�	 �@���&m��#zw�q��UU�孽h�,��U8��YzPe�/�,�PX�+������%\iAֹ�m�NR;��`>�/%5����<��rM�j�6�ne����'w����U�7E����&���Kz=靈�6��V����k� �/���Q�ޢ�#8�2/N��^����k{`�
���[>�c��np`7I����A����7�d�YQ9��{� �t�!:�|��К
�y{�������E�Ǥ�P�L���ƨ��BEQ%��F�9�������ӗw@�-c��gq��),k��,�2i$�󾂯R�����r��@Yk��p4#������;�;-4lD㓅/�46��I@69�����.\�嵪n���<����}�>jh��<�*�t'h���Ѵ���#j!J�)҈�$�R:G�Ou�l	0'�?).�X��
ؠ�ʣ.o�븰۴L����YT�y�y�u����Oފз:�ާ�����X�u!�ﶩ]�������z�:�°Μ& �	"N���H����ۙ!�e�x���<�a�Ե�v DYZI_��_�0��j��|h��z���qQ0�H_h�5�M�`� �^�(�Xߋ����~�NWs3�q��Ջ%�Q)�=
t V���É�h}�v�8Qk� ݳ�����ˍT���(�E��G���@��l^.,�_.r��Y���+�#�cjV%�^C{i��;[� �D�o��/�\��B�%����*p�:;Ӈ�;�L^�<����۱��9St]��39ԓO[7�Y����DZ��a���~�n�=�O�!����*kQ@#ȗ�0��*�ỹ���E��>�U��c����:�#[U��4��,)$k���|L�۩U�	��Ɠ�9$���g�(����{2b��ǔ�ۼz����r2�/�r�rﰽ4�o�r��R�D���(�-\���IWI�DǊ�N����8����W��5�H6�H�&�*0e[_8u&yl�!	z˷h�ca�\���6�K�?�� �K��eLxYxo��c|l�Ȍ��y�qcv���Y[��G�/.Z1(I���۔ܖ.�ހ�iU��+�9�QE�j]/f�3��$@@v�'��`�-`3���'�%�'}��0]+����f�3�:�s�]�Y=�8��_��e$�b��'��2<�����-�~Fh�wٓ蜔>Ͻ*5��M��-X7�)��:�����3���9!j�U������K��nmZY����R�}����i�6�4��VbL��=�Ī�f�y�>u��ܒ+�xgz6X���"�#$u�������:��]^�t?O�����;�4{�����	�	�j�L75����'�!z��E�v����<iB1������G��TB������Z�����ګ"�E;�'��
1�����f�n����sp&`�ő�.��@�7�R��>v6[�[ҋ���dI;<OX�G���bY�V�Qe6���7ъ~b�X�͛���4����S���N�-�����LI��k�|��2{�F��(���4�!5���ڤ�"ME�g�s���Z�.�
�Tٮ|H���Bi��y��d���m����W���NK�;�,��-D�~u�}Du����ʚxY��H���7�#C�+�M肞p�Iv��0\n�Z�������3�K;m�P\���k�U�G�?��G�];H<�/�i乵��e��oiG_^�1`ѱ�R��(��H�_������ڃR�w#%D�SX�ػ?�M��,+gx���j�o[B��K+�x_۞Yx�|�VVHD��!b�_b����w:�^�;���yr�s���k��K��6���s��F�
�1���x|�c=�D0�Nn�`��8�G��w#85�Ж?�б��iq���I��y(��i#��E�6�{�8�?� ��z@'#�v��h������͗������M<�&&I۫�����R�ԩ	:0I�λgʂ��?��0٦Ua��Qg���U)\�� ��mܷmJ�6r��9�����G�'��Iq�	��E6�j�Im�vfew)��	T�N�u���V&�Y�QK�Y\-I�k3�`��D��`�d8N"�*t[�k��C������&)��]8�Ae#��&�Ĉ���pi�lpRU,8���p�&��l�u��.O`y`zj:�g��cVm�NSTu���q���t}}]Sv��"�yCr:8:f�(�4�hy��/�cV���`�V�KV���ͻX)r�> �K)�*˰����p��7uR?��v�\2�����ԷGx��G���7�]19���-˫�[T����Y�Q���g7O��-�.����G��+����
KfC�"�|��Sm�����x|ȽN;J
E-6��&�M�c�F_����޿49L�D��l��B+�٭��Ab���#��ˋ��ãE@c1�+C�O#g�>s��U�@�(�{o@Ԥ*����r���2��)��)��s����L�<L!9i�F �/Qh˞��{�.��gp���B�	ɦ$&�"rm�����{S�N0M��2C�t����w���E��:(�j�h�='=���d���*������.nSV��=ƕɚ�RS)e뤇ń�/�W;j����7j� �::�Ju��B9�\��ٿ���_z ��#W3��󦞑��.��j�����3K�^i���b��� 
ojM��O���*�ʭ|�r|�	>�3	Z~��^Y�����X����w�x��¡���<�/HTRG�V��,�����S�<��P�*��0���(悲�CT���0I1��M��Deq	y��ݮ�r���~!�ضrbY�0$ �P.��fy��udk����VH���P0p�+�<Ğ �&�5@����b	���fLIc��hwdQ��*����\����*2Fnq�|�>����I8z�P���1���Z݉�G�K�Z��Aӻ���hL�Dj�
��Mj���bWQ��Џ!�Fz����j��>l�Q	V��Ͻ!0����o�r�!X��w-w$œ��y�C��q��f�fM����}��gت-��B ��<W�u���C���������'�5̐��u2�#�gD�dr�����u�-,C�D�9��gb/k��AxAЂg�%g�IJ���C����F�$'�L�e�wL1��[��a�q��gʥ�h`��Ql#g�;�Jݑ*�Խ�)�w�y���	'$bٳ��F�ҋ����xm1��}�
��1�����i�ז�sI6+������_j̱V�?���f��	*B�os}�I��b��6
>�Pg.����� \���� bp��1m;m��bA�ai�xzE�e�"�q��{�f[䰄:��[�W��aa�{a�	Y�{� ��/����ރ��f��>w����-n�:�z�Z�v��[R
p\�{��7��{��;Y�DM�T��!�'��!�$V$#�uQ_)�9���$
mx袠x \�M���Q�
'w�;��{tȜ�}w�(��h����/�Ν��8���U�ƃ�]z���F>*Q�k����^q��Mu8mH0x�b'��x1���9��ħIa�Oug������8X��UZF��&y�D(1B�(�-���ߌ�mT��x��H�!�=Ɗ��ʠ��0Q%gAf�����v��=r�E��7��e�A�4�r�qLE	��N3�Iy�'3y��P?�N�׍�=��F9��!����5Bu��G�$x�@�;X�����zӱ'I�D���_1�wR(�ܦ�v`]?�̑=2	i�P��u�V���"o�U㖄]�1����4�%j1B͋����%�N.i��E����bi���)C"��������;Qk�z��b 5%7<*�u�� �/�=1hA� ����MF2�H-ʆ0��c­��6F�ј��q�G�
FxG)�QҜ�$�}D,0�D�-�!ξ�² ���`�4���]rR��B�L��q�s����$�7���L3(��Ԏth�wô�1ꌹ1���z�9ؚ�������8�/v��1��S�`��E��@�++F(2'��w2��=�&���! @}�Z5ന�N���>�<L8�����~|���{?�l��յ�wu��<��@��x����ٝ���(�ׯ��B�����X��c!��'�䬉~�ڏ`�$h�9�F%�9/#y"x8u�a�L*��!t�n8&��u�;t(���+`�� =��J�Jy��\�L��vr0w�ٱ�֠���?g\�*8J�ZU�'8_���A=<N�ܞ�>��Ғ~JY�}wX�����o/k�F��V���N��%y�"��pn*�7�֬9������W��!���E�eY�����^����p/s��� �����T����o�����C�G�l�O'��BH�5Z�5��f����/O��Y+Q]k��L�����+#��t�xKB3�\1��ׇN��т�d��Xz�;g^��q<�&.�c�{ �:a��ՃC(ٹAe��4UK�B�`#�V5�P�'A欰���$ya��?XQR��6o^�x|
K:A'*G�ȏLM ���;�a�j�Q����J�~��n��V�-X�q�a�O`F]�|�O7ߣ>�.���d��)5#T=f�LQb9��v/���ĢD�>.H��9�F�K9���
��a�ǪH��({_8+/%4�I���O���oD�Z�dԙ�+�Y�A��,��-n��)Q�⦫
��58��r�����8�6�h����kܰQ1X��h/;E�՚��q��i:���OfV�5>((ל(V�>B�s�3�u�����(�XC4�A�D�'�U'�\oEE38Y`�Tnߤ�}�+��%��j;~��'8�n�硚iN:��vo��9����M2!��[���1U+��`Z�M}	ǔS^^�2�\����\|�e�٫h4V����6�\n��wpW��C�v�@��$\��v;��L� ��|�O��Ѷ7J���~��3�_��҉��������M�3��sa���L���t�}�]���s�0�}�ΏK��ݼX-d�&�_��N!��b� ��:OJS9����.���1
���~���N����L�6�$�3�tyu5����}J���r�=8��H��q�\�hٴ2bo$Mi�  �1���]�V�#��*U��@���Ч��|���R���r�)�d>x,@9"�s���`2yl�[����)>gu�)P�C�+9��Ko�� �R�64rJt�Kaoz�Dʍ�%�l�ʺegg�7na�M���mi~�Q~�5d|e����	�y�Z�Uw��s/X{3�ކ@�Mz+to�<WV���l7Nj�]`'�OQ9[6d��hX�F'���b������Cw�f�E�Œ���^k�B(��&̭걏l��u�ڨK��?F�2�Ž�;��Q�U��CtU���8(��M���w�/��[�KT�2ܰCI���0�x�3Fm{+wi��������yyiE�c���ݱ;:�Q5�IH����)iʯ�QX_X�%�B�>4ag��8sf�a#���+�^gCF@�w~5�Nx|=��9;��^�N)��m��{���0A�;1(���|񶋖ą��j����v��|Kcu9 �B���.�?��ؠ��ͽ�Y|`��b�4g��~U�
��ի���%Q�hb�[��js d%�KR���Ļ,����%P�޺�͚����l��ޜ��_a��rpt��0D2lN����`�̐�S���4��F�#�g�[�OɃw���/\�]�b�����y���$n	6�~��̤./�N�n�!�AA*ERr�.�]R"��7kd6��ow�� d�KiE�=~��J�w�њ�5�۬3Uu�.��>"2��.en������ð<�W	���0�߬8�Q'`B4�N�7*�Oڪ*3)�.��ڇQ՝�n�F[��RE���G�Y�!ogɝ� ��!)��A���,��}ǔd2*�dX�U\�#��FSD����E��'�q�A�;{Dpj(ʜ�k���.v�#_S.�e���8F�B������,K%���qP�X/��`)Plvi��߶Ġ��ݷ)m
��wh��k��3 �[�w掾CB�~�w(�Hn:7�	�=�%|57�!#q'�]^[���ۺ�����k9#w C�Ԫ:cٵ��-���u{��FAs�E���w���Ꝿ����8�lh�Ffp��e�Ha��>�ua�9�Ƚ�����@��Ш����a���8���	zwDy+�8fb�]�-\ls�D�f9���8�ˤ�C����C)(u��F�y��ÙPlŹ��1�j���n�L~�N�ʳ��p���힟(1�>��1J��'3�Cg�ed	�Wմ�>'�C���B�t
�IT�B��X�B@���mE��h�פ�XS!N�;ѢgwQY��{n�����d[?�'=�?|�j�p���t9�������I���%�[D{�����	����}0E!�~�:	�M�1$�2�n�RQ^�C�e���X5�U�ل��A���q@6tشȁe2�p�Gwpk�؇=��̅5�5#�]j3HCmf�4ŉ�R d�ALPCG{7�yȗVR&S�t�hl͋��tP�kd�rL�KJ0��V�`F�4"��3�2��-|�g��,ڵ@��&5)$�G�]$pw�e\w���u��ה�? @]r$��M�gWQ�iT巡oHx� d��sRH�Cl����ɠ�y����k��[�]��F���}�e�',Ul�e���e����Ý9�������0ޛ ����a�:�.T�"x��nu�7����	��Cłh����u�^ďS��F��B��!R���{�}n����Q[�ڹb��as����]a6q$r��l�D��0�YB�ᒬʭ=y�k���e�Su9�&'��.QǇ��#n��{9����'���/�{��^��AS��b3��3�	�[�������n�j���x��۰ (V��Y��zm����Lm�PA �q�h�Xu�1m��wk��ju]p�!��ۜ������a��D$+�&xF�W����5߷C�������oe��7a��^���DD�|�x|��J�φ*z`	�2ے��r���]�r������JuU��^��L�� �u|F��Z���Fվ�v��RC�-�`�����
��&�����8	x4���>=�����N���qu�E�+�)^-n��#$�7�"䘑iW�GX��C�_[I����K@��� jڲ�d(a�������bGm�v���X������.��7cdlD�)SO�R�7�
��r}�6+|^K��i'��/���=���b�5����j/�R�M���E�m���-_k�<M����{�)'}/��ޣm�8U���6��b�)�ի�p�+����25�A�α_�c1Y�h�a�����B��$���Ȋ��${/�=L��w�i��൨��/��e6����ZU�PQ�Q�Q*��i�oˮ�.�a�˃��β��t��Z!��g-����&�U��C�=�ó�?r9��H��:E���@m�|pw���
�pt�hmd�z}���=�<���gs�y����1�	�^B�s�{f/�Wy�w��F�	�J�k��#�b�Tۅt1��a��m1s����N��B�B�
O�
��V���w�>���y�����P|w��M��Q:���G��R=|<uM�F1�D5|�*3�4/�T�-4Զ�V]��R��lh
~`�"l���BDj+$��I7����I\{�~H��L����#S�R����vH�4��N�2!�T��R�!��у�oD�$w�$�0a4�����n��x�!�Ss�z-�0Ä=r����;)��b�"]�v=*b^���7��Mh��9G,�V�-�`ĳ,.<�W��]Q1=��U�ha���Α���"�������.��7���ݳɕ�`�!4�i4c?0�	f	%��q-��y�n�n��e]���$^��K�[?��v���+��7sw0��V�Z����H3��:��9�?�l�G��w��,��sW��#6A~�	hK3~Wi�.���BL��dh������#�;E��ӹP^B��� ֤P
��ѯyZ�`�"cd���Z'Ӆ+���9��{WZ�G%��/��y�qZn7�Sn�b��w�C�����;A��o^�a�����Dc"{ShЕhb� �#R�����a"���)I�����䐝������B�Tyν�2z&}��'���#��~�����܁��~;S\�0�'�L3i�S"U<9E��������X#5m�ӷ��\^�ĥ�>+F��+TGժ��Xb	o�=c�+��%�M�}k�t��%�����EQ5D� f������a����*�ZY:�0�P/DiR��-�5�5�I�{"kퟣ\V��2FƎ�^I�=$�=43#}M;�WV�.+6Ћ@�;E����$��xm�5Ή�!!�>�3����a�/���N�"5�8�!J6O���"��x�<�x�˛A�-;��}}uhɲר���`U���b�q����Y%����e�f��F�&TeU&��Q�x���f��@�`۹��:�+Ɲ���"!�u�,�vI����ɤMZ�!a67�ˈ��v�-�;Jf@�%F�2+�@��y��l?�i�i���Q�C�<�g��95�֞!�H ��
������B]:���˝~��n�$����f�W\JD�Tn9��s���"[|;i���h��:�� ī|4󂼟�kX�.$�Ad�nELJ=ĀO$�ٟM��É�NiH��Y��E�v�d���4j��}��6y��.�j�{��'�p2A���[����?eE����p�P��2[��]٦�2UQZ�*�4����QA�{����>��ˈJ�P�&
%dW	��m�<m�!��F���o�q��;�%�,Zܥ-�j�J�Z��8�	�~J3So�ڃbcg�w� T��xA-��@bR�����ސ�}��#��PX�2�p$õ�����מ���:�
e�d��D����Ԩ
�$mQE�p����;��G�u�wTA����uD2���"9�.����D,ʿ�0πz~C���*�O>��$<��;�XU]koF�ư����ъ�Q3����5�X�H��]��rg~�́����팋�w<�B5a��eC�AK�Cvh��0M��'�=�n/&"���nX���B]�("?w�q�0Xu3W�c����}��n�Gt���;��S7
Wֈ9��Y��n����4����3���[���U���0���ueg�������i)�.tB�9�Ye\�<e�E}��,A��M�X�u�)�ԙ'��Ҡ�'b�*��x^n�)$.z`��:�,ZV1�w�?��qM�)��h��=z���ks�)��j��e������r9���}ڡ0S�򡒃u��G��-ICQ�6ȸ�*SP�I���,����(;�d�rf�&g�j䌡��� ��@,�s�6|�5�ɚ�w���t��5"VhbE%o�0?4�1/�Iǀ�!�(W�3K��&�����E�Ot��� +@n����:���A���X�O`��/��j�'q�3���������kֺ\2�Z��k�(�`L_������+�6��|:��4@DΉ�w��-؟9wx���A��p�]�g���4��
�G+�/��/Ð�h���G#v�5̸�q��k���9?�	v:<oGI`���tB����IL��B��ͨ1ÉV�UT��s�r���ZܜT�9�x�<C&�Rc��=`=��c���������S����ng�� u�L�:?K��������'.�����ww9�����A���a��2-P$�s��/�uQ:{8�ʳ%$?�J=���\�
hS�� n��	���q���5�n�ɀ�,��O)b���G��_��y�r��}UT����>z0���.r��:�6��)3ơ�h�ms�N&ڳO֢LtukΏet�>��=U�a��NLR3����?;�qf=$&�W+�O�3 �B�M�iP���I��/S������a�BI[���C/�8.�&*�����t3!���N:_����GX\Σh�Q<�eQ� ��&+A�<,F���m��4+0+d�����Ƹ�;u��eڰ`�c=�䲆8��}|���o�A���崱�Θj�?��D�x�_�Um�҇iM�7Dy�r̉`x�8E��s��.�mg&��Cנ�tIO����L��B#�<"�������0d�۟oZd���1�� ��p��C�#���ʌ���B!֫�jb�&���}&i��)W����Tt'��2h�b�Mt+�R�|9~��w��t�+cNe��W���O�G�sFS�@�>���>��PN8��:����!��\J���������ѿF\8�E�Z�R�,Ć^@-Y����(D�I�����IԬ�O%�����_$8?��dH*;��1���:��U̘�v"
H��g-��Ez %t�B��������̕��Mhy.���L�Q1H��T� ��*o�������c��<*��ɫ�����n��5 �2eQ}:)�X�?�>g�X1o����"�'2��m��Ԓ����TT�cՏ����v�F�O��`3Gn��n)*b�YDѿ��9Ks>���D� �x©t$[�	-"~$�!$JT9"�w���	t��
ɪW�ұ'I#U���:��x3	��B�3�	����w0>�Q�41��G�g�9�|v���48��O]RH{�v���u�qN[_K��X*��ZX����Z���b� ;7�
QX�&r��Z���Y�ڎ���E�(s�]��[�oQ*�� �;妅r�HS�4U�����5��VESQ��1h-iku��Ua�EH�WJfYl���̓�A��0</�yC%f���I(�[m���~^�hA�����~����={_�﯏���??!òZ��/����O���y6D-N��A�&}G3z�_���-^O%Q9f���D���H��Z�P
�,���*����$zo_���	�s�?��\�SpH��tz*A�ƝIMQ��O����nv�������"M���O�P#�{�l������誘�7����WVy
i��R-��Ps�����P� #�`W�@���&x�R�?�'�_�R�k0A��W�薄j�9�9n�A�${mL*Q�%���ɠ��t�+��
�ÒB_�(�o�`� ���b<��?�l�e���qaW;���R��k��y(�Й��[ţ�|䑏i6>�C5OKQ��5|HHs�9�P-i��2���VDЂ�����-��*�+�r�J��n�/�f>J�?iUd��e�|8�l��N\͓�"п����q��ƍ��`f�����ps�'~�$��pˇ/ß�p�7��==���b���i�Lh���UѤA��/��aJŰjm0v
���Uǭ�]@�}9��m$�GL;��ڌ���53&��vm+�	NpH��{]o��>�������ی���7Sb51����?����J藂p�@Ԝ:��t�*pNu����]�G҂V)a�in{I3�5!Ǌ�y@��$U
%��Fchnp�Ax�P}�$f��5W+l�֣M���<�0#�K}8���R����w��^�_����2A� ���?��p�2�������
��OoG�\?��A�9��jU�T�������[����Z3�.���L$یI6�H2�XM�<���U�.�3豒���e��B��
�|�X-x\��!ςi|F��I9�ǟ�۽nZff�ބ�m�].Uh��%~��ӱ,;��-�-�;��ٿ�I8d�t�"ԬI�|� AΓ)���y���z�0��z�`� &�MLGVG2A�NA�u��H����P���("�M�1�I�\���sB4�!V�)��t#�����6+ ��#�]�
&!d
	�s{ԇ�^^����nW.��H�����s' M3{�~������
&6�#��J킨{J�Պ�fLf��r{k���F��dY�>��ދ��&-���&�̤;D�U�������#_<�TÄ�/���TW*���I�����"��u��#��D`��ޛ���8؛a�����/���s�`.�?
)M-�Q6M:Y����(�����-��@�6�d���ٳ����}�&�""�V^�q���	��&�WWA6�\�L�a^*�	�������.�}�hBW��o�#_��c9z���^�p���v��o5������L@��0��
˧UL*l3�D5t��ֆ�"�,2K�𝃙�qgl�H+��i����s�R��S`�J�bൽD���l���5�'��Ȝ0w~�k��O����F���7ɾL����mvƞ��I:��PY)C��]����}CLgs�E3���MuD�dt�x�K�����h��~�2�d^Yv����c�ey�zÃ�ay1ܻ� �����J���R�@Ά�!ni+����%�&����x�rc �:]ZA�M|ݛ�@ٓ������j�i�e�1+fQ�3I�|��l��h��¥�i>���	�VD%���i��/�_T%�,����0�7��L�6*�B̬Y�7&\�C�-�H���B[1�WO�Ș b�pe"���%�A�2Q��gDJ��gP��}8��y�S�W���w���󂣤�����C9;C��x�h}ɹ�yRO����2̛�ѮhB=dM@���ް�����Ö��XI�v�x7�H��2H�|�a8(0>	AUU���ق���$f�t�]'�ʚì�R��\����[�(��6�4���><�n�*��tY�'�~�x|<a�`�~�YdM�Fk��{�V����7=q�]����RV"X�#�3��>�<umY��&5M�^B�2��+}������%�+k�8@d�#��X��_﬇%���>��'��q���d �C�/M;j:~�.�4x�}��S��"���g$�5�8���fk%��Z���PĲ���g�m�y�~r9���j��tw���[�����5d�gl$տ�O6����IB>��;u����^g�g�0΢'��K��B��U/l(m�ڱ1�qa��D��MD���@T��q��h�b�_�� 5�C�9VLTP٨��g��%��~ُ���
i���o����M�p����EA���R�Lo�����e4��"&'�.�l����u)*�DbC�H!��^�D���K�y�gg��ڟ�ZB���'=�'|$���#���n	[���u������?����0I+�8�R������h<�Sj�G�"��B]C�FB�	62�q��
��ʻ�
`���J�^Ѿ�Cb�?��a̅��.�0K�9idJ�)�v7�i���{so���U(oޯ��wH�w���(�Q.���౦)^U��rf�3�L�g��'�~�ZoD���3�n�O��ݤ"�� �	���X��s���}���������,p`]�F����p���2#���r��Yk,��q�c�?�39_6��4��8>/��.kĝ�q&���/z�c��â�}�	�kb:��	n䄥�y��~�i��]���V-n��ho��/�<5����O��Z��9r�q��
���+Z�+v?�$Z��4y䙲�JI`Q�w�'�y�P#@E��.�l���>bnז�	9�e�>G�:/�o���z;ȷZu��n2Ԏ	��z��74�9�_l�n���ޡs�z6��_�����ئd���XS?LH)�g�Y%,S`���դt�ĮK���>��v�ض��O��50�k��S�HfL���?A����������Yh��ql��6X�{��c.����J&�Ĉ�c��2%%�h䆚��̲�'�1"&����߸ϥ��}f���n	�a�}<�Z�Ŋ�Z��`��`9�iY�Ht�}�*�`]�$F�2��E�Y��G�}��xE�f�-U�;_lu������<����vF��A���-i����*����Ř��d����R���Ϩ�2c�����w�2��g[�us�aaZ��8��-����l�d��'K��x'��Wh���&A,`(���!D F�GQ��{���V��쳥�������*�!��i?�����z�	v�(@����T�����,�I��Y0�%����Ed��F˿���D� 1��H���>�����~�½f��F���_��rE�0O;�܀M�.��\]����7���Υ;��!�g�d�-�ײ`��Riq�Mf��t���;K�I35�a��8lR�ϫ,��Ix&��X7K��|��./	8���C0��)v�#q�y�hHs9(=�ӕP>Iw�b�#��1�Q�"�TU�#؍d����9qQ�xA�x'A,)g�ݏ�0�g�̓�y�\�=Q��I'���%;_\�Z��)u�M��w}�8�GI$����BDS����r��	 i�V�C����*���
;[�Bˍ���<�m�j^u�vZ�C�h����*�l�,(���ZM��i�l0�l��n��|���a3�;Aj���@m�EK+�[������`���#f����}�cI"7�*�#�H��RW�@ҹD�Z�R���UUZ�zǣ��E���A�㈫��@|�c�4�,*�����h�.�`Wb$z��R���W������R~o0���d��1���eϞ�Dp��v�d&O��Y�%]G'����]'��q�L��#��b��!]0��.Lp�t�JݤE0#`�J-ᐁmߤp�e|����Iİ&���a�Wh�r��7�%�]���Q���2��c)��~��z�D}�x��P���D<�,U�b)1�M�M	��$=ʆ�_��\'����>s�I?P"��^�~������]�v1>���c&R�{D�h�+ɦ�1R��G٩&F�_CV�՚����a7�.�5�"�lo?�R��H `�)8t�o�E(��
,&Gã��s�pY��g������Zc�Vj���
��3]��#��[?z1�
��Y\����Wݼt�YNQd1$+h��Z(��xu��gI�P!c���R�He^�ن����N�@1���z�nu5E�\�j#a�0��W3��SAy�&wA���^x�O6~G�K��~�Ξ���˒�?����cz�N����\_]�����c�����/yz^�	�FY���:t�R=X���S�__�j�9B���I��9��l̕?,��i�E���� 9@ƿ�	lll�"�Q0��X0����N�uV7�^����]��w�N���ң�wy���
�On�&28���c��z{kCK��D��� >�p����,YDk�z����L���+(��:�u�ߍ�\��#IH�g��-m�f�30���#��\��j$�j#��D�#��x�w^���?���wqѫ��*��V���&bj�FX]�(g-�S���X
�(e�y��mb��dU]�`� ]"�0$: �2"�&o�k�$��͌�tm���bc
&��q����j4ܶ���2��t�u9/���٢�d��"��uC�E?���$�hK���#ess��ٳHNla�ոw��{����u	/��b�$�1�S�=Yӑ�-Gc;}��-�/X�T+�"�ڲ��>C<�}��?{g�^�b� V�qp������?!$F�d�Q��¶��º�
g�C���n� �,	1��7���%<��G9��5��(ߢ����������������C�t����.��
ȅǪFnLίe�˾�?HL�y��/�^�M��&�)�_�.���T��
��t4�"&D�z��?�$z������cQ����$l�C���{���ە<߳�1����2�gU3�1m(WxG����f:!�e&{-gY�E�/K*;�`��t��Tۚ����6�� r�����U��<rÞY��!�^�ă��Vf����ۙf.N#<�`v�����������!N73D�^�ӧ,ȗ��M�8�s�;�\�ʚ��$*�/��#i�!�����i�l>%N(�cTY�U�j����BhP:B�L�P��؋��Oc`:��e�Lٗ��"а��)js��xΊC�"z>��x:�</Pq�U'5{�	s�IB�Q��LHk�x�o{ea1-0;A�,CyHz!���GO"��l!yn*e����EF.��ͳ�a�(�����+����8�n�0�\�@��G�2J�瘏(Xs�<;���pS":}2	��eO��T�� �w����?��'���"�GF?m£���c3w��/��Ͼ���k��B� N�s3c�VM��L<�G���@E?p�p�qh�E��45��b�a$k�IU)�	i��:S�ߚ3�V�L�5�f�Dm"�s=Le4=N~�U�4�~_�ɱ��q��,#c<�1�%��&��GU#� ϗ����V���ot8��2���p��ڹ�f0�*��٤�Ն(u�ѮU�b�c�\�źpF�l����5v0���\�F��2����lc�ҵfX����y�/S�4�9�`~�:~���=̿��x�^`0�G�O@��܇�}i	��� 	����A-�����v�v���+ʃ��5��|���M���M��C����`�3��X���H���~Y2m�C�خ�f�3��S�����4���<������~-^��`�1[KLM.9	�KR�i����>/Q�2�6�O�c0L1H;��
�$�񞌎x8�+D�	����H[	2���� �W��h $�Y��8C�aT�Y�D	\Ä��f�Q7��b��Mɛ�1��g�+?��v$B�wC����o�}�ٟR�э�l@i?ʷ��[/����������pr6�k<�yvL�z_�P򪰕����N��a�D�q��`��(�(O�?�w�)����^s�! �I�+bY������e�_*�<W��(�CY�4:bh��0d�ϕpу��bL8������^//�������$QmYPλwF��7W9�uc�<{S{a���A�	�e����P�Z�A}�"1���8#B&̙�2,��8-l������ï��߅w�<��,F��9���X�fZ����m� �1�/p�h�>���$�l[G� �~Co��9��֍-�2	Ur}DA��X7g1���T�7���g&��[\ׇ��'��AݐYTc<_`:[��}��3���(O��`
�~H���NG�l�(��ψȯ�!��}&�Y-?'\�e�4���u!4�^���:2���gc�L�S���M��Ў��LT.-�I6����8I[�c�(��U&ǖ��F�1�n�*`X^'��:�>�_���O�����=*���G%��q�]������09��0>��x8�>�g�N�e��Ţ�d���é��ll�Q��۔!K�s�R&p��m�4*iϻŁ�Th|T�Q�J����n�$��٪:��0���ʪ�<^;_�hI_���ٮB�ÏK[IK����6�E~_7�%��R~i]0��� �"�r^��BF�P8�籮�u���y�.ZX7�K����²/]�jc$�֖��X�级�sfR���,�	��x�w��_������]<�U�SxU&}�r�6��K�����b�ĶKpTa�R�)V*&�c,�u���X͵���1i��L�6@�Hǜ-���T�n���؞!:g/0��84��X�`o��i|I��T��AQ6�,2Ng�T�C��Z�/g������ȲJ短%�J2�M���|t�@fFxEI�@9i�St�C�����c� 0��Yo�ir����ҨH�ܲ�L_�P������PШ�JZ^s�0�ޡC�\P!a#2�8O!���
� ~��/��ף���������%�G�f��]���:�'�饪�?>:?s8����=u�����F�7���8?*;T�f����z	�l��܂T0W�(^b���&Ҥ+�;�ڂ�gP���B˥-çR!��
��*<R �����i6�t+Υ�%ѫv�8�w'ӹ��(��顔g��ő���ƻ���Q,k-!�G랳�s�{��֍���9����;��[eԩi�������&�.��L�Y�Xvrti>�Ⰷo~���q��Ც�3(��ɥ���K s|C�,��� �.��ɜl�Y���5Q'�Ik�d^�rct@�P��*������f4�ƌFU�F�i��G� M��ҿ'D�Hz�F���T)ÒLe��;��,�p0��A`$c",%���Y� �v8���	s~$I���B˜c��%5��,J��� 136��CT	��A��.�-�"92�L� ��Y�������M�m�[f���\�93C���a���D&_�q�B� �:b�6�}�l��!J��)�n�q�6�����kх���&j£�����1��F��?����g�G������&�sEYn�Eѯ�́D�,�l��(�����;��K3�ʉʗ�gp����|�i����x�,K�����B�27���k0,)���w��^:�v���H�NG</����T�Ua&�1�L�JBp��DO��e�N-PsJ}�6��
Lq�z�a�Z���#w����.�,�`�-���x&?a���j��4T�\榖�L/�8�������?�y|�op�^n�I�RINs*I�v�m8�$�	=�/�/��F��?��4`kP{4�K�Z�����,�s0R��T��F�;�/��u��]/� ��=�<3M��i��ekl������5y�>�E���X�"ɕ��/�#�߼8�}��&��^Nnv�i'��D��Y �Ywb@%���@�5'˱w�]l�ԢHљ��d�ʰ�'+�%�c���.
���QK����1(��⹇�\R�i1V_�8����!��@7Ţ�c����<��O���|���'��ô�QI��U/�/��ivi6�]��f/�'�g���c��-��ۨ�:��M�A�^<�A`�p$L!z��s�;j��|�?�^����e6L7K���-rQ�d7���0|�\v�$��t5B��2���x����� �P�f��!�OK�W��`G��$�w'�ד�뿯G�����CNǍ����4k�8�4�3#wŘ������G�kl�c����O���~jl5%8�qY�&t$z�� P�2)���dE�Ycc�-��`�Ra��L����V�I&���[� �k�K�u�E�� �WO�{��6�,���]�,��Q���6'��[���u�(M��tP5>k��.b���5m�BXj�$u�@���X-6�o9����m�vrDl��.�3���Pޫ�c���!q���x\C�؇�
�s�h�F�J��0a�F�6/A���9cD�1�$&��ۈ��V#�sM���|������A�ԏ��-�M5dta��o<�C������W�zi£��p\�,o2AZ��D�������{|z2�}rQ�'�,��u�k����%]��g6g>�����.^�g?��r��*����D^2���̦S1 Lr2�ia"�J��4�>��˪׺0ḝ>fxʆv�� �C�隥z� �a��e;��n&�x�������â�FZF
��x5��%�	�X�,�=B�tON������v�A�~����f��]<�W�V�4�����J&[es�����F��!�!.��`�Q�Kz��D
�Ls99c+{9k�pB�A�kL�s�1�@I*ɜb�7-��I���1�����Џ��28 �c�W��ŵ�	��	$0�L�\ $��@�NJ�#_�X}�K�����T�R�Fj,���ў�_��F-y���2��L�1�y:����!��,}�$ �N��$�yH1��s6�_념��T��\�H٨��%p*t�i���N # sx�*NQP�qz�%��������4�n=������|�U-Bk>��A~�Z���|>�F�u]^�ϳs>1ϟ(�b�p4N'�YRTM2�L;�ɢ��zx�/���3��#�L(�,&V)S�s��E�B�0�:�(E�g�:�4D2E�]1Z�~K6�L��u����"���1�P���ڨL'c�_� 2u f��3�0<�����1	���^��Hx\O	<����P�J�Ք�%ˉ@Z�A��gY�����g����=<F(FZKBwd�8�jXv����A�03LBU�gn�U+psLt�Fk2��,B?&2p�sd�Г�`RW�)�\>b��PT�BO!erTit�F_y�B�XPʅ��1Z"k;���5���A8Y��s�����I��WwU�s����I��ٱ�a�sXN�$p�8B�A��p�����6`#��2|DvlȒMIuP�(��H�\�Z��K�3;��]]w����f�+������k`1�35�U������~]��=D�
l��|W3�贠ǱE�͇��D�^�w'��Z1`@S]���&hx�����H��D��\=5�tA̎f:����(����!+� �FH����`y�@�I���?�(	��FQx�4��@��XV���ч�����9���"�fy��i�+W��;�F�B��Z_�Z�-��M�m�iq�������=R�� �i���~xцR��Ǆ@2���0,Ve����Z�T/g��L �+��U��i�9����f��A�(�~pCj���07D�f�mb��2�E��\=�f"2�c�L����iQI�=� lT�Ƚ���/�r���C�矑���#�j4pt�ecT��Z�"����	-8"�t ˄����tǍ�w{Z��^(��#�9"�e)��Hmv�p�8��a	�g#f�H����!��
�K�%	��4�*��Zr$�iF-'���\�J�H��*,�*.稉�Ϭ�t�C�6��n����ʯ]�W�e��b��q]	Qu~�n �.�(+Z�ʜh٥�/�ٺ���E�w�<�Tm#�	����\��@�o�7��5�}AB���et%�����S�P�[!�YV�p��*VWe����+g�������ԍ�@�t���@R�
8?@���?��a���@D���l?��^i��W����7��(l�oH<��e����Fٶ�^@�>�NH*��x*��5s����M,q|� wU�i��`�0���Km�-��ؗ�ǟ��?������e��M�B��	jH�T�Vb$��2t�����L2�s��M㥃�٪�m<�I�Z��i$�@��8O@2 ��ʳ�y��V�f2�G��]����j��� �NE逴�6��n��S�!��{Ew���I�{$,h�i}b �$fTGH@hub �:�mṐ?���T%_rZ��c+>�u�k�8J�*�h�	���O)��y��<�(54��9�G���\&����$$�V��ĴU_^�����d�s6!쀅��x
�"N�����W~9+�w�3K�4��r���D�$�L�e^����F����7�n6+b�06�Bg����!Ȧ���(�F���6O[\mg�V����Vj˨݅�"��E�=�8u�-!�.Q&f8�Z鍿�I4��X®���U-�H.��|�C�[�s'�X�I�H�����_�2�9`�� !���.`@����U�	�c�`��)Qn���h�	T��+��D����ش����Ъ�V�,��Vh"@b���U�O��Q!`��xba�\6\C�Ο�{o���F4�����S+(��g$�u{�A7F'f7T,e��"I�7���m+��a=�kL�|�BЄ�Yn4�v��!��|�8DG��� �������\US ��$`P����R�=��
!�Q؜��mo������۵��vEv=/*�+���\����WF?�z��E��6oh��H��Z��-�@�K�_w�mR�$��0��Z�l��43tnw�܉q)�W��g�>�n]�j�ͅs�9�l�l�(6�F��cC�ڨ@6��3)hƁ���Z-�j�,uc�{}�w> ����h�K��(MM>�����zJ��Rڐ� �0��1�"P���Q�,���?6~n�)ʦ�;�X��<j!������Y�qh[5�^P��vU��q��sģR��Ip�*�9��;,��!8��Z��J�h��Xq5��.�B&0�aK���0!�σ�A��`+�� [E�pmL��A�v���j68$K ���*R2E��YİB��* �Fۈs|�qƹI�| H��/��~,M'�H������tph���Z^lBخ������=�:��/�����ʲLP���@r�����!�r�8h��	��@��
T�v��Da�x�@���Y ��t�:2��ܽ�<f�B�3�:Ql��Z�;m}����kC�a�5�J"!Iw���`�mǴ�[�u�BRkA�F�;���x^��w?$х3rcH/��w1WM�$r.�8o%jIc{$��p�"��U��%�1O�L����舙�J
�A߇�a�p_�q�H!c�ʭѶ�D��d�됸��� �5]b�w���C�U��l��+@�b�h�@)	|����.Ґ�����������t(�M
�?�oHB #C&�<��Q�&����$�t�Z65&�P2��V�@���rh{�wzΈ�#��H؍X!��"��:�B��]�e-�oy���$�o�i�py}c^��Z�t�����y��ϭ��#��(����M���3!�Y|�PU(:�&�i���
/�l���p�ܧ12�3�Q#��E�����	�`ބ�nV�'�V�PZ���z��ߜ3l.l�8"�����Y�l"������*�N��� 
er�e����d/�����@[Yq9�����ܳ���٧ `1c~�^:}�~�29�E��!��5�nߌHu6+(�����q�鱻��ɹ���bf���4^j5�L��I�z�����c2mBuY��j��&8��u���$A�)����׉%�.�f@�b�t�
�X8�eE`    IDATB�bl��YAB�X$�4!��o��p�,lT\A0�������ݨ�t� 9mT6�Vj���z1B?�f n�!O���۷<��O���Om��a+���.~^��O�<�#�^>�c�I�β�N�l��:��� @R�ӏ�Qdm�܈��ڤA��UJ��Gv�,����r�kv���a�n�2�S�w��Z��&&
�Z��Q��T#me�Q�6�iǿ��M�JV��ȭ�x�:e�*_��?��O>!7�cY� ����4�k��5�bo��=���i����a���PI0�r�Y�I�\0A�*��6��y��p�h5�f�,���	��r������������0tB�ΕI`F�)8	�����R?T�AS0}]"�q�����t���w�0(B��M`�d�C���x}?�e�������}Aˈy�$�!`^��
��"r�J\�=l�Մ �1��{O�(��=H`G�v�o��{��,��ݮ��&����y���\��X]_�u����Iz�x}����d1Mӹ��<,:*`�I�m4鍬���r����A�����j����ʝ{K���!�İ��[J��n���!S���������lBh���o��&3}��۪`�Rhg�����}}W�i���fU���O��>"7���42!�ږaB@�]~�rȮ^ϭ�(��,��T�����t����!����n�ڠV���c�M��\سWT��X�m�&��F���ǅ�@^u��P|&Hc����}m8��x�kb@2 spT��Q`c$y�Ot��BHh�'R�X4�ǀ��C�V�!��=�� E� ���Lkм[�:���(grUz��lBQC#�d�����1	�ˤ�0!t�.eGX!D�LC_J$�a,i�{����{���9�]ˋM��7��6M�-/K�(�G���n��r�ޕ�+���F�^Z^^�p�R<�摑�@U�J�u<�s|��س��2z��E� ����7�E�h�J�`6�
��$2<�Ѱ����id�(4�a�Nd
�U"�����n��6�ƂzU3�7�U�w�-4����|9<7'_���W�⣲߭�@ Q�LB���D��wC�EBS��-�Xue��H�e��L�h5��c�2�.�n�j��*EU ��S�q˫��c��qSH�����<�w[���ص��V��r�#��ba$�:C�SO��}����
�F�~��Ԩ��ܘ(��Wf!g�\$p!L���;AĪ�;M\/����M�N����2�G
���_�
�!f��|�B)<Nkd+!	i�!�Jit����΃�5�X�b
b):�d���H��>�>�qV�ky�	a�"�&^X��F����#�����x�T5e�4�[W�2��4n]~Y�A��������G��?�N;eY�AG�%Q{H�( �A��[��t��vX�Y`��"\u���h��#����|�KU����Hy���c��L"3��v�&$�Bg�uڷī��'Aj+�������׾,���ߗd}E�v;����X���p�0X��#�&��tj�ר��BՖVN����(�Wkݕs-6rX���(Y=*$ѲP$Z+U!�[�o�Xa���5�.t�����ŃB O3��mĻ�9�	�5AӨ��g��4�$�<ɣ.%�=�#}T��{�3 >X� ��tV������G�0��'E��Q
�m�)J��b��ZeSe�(�\U=�I�ufQx��JS���;����� ���ͨ�PY@"&d�e����¯���{���8��l��&�m	�}�׊�����{�ʠ��[]]�2�L&�8��a���/\������G�M�dzd��{�q�b��N��N��Z�i,
j!��!���\dz��86T�q�`�x���?k�Bh���	�ռ��B{\�l�Ntӫ#���Qp�b��v����G~OV�?.7�V>/�/�=��
"k��	����y���>>w�&!2��~�WV\kMo�$r-�j�ZV��=(��E&^9%O�EU�sA��Y��W�����,f���a ��=9�4e���?�tv ي�$s#IaqI�Bȁ2�XT��?��)��m
(�		!4���i��U�N2׭1�ىVdLj2hXhm��A2�mqy�HTD�=��	1�5�BB�v�Z!P
#�:
%KB�v����n�ws����8��ZalBخ�����D �(8e�Ѿ�,[(��|>��E�g<��F�/./߼���XU���(
���}�BE9�%os��^�f�[�4�iw���^	H K�=�ĶY���3nүrX{��`�Jp�
�ecPϑ�+��#�s���������2�Ū*�B]��ɘ�v��n!��0+,`�����V5�!����$%��C���Mxi��dcqav���,ж"��$����a�a��s0u����$��a�϶TN3[Rfp�N����e=L��1 L4d�s,�H:� ���&T&�=ñ�i�3$��
����4�yƉM�F��&�93PkM
�c��*#�M�6@T	��Y�HIܕ
� Y�X)���E2�]$��w|�����>�8�:m��&�m�}�k��rY]���˷\\^�c�:�keu�Nid�gP�U7��n]�@Ʈ�v�!��/t����``X!�|T��v��Š|�4�����h#}!#��R�$Q(���+'�-_~�c2>���Y�Bqӌ�$���-il:3	A�6�ID����
�D>���SW;H�i��-�B���	�p@p��Q3��4e&N�k[��A4�ݓy�m������̢���9�^!¡�8�R��٘�"Gq�X0��톒��\	�}�3�m�NR14���֓��$u ڈ�2~`4c MV}1�<<�Vh�,8\���6�A}1Q�v����6�F8�E�?�:�&q�t�s�cZw@X6�3��0k��H
�gF�L�����w�����O�M�]���-fx���.a�_N��2[X[����d���=UU�t����4��e�����㢨� �0�]����3�B��L3d�M�������Ǆ�b��$+*�CH5�D��|����|F�F�x��� e)0���J-8CP�9:c@��*à�Bw����U2D�;W1�0��`��|"��Z��"p�rV19����QV.��[�	���B����@���j�Ը� ��gB>�jB #�d�cq"+E�&�,���A��֮�
� !� 	p�c�Ǆ�*c�����������4��+�7Z�#��L�`��xP�U�L��eu�_B�4T6H�4I�ʨf{���I��7q5���H�Ns�2<������;�7P~���u����V@+�q��i�w.�ҟ\Y=p�����h_Y�>p��iy�*�cU���fP7�)ꪃ��� ���Io�^��jg	��#�'5<wB��mTIz�<�O�ڋ����������Q*^ ���m%ˡ%�����Al%�A��fMHL�pgVM���	C�C`d�Q1��]$�J�\���TW	�˙%��,�B:��,�,d<��]y^6�K���_O'LN>��+�P��q�&_Vj�K賃3 � �c膡�Q%@nm.��Q%EB S�T��d<�٘��Zɟ1|�m<�I@�,�V���T��_Dy��p� �M�C���K��n�` p����ՋdڍV��y�/t�=��s�lµZ}���" ��y���.��i�����lR/eE6L��eV˪>������AY�ݺ� A�	<��ۅ�E,mp(Z.�Q#E��:����8��6�\�o?�|��J}qEn�K��x>� �>�!��ɶ�*�R��j�l� �XErv୎R�������*y�t�0�me3�44������aG�ݾ�������o7\��u�c�PW2^�"��HҬ�0����p�Ҕ׉�����HqG�ڑKU�v�@~�(bB@r�� 3����¿ �3"��S�[D�V�Ր��k�Ϡ��v��EO��+�k���l*�J�_��װ�4	A�8�w�TFB ��ф��<��Ɇ��G�q�����Ƿ��d[F�a���.�{E$�,��r��͊|_^�K�4ߗ尬XY�0�N�uӯ�:bҨk$�~�hix�t��󀆳�Z�{��W����<%'�|R��u9��� m�tB�>��E��-z��n2 ���~E� ��c�
'6_��:@K�(E�>tv��k�94m�̠}c�ǪhZD��4��� Ҩ�e<Z���5�|Ch_����f��7�Wd*�]���>MfP!@�b�nd-㋌;�|�Ɖt��"yH$����.14�#���7*�VZ�	5����΄k���1 ���q�˚�T�?���*g��B
0�}_���z����+yVK���2Bki)��؁_��v�W������0ل������� ��gE�ΪDU�v�i=_���֝��)�|����$;Z����t�i��iܮ'�@j'T~v��tBO&+��/I�_8!�@�E%��&�$χy�*��l��	$(j)ӌ�,.�� J�C�@F�'@��;���J�b�v��6�(�~8f
F��Uޜ(�V �l��9����!�Q���_7�M`�E��$D���D�"���1q�����=�E��Z� ��;��J�2�@F´�h�c�k忉�2�!���D8��V�������1� ��E����$׎R�H���6@Oy �AI�������G=Jd;I��Q�#�ȑt>\_�����w��v�M��Mo���^����AEE�뒬�Ӯ�n�����Ln\�Lo���H���M���t2�������ҋ�7l~�ʙp)�dOS;��Ϻ����q�Z�,��}�Ek��
nH�jr����gX �Kв�[��6��A�b�p7���V9r��m��&�L��� �FB�s�B��Z7�t�Nā���X�\� ��I���$�p`�E�ű��LkO,���P1;�>���V{	��lf��^R�_4��\����*m�n�"�C-7�o�Ti����C�M!W��N����%��ݰ/�ēr!����n�����^���M�"��5l�0n���#��*�7M�=)� /���ϼ��G�����2I�� O�S�y�@^s2m��ɲ�������O;K�'�~ф��By��P�<,� a���0U���V��Rh���Ö�ym�7��Dd<Z��ш$@��8�"N��t"^���
�`�4���C��2_2���L$-�vݮ']�۶�
�eǨ���8�R��!]���Ӽ��f$�)i��i�	$�i�pN%bE��R��A5���뱺	��4�wbɺA߰�����:��ſ�[�o|�M��'��6 ������>�������_~����u#=��`�]L7�"P$ID�_uNS��Pr�
&��ʫ2g_��h��WՔ���APΑ�Sj`7;�b�H:�X��f�Z��T�ɘ֫yY�ﻬZ�t�R��4�ΤE7��	�l� dBH��k�e�2�;�������:H����{,�-Y��3h1���ZFRt���	�u)%����1S���H���|)=��(JxV�f�ܐȈ&l6��0qNV=�r����-�On����IF�}�ڄpm>��Ul�khF��_���~�G>��_z�{��x��A�8�q=		���`+��X�he���W���p,����][$�=h=��� ;sz�o�F�;�M���"a3��X���6{�F?�\#ͦ:�|�|^�S�Ҥ������ r�$m�2e�2��2d����2�;�����8O��o>�I�g�j�\#i�
&�R@ۈ�HTb��2�·�~JvkB@�@ �d:�9���M�j�΄��JpB�b|��_r$�=���Z��������w���W<�M�*��ul�� �it��_y��?~���]8y��ѥ�{��z���T��UUr�t�Z��יNٓB���~h�J��'P-(���.��I�I� ���k����r6�#�<5���a�/����>]��E�j,�E!N6�O4t��#gB ���	#)݄f�����A�yl�|��E��Z��R��h^��=�ӳ��t<��y&:��G��#�ǅ:w`" IO����:���QP~$C�tz��
t䯓���i�t�ve:�W�����w��vsl��]�`ڧ���h�&_�07���8[,��R1���|�S�ƋO��~�ɧ�'{�\4�	D�Г4�
T����Nm#�C�-&�jٷזiД�h���Rކ��Cj��Fa��	�Ȓ�x-�(�<8�Q�R]�`G3�e�x2�cMB� ���H�z�c��:2ZDd+�2}�4�t��l-3&�v�1�(�]�����\&���W0	<�ل��
zNp.EB�<���� ��~ؕA��
�R)���B�(T���(�D���;��~g):~-�_�B��Ѷ�e#p#Мk������#�����9{n0_�����\]��ߑ�,���(e���O��2pILS>�Z~����AƢBikzc�0�6�V��,�l��	h���p�[��2@���0�aB��N!9�b�6�ow�
%�\I�`�h7a!w�9�,ĉ_|T9���F�C�0��|6���	������**VEF`0p2���&y!y��s�U�d�3��ҔC	� �LD��i�=Y�������Ag�3��o��Դ���o_�F�F`�"������C�{�C�����L�2�Bz���W�J74���,(˩��D@q?0v[�N��҆�Fe.�P�!�qjC�`E`��[��~�>��'���TT�z@�b@�y-�iF##��J�b���c���4������F�8E��%�>�\���c.�h�Ln�oCmY�02�I�Jh�ʂQC(��V���e%Y�]�z>e�A@�ŉ�'�D7_�������R��2���ѥ������g���Ok+�kq�z6�0�������3���O�O��!����q!a������5���`-� �u�J�T���Z���,�\�I�2nv3^ֳUj&�P.ą�h�/�)���v$<A^���~�s��	|"z"7�#)�@RWd��9�6�-�.� i�z�w���W6tG�\�\1�������K� j��&!���5���@J�,%�Q�䅁1 ��}���&	��w-����sd܏.|�_Z|�]��8s۵|؄p-�m_�F�G P��K�^�����S�|⇾������7w�J⺖�q��A;�wSxK%i��"���MR�N��JMmټ��$Jk�T�ecg�c��0d<��Dá�I_-1!� ����,���2��IV�*�B��0���ɸnd���-iʬ����?O�^(]7 \V0�F�dD�p�` ���P�TF�jN�^�f��1D�JV�
�� �<�^ғ.�:]J��ZH�*�`��,�J��w`鑛���/�����U�r6!\���״�h����=���?���<��gޙ��x�YY�!�(�\D9Y��4���%�7�;� �� ��W�uk�V����^=�\hL�h[I�?�$a����$�[�ӗ�#�a���j�e�N�8Kp�s�j�HP^@����eڸ2Wr��<]��E�|�N�I��_��u�sT?ge,#9r�@��M��ϔ���s�j -s�� �9��B>-"T:�1�a+.�|:�����Ts=)g��s�_z�]�}-d*^�-h�u�`ڗ���h._�������?噯�-={�`5^���� H�����E*n�Q<��4�� �Z$b�`���7j{m���s��E�6�6R9h�&�I0�w� �"��j@a+i�L�4���h!�� �l�� ]�#�L>�o</��x]�aEZ�$�+]7�<0 �@|3�u�A@�c�PUe���~Q%�V.<�ySKڔlA�<
�']��8�a��84�ʏ1H�8?��H�$�ji��o9���r�q�_34�  �IDAT����C���'Ӿ���u� ��_����'>��>�������[�ӯ�Ӊ��5ܔ⃴�a�	 ����H`=f'�u�흶%3k5�"}|7 �7��MoN����9q�P�VY@O�T�,��6�0`��I � l�P ����İ���+w�6*��i$�@b0�=�#[��5�Ș3 I {kJ��1�b�t|k*"�hm(1n�ӓ~�HR���sp�;��Hd"�HőTn,E�+���z𮟏�����q���et�o_�F`'D �!;����?����K?�◞|p�ԩ��d�y&	��i�{T�*e��H���q�Z� ��"���J�t%��#��q��T�.PUQ�[��������#_�<�xn�W�#�?wǝ�M�g�Kd��l�=��HF��It	ٛ���y��]��Yw��{������y^�x=�[,>�QI�r��4\tQ���u�dX4W]��}7z�����S5��)�	�,���G�a.)*�c��ʭ���T��j���́݇$��
V���?1�+�F��xH��[���o8^���,=�h�������М�W�+1 �([ŝ~�w�$/;��h������g1 �m��q�*�7�-(J%�k8�CIE���)�'ԶwP��X�	���H��H���=ڥe�c�Aɚ�!K$�m$ߤ�*I�I5�G��W
J��,)
�e
ш;�zNI����`�~D��Ԣ���ӥ�J�����X�o֠���m��C��4�*j�^A���FJ�̓Nzfm��a�.%v{ʔp���P�2��飑�`�h&�q��R ���gnm�\l-�ntŇ�}�~T2�r����]8Uu����+>KQ�7�Ā.ꡀL#����V2{������&���{6����Vx
���\3Nzl{�II!5���@����d)���u��s�$oq��s�_���c����w\�]�;k�����32H�e	��H���/�
�&��w�­��T|^[t�5����at�kXow�^TP���ꅝe����>�p�L�M��l�<U6�f
����t�������!��h�sV#J&*��P¯�~4�)�'��T�i�)�']�k���GqD��� �G���,���(�k��s,��ӳ�R��Sn�+V����G�{ �E��NF�h]Wx�1g��6#��))���F���o�n��#iC掌����~�:�ƽ��H�e�:�s�xb��M�/�Q�yD���c�t���>X���:�9?�:�X������IF6��k�Gkf��5]neE�N��/7��ۮ��ZY%J��Cu�cV�
�ǯ��iTO>��)�cUL�ߗ�>���ţ��o�q�Q� �iF�@��6g"����� Z9��
�S��Y_�!��xL�
�3�/�q�gg&l��E�"�pDf�d	f��)޵��
��}�ʄ��~h���G'A�J2?[I-�`�����	�":���M}Bܷ#3�<�qj^'ޞ��3�ߋ�;6�;��-��Oo�!\����̠E���jP`C��7��r���GR,��P�J�D��g���8����7�0O)��V��<%�.���(J����K|&��5�e�*���*�Bϔ����A�%��1ԜN��G79o��k�u���M�a�Q*����΁��`���_(��8D֛~awv�h?q�k�=gX)Z�Ż�R;���GI���1�''g6��W&E[μ�ζ�*�S^�*y5��'P�=���b�i~ߞ|��{���rT�j>[���K�u48>h�Af4���[{��,� ��g"�[�u�R�W>�S�hY:�w�LlAP�x�ehϕ�L��;]y�F�":d�}κ�r�����B¬"������0�g�9|iF�D�5�>����m"N3��Iav�[K�*�>"+��^���J�Gq��8�S�����u�v|0�xzt�O�d������Ԟ4�+co��t-�����}�����+��L�"�X0*���WcX|�m�̽cɅ�{�wp:�����!���&�{⦛ur ��*Uo�����)0�2h4tg
	<+ATr�M��<n�b׌�@T��H�m�j`S�b(ШY-c(׼W1Ƀٌ���>��V{fP�P�o��s���H$�����	hS��Z�ڎ���F����Y~ۨ���c�"T^!a|!&)Q|��wX���,�@�V&芬ǋγ׀��I̓�~	}S��x�5^S�?�:m-�B���J����0���M�$�4*�%���i�IN�@���ܱ����+k�z�|����jX`Ă@����_��^���V��De�:>sC�k�g���//!8�hG�y��"#*���=kX�����T���IX�˓�����u�@���mx_�n�U����2��2�;=Ʒտ�.=��r�1Y�N�����ҿڇo�I��NK	���Q�[�w�{������������=��L�F��"����Af`6���7��Λ*����uI�q�D�'�=S`��v�ډG�8�! ��q�3�NS9��!�~�uz8u��H<��r���y������q���A�+x��|��n��\�m\ؙ���4ӽWY�/ץ�fG�o�3�:�ee�^�w��J®Tѿf�}������d�9.X�r�s���ʴ-;:7\L����e��ugc=/����nb���7T:\[ٝ�k��;�3��h=Y�1W�Ĝ��0��:�y��\DRa���m{j޼xEWa,C�h�_�� �@�����!�RF�Y	�ݙYqm܊@WI��e�m����w:1��:�K����͢\�Q�)(�T�m+����*�<����љ��<�����!�h��ۡ�ݘ�)�'��{i��aD%f���\쌺���j�r��2��,@��Wp���6���G��zdO�h���>G�v���'�����b�B��{)b:�0p��D�RoZ����^���f��l�&�y�oF���2��.�PF��(�h?��h 3�Hs�>IM2�CM,�,{��1��I��y�A���:��X��v1�W�!�[`HV����x��P����T;�����Nr[วϿ1t��d��6�O�3~㺎j�%_�� �&��ɰ�����qX�D:��l�~r�'�$�E�>�������$�F	��0ao���ǀ��'� ���f�a�r�!ҍ����OVԅS� �cy�r�8��x
k �.��=5Y�m�y�0�n�&y����P��!�8���Vv�k��u����уZ�Km�yz)�u.�{Ƈ����GW�?]�i�,���B[s�x�����fK74��1)k���ԔH�7\7
�-H�Q>�=��mM�BN�/�	��c"��}|n�����Ы��Ҳ�3�P�_��ŬS���X�
>����J`}Bv�	]������ߡe���&���$r7(�<�f�ᓷ^���5=���[)��K�v�,�9���Ϋ/gXEꖕ2/��Ҩ���'o�-��:���ę[��U��G��w�N5Sd6�ƴ�{~?+Bv�9?�TY�<PavL�TMt�E�_U��J i�B�o��p���G'W�����/Z7��g��z���2�p"�
{�U��d�/_��G*�)=N3;��Z)�vuKxIgw�V��յIZ�r���������R�M��r�0`���'��<���'�y���l�ֲ
M~�C1BZ�R��벾��+ٻQ�lMӍ?D����LL5L���vY��.���g��ߧ*�Z���༅�����'e�>Yuu����E���xH���NU���Y׉�ƫ{'��x�.�� _UW�	��a۸�c�0c�+�nb�v��@.i�;M&���9xgb����(#k�d���CQs�'C:���ߚ�'䤐����@�O�u����&���;n�N6Ov�.h�������L�L�'S����&��^��A���UGȳߦi��En�����5��	2\�7\��)���C���%l��Ǟ�@~���>�ۇ�PK   �KX�C��z �� /   images/cf548ed8-d697-4c12-ab8c-ecc45c0ca7dc.png|�eXU]��(��.�N�A@6�JH7�H�t�:)���n��ݍ�t7�������9׹���{�k�1�q�s-B^�(����@��T�Ah�ʆu\��q ���\ ��<����=�H�*���h��a������v�u13u2�u|c��+IAL�S���g�v��/y��_��y����PQ>~�'U�]zu��i���;�#ߐ�ʂ��!�Y�Os%�l|���1�Џ�(��7���>�So.S\N۽����o�KJ����?�H1���-9����OJ��v��^JR�e3��P��P[$�d��Պ5�F*�� <"@U��H}��:�d��E��XPF���?aF#���^6��1T�b�Z�����y���!3w��+��B|������-�S���E'$�p�մ��չ32JKO������ק���Ӭ���
���g��4t�Ɋ��c���ț���		Q�����)faem�WE��
n��������a���w�*�Ǐ�?�W��:��,/���Ζ��uH��&/��`Н�<�igZ(~�a���������ז�+��N�3w��񰱱�������������T���E}��s��s�!k4��Kɻ��<��-�0K����[j�}�5�|�,?Y��M���BLE�Ar�zqq��G^>�O���r��`�1�Du=���c��kku�Fs�������-�'~x��:��7��nnn�Z���A����!%6�	IW\O���]�}^�����Y�ҤrO15uHI	�B~F���<L_�[���xa�J��l�D}Û�����|�tbﻻ��m�AGg��������Ȏ�q�e�������޿G�DV�|�k�F��{z����=��͵�����Zh��r���Ar�ěN�]I+����}{;LSS��Z������������W����^�U��K&�	����<kk��^�1��@|&��pHk�3���O��o�$�����wc����-��Lw���+*4�ꛚ�6FsI��x)5��2����y�����DddyF�ppq�45?>����O�3���?Y"=/�{����Gܳ���c�oF���w��O���^]�mh�����>���"�̌r�g��9��f66����:cE�w
������2k��u?�
4��H��#Tpk��EͶ����V~�y�$��8�ٚR���
k��w��X��|��=
J���Bwf����2�?:���5�$}�^ԣS	OĘ�G��@�̎ w����ETT��_��質��M���T?I�Y>Ub*Wa=�(\}�� _el����$�?|�*e>��R�ڞB5�ۙ��p��^P5���_�P��E�^�/1����/��U�M�	0FA������n�����SO/�Ʒ���Ab�X߯@�=1�wJ'CLJ"��Xz�>�Gx ܡI�ſ�T��EC��k��x����6Z�)D�6!��!.(����̧H���D�b;;������mc;��)�}�|����8	7�ްs?�(��?����#'�V�B���g�8c���͚��j-x(:�fP�Ү�^:�"�D�:j����ڽ��ڃ)d��`�0K���̧��[��v��y�2D)���|ԓpE���8��D��;,���Ѱ��g�1�4���'J�1br"\`�^��@�qMe���%2�g�=������QpZ�(pY��P����Hg1�������xvp0<ङa+�Я�d�Ǡ#���v����IU������2A��t'�_���{�QZL!3���/G�
���yDP0����G�nL��b�O�`�=gޗ�H3d�Nw�X�1���$먧q ���$�NrW�F��z�+rٌ�?5j�9���g�A�X�P!�k^h�[��'��)#D��z'5y:|��J-	����h�~y9����x���(L�U$���#�ƖUW�����m*�ʧ !%���ʰ�M�W��c�������C�ٳ2�������n�T�&�R�heL|f��D��n�<�I���6Dh�����y_��Y$���V
��� ĵ0�����gX1�%[sc���y�Ijd���H�PT�9����V�&�ԧXG�{���b����8Q,��=N�Yd1"�G��EE�N��۬�n]��0���F���b����S�3M\ ��&�u}��b��ID�2�����%�}%ݜa���OX��l����QJ~��F[�Ӊ;�o��+�aF�c9�QA!����P�'C�j@�h5��S�0���D3�;��������y��7���cd��%�������p�q��׷��1,�2Oy檅��������ҧ2KF���I-AI2�+��E^!�xiiic��\M�+Z���,�� ��e�D�>/�|e�S�w)I�Y.p�i����cOϚ��4( �+8�"=���x�����eG�Y,��(R���y���EP����w��D�NBL��ht�ۅ_�����'�={FDB��œ�칒��Vm����� �۶N�������YY�Yw)�h]�����C��J�ݖ��_���>�Wt888���y��K[[��>G/��6��5�5^8uV��KN^�L^���o�.�/+��8��Y��
j�I�n!��\��\?O�/���3^~�hp :�7��>^�����s�T	�+A�4]l�~1�4Ӷ����V�Jb�EN���b��P_,�>��(		�2
-%�p�~�4�$:�)��x���#������B��-��pc��,��	2�**Ex��p߲�B�x/C
�ٯE�՝@�S�y�́o��Q6z����|EY4��A�uC1h�m�B�����������p�A�(���w
�SO��J)c�߅��*:�1�Ͷ�f;0uq�I:�2�5T���'�� (+�t�ĉ���� ��`��[���2yF�(���Ѐ�(K�E
�N�$�������DǋJq�&B[�A�z�tk༌�������`�S�s��m��%��ĸK��ъ��5�[�����;����1?��P~hs�y�I7�xQ'�%�Cݿ��*>�:M$�裝c��?��������ϡ���BM%��_��m�>X�� 
/�D�����%�Ei�=|�x ���1Q�9!#-u]p|�Ϳ�>E����f.�B-s�R��A>Ә0F�F�P�s3C��]�%�F�z�:��&���Wѵ�hjZ�%��8�W=Zi�5���Az���99y�T/��+�c�Լ���ׯ����w0Hˣa�p�����aڇ]5ޣ���s`�j�I
��m�ыLK��Q8��c��]
}G4�Z�J�*,���5������4\�B[�
��N���ڂ����k�����`��c�.�/ɐ8����E������3�F[w|O�x�`-�B�4o����&�S�w�u#N��v&l��ޣV�][��g���~�JW*��"�c>˔駄�����?�<�J
��������@fe:'�L���8��?�7pI�n��-&�3gøT端���זR"�]��}�f���X�!h�q@�1�Uv�h�~d��Pl�1���>���ī��P�b��F(��̙V��CD��Nh�q!ΐx�諯}l[��n{�{�c\
*m昦m�;E���(�'-w���$�����"N��F�$��	������\g�Ej�]�!&ѡS��Q�/D����2	�;O��m��BPM� ��/*"[�"2��^R)��tJ��7���C��A�wj�%%>�e��	|���_`�!T]?Ψt�T�*4Ę��h�:C6XY�ԧ�Vi�b�����ɠ!�g�d�V�=8��j�|	}��F�uZ�c��J)km��C�Wկ�ape��t�)��4>��>!��8��K뼡n!b�$$�s�[|lu����� �HD���F.g����R%Q	u�����'@�����1y!ϟFϿۿV�<����R"t���A\��M�yh͡8"���g��0RH��o������zdzqd���!6� ���d��-U�+�c[��~�:��=�w�MM%j_�f�H��~��g^cJ�>������Q��}���i�\�3V�9񉆬�N���:~C��a����|>�:D��~2����P���JS��ڪ;*��p���n��<������B�!k*���*YF��v�}b�=�Dj��	�#W��"`��7�-X�l���>P���&1�.p�T���AV�y��a�?Ň�gv��}�mu��/�ܾ��L�2Ě��+�b��� ��d��-U.�����ՂX�,�h��4����,PCo��m�S���mW~�%7γ���gB�Zޕ�?��1yG��zc���5*��O�w��m����\M';�Y�~
g^����	��|Nf�㙽�M[ٚ���Z=�E�H���CM�ܛÊM�s����c4Ŗ��?..����z���ʦ@���P�=�� ��	NG��,��a��_�a��٤K�0�h�*�Ϝ�j�Ԉ���U���S�a%|��H��NO�����'BY/� �����{Ľm�癟ڋ?si�60�:��~�Z�b����j���#� !��<�,d�ǽo�=~�q�eμ�?˾߉��dK����M3r�����^jX߄�hBhV�es�����l!D�K\_�r޿�E��0QL/E�c9��=89�h�F�b:���V�H�y�:u��2�f�o�7$B�=ŉ9��{lh��e��RD�v����%����/�}BC��-Nl#�,G�l9�Q�܆��!ۤ����2߲G~�7��{	T�Z0z��ʒ�x���1�x�w�D(+�_�eV� �ǝ$`�P���*����U�C>�����V����S;I�Ho~A���h�i�"V{�TA���GM;kzq_�E�8N�PF��C��6�Rez���G�C'�W[[���1��#%�GMMM&!!r-�y)���#vn�cW�$		�x>�S�1�� /[%����W��L���xrv�2���^��M]v�YGG��۟�/��$Iz�dff���j־�q�GΙ��
��'�9���
Kkz�s�8/�b�������>���տ�`T0CVsǓNr|�f���i8�>sB�n��ҳ �A���_g��)쮟�̈�oS{Kcacc��|�Cޞ��x2�gc8�����y�e?Ӄ�EFr�^���%��UuwVI��������/����"�|}3$�lhYZCHٜ�֔���<6����YxC��8LDK��D6���,�%:ZMO/[��.�����q�������(*&���˽����������s,�ZAC*8�\Vy���ǩ����5n����������DjN�ӧO������G���.��//�S1���=�p�TAU��s���X�h��Q_�@4�1�@�k��I::Uq��CD��,Ы�V�V����;�������+��{/X�%g?J���a$SH�(��t�m�J���P��HO���c�
�f�a�v���JĎ?5���*�roޔMDd$�/x����_����a���h�Ap
�e�����Q����bfO{OO��W���T<i�;�������(�&��#��fR�����Ғ=�g?F�ӌī"�DE�K�o�3�#0`�~4o�#fໝ�$B3��Z9<�(��=��Ys�dd�G���)sS�	sR�z癆���7�уD�]m߷���~2��)V�m��H$]GEv� _.S���O���D9�������W���YƢ��	0�x�'S�(ez���j��ב+�m�U��*-+���U������g��·����4��ލ���p�r���l�������Hd�G9ly(m����Q9��1�p���e���sh8mLeS���Y|*��
�Oq�x�߷��E��u^Zie�p�W��S铁E�TS*�����_�	�YG�����΅�5h���'�C�������;�%Sv�Ј�̳z6z��*:��JON�������R��vh��F������k�ږe���P�C�(��E���L���.��a����M��w��ձ.����d���h�p��(���N_D���*!!o��0�&DV�9؏�Ã�������t�9=��Q�� ��2��k����r�W0�#o�x�g� +%-'��ٙ7#jw���\�^�6��߿I�A�z�r	�z�x�|a��M�l]l�a��9��f�zk��eU��}�'����+Vݜ�[5Ե�ɕ$��		�e�M VyX����l�:��˽	@���|^��A��ΖĪuTQ���
Ł��Ρt�d�է�nD)�53���������/�B;�n�8�er8Y�̄�Ȥ�G��41
��5oVCg��Q[IY�vrkRH6mp�T�������g�d�wò������Z8�nz�M5�U�c6�Nٰ��q�]�*Z{S�H�v���Z�/��O�d:~ja���8�G�<�jd&�ci�NI��h�B7�1���>�G�򪭆���W��P�bc���3���J4�����D�
�5+���Rk�|[��KL`ٟ��dkB��:���M�y�N��%S6�>�u�<ݧ�����A> �Q�r�e
>H���7�N�n��������-�A4��Yˏ�"XP͸Zd!��3fb���u1�
0�}�c�d�H�p��u׏���xo��./��	^�M3cY�;;1=*�#{l8�������WZz,N.�cl�O���'�͓�V��[�:�^B��X�x\<[��{i�)u�\��;��y|l���a�XA�Ƿt�f1�(�_������~���Z�GVL��π-T�)w��U�*{�yz�i���//Eg���}�k�dMY�Q���*��7I���$)�X��:�"h�����2�o�n3�"�ޜz�>k�{,}Ьڴ~����	��B��n���$Ì�Jƶr������5��t�/��Ma�/�rfsC�]��ة,>�r�{s�_N�����,���I4-R᥺����ڵ2=VM�4ք#�W0w������{>�_���
�x�O#åC��y"
��;G�y����j�8�c-PTga��������/(���~_%)�j�~���d¤��vbT�������EF0yyfnn<�u]�ݏ��i899�V>�01���3KK�P�Vڌ	����$�X^K01A?~�H���U�E��ԄEHH���ǧ��i��{L�Q}��������?��4�D�A5����3�%��͙<Y��\ZZ*��<:<L����/�10��V����ҽ23#&'�`y��M�OHw�����[,\\�d��^��~�7F�~��O�ӎ��8����ۙ��)�i���@e��·�����sƏ���s˔���Imh�-�ky�eff����w~u�
H%�JQ����ٙB��)���l�. �P�4��*���@|Z��ŭ�0Z���Rv!Z����&5N�����O�����O���C$��q���[�|A>�Z^YA.{�$--0�6�;N[�<�1�/�J��xA�_eg�+��B�0߀|P=����>�*��"*JU�0��{/^�x)Yq�OKc	�n�! x�?[�ܶ������k�c{���h���� "��� lȒ���J`VV�$$$/���Fs5:�����M��i�����E� �WR2����u�Ǭ�7� �#�#�F��$�f��*�/d`�vB��X�7mC���H�-8�(~/��44R�V�z�eSᒴ(�<U����1�&i��[����'��p:(c9
sQ��}5=4�ڥyq��L������<i�S;���I�  W��D�ݸc�ˍ�
�
N..�{Ϟ?�����쌲èɷ��x�����OLyS
>c��Y����`v>�O��52�:�Y��ן_�zջ����b�CFA1<��c=��|���]�׷�c!S.�����~���\���E��ͥ�
 �_{��=x��|���D+���[W�A�����ֻ�����?}�4�
Ro�������w!�X@�a��Hz[a���F�PrWd|�OWX�����f�F}���k���P��J�Z���mRg�r��/9���x�2'�v8�PPP\�ϝ����27��F�U㴄Z�W�����3 ��`����rGXhPo��&�?�=�MG�#���S��&oo��MA�KI%k>MW����aU�1Y���]�{�am�U~EE��Ձ$�OsY{!+�����<��B����V���r�WW__��z��c��V����=@fX���$$�Z�gd|��>P(on�,.:�� �0w^�ٓ�(�nLy��	���x�}�S�$��9�<&!�Cm�ap'�~W���m�...,FR�|y���"����J�Ao[�F�بL���ֶ��5f^�H�GJ@ ���X�}���қ�߭�HQ��A�_����_n��{���	jkLb�s@Q�Oчș���C�WP�Y�������V�v���Ҩ�+���\0�(���B��Ę�F9������v;�
 �$}�B�_���1�H7cm޿�[|�,GV*'�I���=�;�� �+�+��������h�sʄ�&���־d���c�Է�X|��J�nw��(��W� �CӍ>��.$켼Yҷ�潷xp��\9砍��Oi�Hz�����)�f��~J3����*�+D��0���*��lƯUI%���r�Pq�I��C�c��$f}̙�����HFLL,m��Y���Ç1q�z�O�nt�����=zvW�e�Ս�U@x��T���s�k��^�5tn�c�����@\
vDu%���t[��lmyZ2��n�����_z��eu"��gǛ#��ҭ�/��;�oD�WV�0+˩��"�pG���8&�M�6�83cbc�&K��%|	�# d|�q�+�R����RT�|�j��ښ��lާ�*z���G%���d�u\�u$�ɑHv,�<��/<��ə�3�k٤����a��jq�mw��;��[�@<�^��*{�2��|[�J���WWՂ跋F2�/�����O�^/4 ��\w�q�$�������CR���Z��ηGz`!2�-ѽ�SP��o�x��3@V����$���S�UX��O����~�:#g$-/�{j��S�x,b� �UC%I��$AOb�bcuu�u����n��;c�E�a�m�:ď��*�F�H�� ^� �H�J
ajz6�O��2�������?�~ۥ�/��V888D��B��{Mm������"�������|��e������?�si���<�3�4ֽO�C�V���
"��;����}+FFF<��X>�ۥ�[ �ܕ�0�F��}�+�0]n9?�d4�k�#Ta�����c���s�GPAW�Õ���d�5飫��_�(��Ɍ��S|����uZ i�k�������˥C�B����yˏ$���Sj3�Yn�%�i�E��#z�,�����r�1 �no8�հ�{l��ݻw_Z��d`���*Ը�s���`5��՟����f����2���k���v��
쓭��A�7Wgf`7���f�$�ջ�	��HMe�X�G�j_`nQ����C�Da|�.�F��ԏ.�]��?��Yx9^�gі�ȏ&������h�}{�/%���"P���h��gY�t�Cʦ��M���Jm,�2%�����|)�qT�D|��vln�"�X��&��ڂÊ �ӂ2"L+-&F������_ �9�h,Ws��(�m�Ҏ۸����u��B$��������<�}�;xû��d�_bO4���9�t߁�S='^��z}q$���6�@l5����ރGf�pY�K�E^ꢖ��YY���8��kb�vZzv��Q�F�zu^a�ɗ�3:q*( $�[q�\�SG6?��g�j5�2�}�瀊���������<�������B����VD/K����"9�b*���.�{I�c����F�q)ѱ)�JE���v��ʒ���`~�,V=���l�FB%<v�T�NȤ�?��D�F
#F�qZ�eg$�pD*)1��X��� ��:;�{�Fv�+�M��6G��Ϩ���"]ѥ baaa���SE��g�؋�=�F�!��6�%�(�#�t��pɊX���(��F����G9���i�b5]�f4d�|�E�e⾾�ؓ��|�O�xԏ�%���MYed'<�FB�N�L��mEKeE���d	bbbM�
6#Y��H#�����A 7�'�[Q����Z_A����� �B��d	���J{�*U�����$[%��� [�]���M���������M�����R�����'��t��X�j�TM�� i��{���8|q�n�E%d���|{�<F]i?���ֺ�/���[����
�FЊd��А�u�\�9�<��������y�+��U���g�������81WZ=v���T��|�Z���-`@�)Q���z�����niQ�
���T�/�]*��X��#O�Β�w�17E��&*�@i�yN���1���M��� �R/O�4 �ټ9[�oԁ��Β�T<=k����\�zoo��'�{.cO7x=���k,��M�1�u�Y�n��W U�DFJ*���Ӈ�T���qS^ �a�,���
.�f�:pԮ%�nM�C����S}��$�hl9��V��Ѐ��3vs:ٞ�x�����5K��ʊ\��=I�I�M�Ա��d�b!���B�n��n��:������?Nڗ�F#��"��=i�u�ptt4y�����8'��ۓ1�U��ocVf},z��eU���+e�	7�P�<`���{}Ga0`E^�Mp�	�����o�w*�3���cB�UF�Ÿ;8�v���ly����9�@r��Q
��(;�M��oLb�x�`Ttb"�-�S䫤Suˀ#���!�,���t�k:OHjD�9\v���1ȫ�Rhh(lK%��)���yM9 ��8AR�s��~�;�_�f��v����C�k��x�I�Al��}	P"7�4S�?�ӷh[X0�����.(z�KUM젲l&v=�7�'�x��P7���Υ�U�����L�|�x����?.���s+�Ȼ���Ks���Ms��a%�|����`&7#�����`%TcО�|k�8> W+?�`e�B(g�����Y�r\LLWk��۫���n������j��cS*k��� �QVg�9����2!ȅa��aK���ܗ���2�"3��������Tw
Y�v{{{��,uˠ�U�͙�,���ny�J��t@��Z/�`v�1�V��]��,M/����Tl�;H"� ua�@]��l����V� �-����U?9�����H���^`�a���"�$�~�����U��r��;^��<z��o2�1��p׉Yːr�C6(�=F�A��5��(TW!b>���#A�Ъ�0]_)`e�����x�k.j_A���-�~�֗&z�<�ٞo���#��^,wX���,�R������~a�F���{�ۖ��_6�$+��2)@lMSeY�r@��)�]�>�u �*+k�gg'����k�N�l���VS�YX�<����F�3d1Ns��ACCC���BV���}����D���1*���h�i�P�;�r��z������o;ee�x���7E>�Լ�sA���b载���M���(���]�W ���e*\�XXP?Iw5�exuuu �\�uu���j@�����4Y̌7.�1h�IKcA���Ix��O}���BZ$���5������OҼӫ?����e~,a@V�9QV��.�WW�o�ަ�pi�\̣a��4���I&.4����'�}�� 2�����l��3Œ�3�:yvd��2~��x;�P2::��ֆ7��S|���T����k�օ����V���#ȃ��ә4��9����>.n�ˀ��e7(-����d�R��g>�_�X�Dx@�(���˽���B��J)�S�g�4@�i�Є��܊����=�茻R�_z�x�j?SE����:K\��!ZI�@��%>��py�I�_Fg��2�p~�M��
��b���KeV���X���t���i?�-Wa��n\
n�sP�a��T�B��P몪�\��E(+)����Ңc�⫠˚�kKK4�����j�Ik|5H��u�4����Yb�G3T��Dn���рY��n�+�d0�-��6u��$`�-�fȟs�4{��q�����V����gۢoK����
}����7Vvv���������{�̞{^�ut�}o�G�Җ�I8�����A�z���o@�P��p�PSS�z�n$�{}��LdA�ƆӢ���yo��'ȭA>[���o#Ș����f'U��"�5^8��ʈ|�%�3%�mw��*T���kh8��R�eJ~���%�ׯ"���&�z{�$OF5 <��ބ�R>USW��.k�?�s~�����t��O����\��&��C"b�wb.k�`�[?����G��SJ'���I]��K���s+$�/����d}`I� �n��XOO�s�&D�$@z_��s0�˗�.�OLĀ���86GH���<�3VV��m
�";//E2b�܆�����t�ߥE�hkS�6]9@�]C�
f=q<e�Fu��b�Վ��I�N�<H���=����=�J9���T���Q�롵��o#gg���.�3c����y�s�r�]�����/6br�{�;%A�!���� �TGH[қ;H��c�*'/�2+�'C���Sp	qՓ�����YA��*����%T)�@i�ȵ�c��q��I�ˁD��BSHTq�f�yO4p4�*���"�$�X�~�o�+�kpW�J�*٤ZM+���w���ՙYn�kg"����=£��k<&٭]g0S�Y�p�x���!jn���p�����t�q��@d���vb�k�ɬc���[P,i,������qD�Fb����[�k	))z�b���z�j�x<�#��w??`��}���)|վvu)-�W�ӕ����	��Fx��YY��S�z/K�zj��\��JD�ԗ�����ි�J2�0\XQ�����.x5Yb�1Q���'С@�ִ=���%��e�;4�P��쭣���J�E|�*]8ٚ�R���e���W�F6�;
ڝ��N����[��d@������a���U�m��3J{��LQLP�H��B�>ۍ��w2�V}t����o#�����q �r�#��-��<|q223C�	����齆�$�����g>�9ֈ�f�����[l=��*с��U_�$�(2_�DfBږN����{
	�t���/$�.v����9�~P� ��z-Õ-�k�C_�㣕��Tυ�	�C�%	�?I���m�}~��=1c�7oU�?���R��o�7j��_�<�w	���`��E���ϣ�c�`A����h-�؄�WLN�NmĔ=MAs��%T��4�Iȁ�-5�$ʾ�����H���Cd� ��*'�]j�qr�$3g,{�R�5���X�O�5����|����|	se��!l��oc���򗧻s��䔾a���~zt�e����`�'�/dN���)"�����뛈c�Ǐ�F�㞏������LYg���.hz0[벾����ܼl?!!᫘�}�s���fQQ*@H��>��cU��u��.�����3R�p�ud�?�I�2�;�O��p_`��_߆�}d���8\7!���� �v�W�[.��|�&����Ԇ����K��_K&!��ďD5���G[�A��"O~��"&%e����t�D����%%5��p��0�C�cPPX馫x�
t$xma����)�:M�&6j��={�IsSN3!ȋj�bY��R��>��[q�� ���r�Wqy���qV�1������y�0z<)��1+xdf���Wj��H�N����x)^�0�,��U@L2@ ��	үW�E��lB4�UBh�l_��/�g��H�����C6��� ���,�����9F�J�{�Wk}�SF�-��U�o~+�#���C �|9]a��..���rl:���g\ZZ��qf5�;�Z�ݙ�N�؛.L�����&�o�cӻ�b>�׶>cO��fk~P!٪��	9(��v/@�
��]]|I��b_�S��>�?6����=��D�G�O!{���h��ځH���3�y{��s�>:OM˩ư���|��-�p� J�p^F�>ݶv�j���ﮨs���B �Mw�,��tgF����߫��㒿WW�	tṔ`�"kc�w�mh��Q�$,dbb��jB�[��@�]��ZT�T�1S�üW����B>���4��=&x�8o�|<㼂�Vx���x���u�f�SEEŒoA,�����/:�R7�n�[����>Oe�J")�� �P���l��k��9H �Da�d��!��~��?�NK	��"�ľs}w��Gޟ�6:P�Iy0|��f�ۮ*[n���#///<���E�v'�Qz>KA��u�"�4`vXXX-�s�?���X���o�����<��h-4h�P�9��N+*)�ֱ��C/%��x�zW˓��ޅ��BtpSD���n�OC��
�>�H�9�u�%.����U�����缼�pc���rs��XI}�S�xDqQ�������s�av�'��_�%~�ʎS�ِ[.�.&�'������hv���r=��٩an^n��ACZ`���P8��r�VO����[�����|�p_�L\J^݆j)�Y垊ѣk��������Xܪ̔L|��RU��̀�kij�pp(�����ڷ��/���?K���Z�;��å$#��c����<d�Ovߙ�2.AH����NUy:Sng��>I��pZY�T��#��v�>�Q!�\��1		8f�����v�c3��H�o@.�����F��]���.4�vHި�1�E�pW���l]�  y,������I&����&�)?� S���Wn�ᝋ^������g�4�C ���S����y���	�}~hOQ���������������B���{�6m럹@0�l�����k�d�ӐQR�zo��p� (�X���E�����6**���B>�#��_�ձ�/���W���g�L���u�Sj2���V��<�8D�<��uԨ��J����
�#OA.�l�t9�T�)��f�{�~�F�GnO�'˷;�Q�3OxZ�Eoq��h��g@p�S���Eu
8}`�=�P�^����C�
�# t������Hz��


aYe���R?��1K�n|��	�k�V�|��h�P<3�
pn�*�љ����	33�n�U���;����}�w�[��"Z���wr����	Z:�(%�x�MWه�
��S� �m_�YXX�Mvf��l�s�J*��XX0�Ҕ/la&\��@�=:��|���@�>+K�ۖv���D�t�w����3��:��j*U�ۨN��! �@�f���>tߝi�@B������ BF��ˆ�~�(��9ggg��W�F��'��_��!����bx���}ΪjZ��hi�.��(v�x������3��Me�OMM�%h�&���鯱���dUX=�����L�����שee�*�ҁ�����	�e
j���	�w����t`j[Q��ii�(iL����v��a.Pҿ��.#p���w����L��ȉoV�05uP1w�)����?ܶ��^�״�pK�ӊ�����s�����/\��7Y�߱�V�ud��V�as$���W����F���!h��2�fvlfv�f�Kx��Tf�aT�;/���lӱ>�����3~���4O
3n�/(��9J9
��7�gB[��
%��Q�q���P�;��x�Ļ���x,-/h%eF_��J߬>k8��I���?)P���ЩgVV9a!!�g�s���V�ޓ�׶�l+H(2�����,�m�Eߛn�*����0Y��:��!Ec�&&kS��".m��@3��'`����������.'o�zd������!�չ�h���]i-�88���66�f=���]s��W2�F'��X��
�H��q�F@�q�[���W���%D?�..�D(�m�_�qn�%H ������6�&a����VϬ���JA��Gto��k
�;aC�O�Ɔ�Z��h��]0�4�<�'�F�ܯϝf����l EJ�j�)A��*�WŠO6x�[)�¾?������@}jj������'3 x�=|�{�j5w��_�`s��m3���� ���y̨XZs��a�K��t�d{MO�i�ݚ!X��Ef��c//1a�I���Í>S�����su�HHI� ��<��9����)*B���O�d�;&vߞd���2C>&�)���{vW<-=��y�I�(�64�%���˯EӀ5B�А���X���O~ڡ��^��&d� Nu��#�8��VV̒ny^hk�'A86�0�`��`%�YT��ښsܿ9�ё�
"y�r��`R��QP�T���?H��k���鏹d�r�m�`{��>;�U[��s��9��y:���}G���:m��az7C!��;?�,;��f{R ї�3P�
�~�u��N
ŷ���	#phO�tR�K�1�Y�D��#����tN�����+!f{%��.L'�@k����Lz�ڠ-���~1���=$��$%/;�W��y@�T���B��>g�o~c���M�w��d�qf�X?�!�,�=��?x�&K�]�ܘW!��:�Y��x;����b����Xv�%mxX]�s��Ǡ*|�7A�V�������(235f���� ׋����%]��	Y�ga��.*��4y�����&���n��w�4�����j4����~ ��Ӈ�JKK���9v���<8�X}^xGBV��iNUܪ�U�����������}�j(-��6Z�G��R+�%�{r��F��Z�;c:&n�XY.�����ic���*D��������VV�Ib~W�z^��~E)�ǂ��������4M�[퉷����Pz0M>l�(AZ�*;�d��~�{Y���&�_n�!_����e���[��D�c�fll��v,=��d	X�`����o�<���t[*�1d���Y{��R� }���%�ďUY]�踸'��ȷ��o�AZ\
n������� �ji�=RR������n�.�C�S@D��DD��Ni��.�����~���Aϳq��̼��ϼ3{�6����J��E��m�,Q�绯fN=@G�hjj�(�����p�'-1nɀ����f������(~B̍��U��;�Z\�̙:�]��mi��,;Z�Gc�Q�7(�g^Q
�ys�gy�]#ystSV0���7�C�9I�����·*�%slv*��g>��Dت������6�!�;NUO/2�E�y�яru�vp��T>3\sl�����4��r�a4+�LQ�B-yeeL��CɁT�a&����$^;bh.�+��Ԩ�RE���i��HH���/	�p�Wcĺ���=L�ؑ -�Ï;LT��O\<��E~y##��
�TmflRR�XS0LS%���ښ�@�2I�R��\ӵ�JO�V˕)jV���,��gX͍�7I�ɩr8if�ύ�/���gfw�fppqq-0;###���.t����?��'H����/��#Y�Qb?߰9SYh�U�Z걕�H����qk��v�����nv �z��������4*�^*(t�dK�[�W����>�Js^{�Ā���E����ԯh�C ��g�A�|�qh2��Z]��*��^����L�E}��q1S ^+N hu�TZ��4���S���3�'/�<����C�YdM�ڠ���a��ݭ�:���GMJY.���6V9��i��e�m��FdT��F�����w՛)ʅ�]���\^�]�n �@UQ����R�	`�W��ݑ ����cbD��jjR�##�f\�����TU���v�A����RΜ������U��>����\����t	��s�Y���k�s 4t+,P�N7A&{5��Cm;���n����H���-ׯ_���۳M�����W���i�l�Xu/3K��s%�NA+
�_���<�W����Z�]���ϯ�����U��<��Bk;�\��a�	�EY��[n:�����~�K5��rL�="c����7P��Ƿo055yy�X`��G@�wnO^?-�0�H/7�C��B��6m��J'���Նn�k���Ȗk��P7�W���G�����7�'&z���ǡ��rXl�,o@G��O��yO��CK����k:0p��[�w���

��}u[�~����} �����oL\JNI���u?T9ԋx�Jlll��A������6�v�Q4�R^`��JK#�
���:����;�{_�w(�(�����^��Epuu��ꉡ�q�}���c�c&LX���P	;�)@K� ���9���,l��Gd��B[P��a��u�ٿ��JHH@S�#%�|3Y��@�_���S7W�՗��cg�R��;99j�A���E����)�V��)�J�Zs��/۠�"��T!�S���v5^��	�Dv[�kB�����g����I!��ܹ�$�$� T�'8�X;��t�|���s����c�]�?�����s�8Z����'��=ʇr���'<��S�'qe��ۆ��^��0�����L���rb!�F?�Ǟ��h��A�=R!���6������?~�QTĀG@ i<8����,���&~NN6>>b�r8�����y-F?�P��d_�z]�����=`h)Yَ�E
�tLB6�F秠w�GF��ϖ76���9J��2B���m��$���oJy5AoAd���&���ЏD�q�V'��?�G�"X�N���Ԙt��}������g�:�V$��=��8 ��/��|��?���'K���}��}�+`� �].yl&�8x����#dM�M�Ͻ��eL�>>�^�%�v<� Ԕ��򦶇�������5+99����^��v����%E�֣�o:�"�:u42pҽ=��K+<2	�F����&wP�1����N�?G���o�����o:�`Np� �����C�����щ/���c/��'+���~��ĩ�R�al���U�r��=����~���'\�ǡ�Y���/q��v;?�y��Ӿ�o;>��g1��[(%,%���N���٩�H������|���N!zuۙ4��DI���~>=b�3e�Q��Z����'ay����V�E���N�܇$+:�[�R���;K������P��ow����f������E����Oel�Ҩ�q���x�=�X�#���?|g9��eF��}�����q�^��mh.��3�U��K�?��v{]��dD�m�/�.N{�F���� ��n��T����>�o��>g���5U������C�L��/��s8��f�Dc�Vr��3�����1[A֜��n�#Ƀ���>�s{�_i�o�yld��WE_�=���G��YŪ%�h�o~VK�a{���'!�p��sX�an$�M��q�|>��}�`v�z���HC����#t����Uэ�{�_D�k�Lgu����n�q��z���?<u�+�8�~J��� ��M�W}�x��T�Y̖-�W�$�C��级's�zt5AEO����f��4!^6b:6�\�HS�(��Uv5Fz>mQc~��}�+j�y����C:%����_;�EL/�l(Nt_�X3���[2��(Di�	�%���	���nj�c��Q�kͻ~�y�1��� {����4�'���g�ft�8�&V~XiZg&Gъgq��Ͱ�SN���N"���{��X�m�ׯ7�3�)"6�D�����9&o�ꅺ�!��2�<�΍�@$|�>ͅ������4��~��'o,�E&BZ�'Ǳ��2J�i6���#��>ޢ��b|���ll�{��)�.��>��h6%������Ǌ.�9�.hx3�x<{�^J'or}�j�R��Vr4�}���c�Y	n�#ƭ�36��G�LGD��@��U���2~��ab��j�<���gI�k�ҍpp��}ɹfO���+��D���;ׁ�jb$���.}?�xqխ/B|q8q�q]�u? �곂����[�G-I�x"�OlΞd����R�8 �CA�
�{
d�t�;�ES����1 ���/g��#�|&��̰aǅ�c���f��2�����]�Z}�ݮ�c�AP,PEL{;�h>��[fΩ�l��e�Z����m�I��3��J��� ��->� ~��<uα��S����r�z�7����|b�U��>�����8�]��)��]��[&V{���Cn���tnW����3j$�!b�Dy�ށ��y����^J��p�N_�'9�W_F�AW���t9�ɊҢ�/�i#�Cy���A���ݔa���x�vq�����b���_�G�����vh�A�f��'\�}�[="T]�h��78�Ȝ��H㺛�F�)B�"|��>��y,�M��}py���1��4�����I�[Ej� 8�`r{���s������o��o�/̳m^\ʲ̚l���L�vWd�v��<��1,���kx���\��o��O�뮅*�R�[F��c����ulݩՋP�JҢ�(�ώR�=��wML%,�푁_�.�SHj�M-�!�w��M�q[X:s�Fi-�E]�P����32n)�z�X��Yy��P�:������ђ{L�$��DSF"1�~pK$�݊#���u>ҏrr?o���b�v�*�_�!zd�Ԍ��lU���>'�]%���`}������p�5!DX��������_����"�~�� v��d�md�F�U_�L������'�F`��_��H03�YԻÁWb����R�N����a�$��w�/�&�y�7Q"�.TT��T�	�mjac�>��[ͷ,U�?�s�iy�����@#�)MA���y_B>��w���ѝ&�+������k{��[x�G$��!���uvKy��l|�H�����QÈ'vy�Sz���X�i�s��ck�&;V�iH��^h�˫E�x�÷����J�%��bonP]����/���H��]�ݓ<�}��L��8�_���&�	��!���Y*���x3)�O}u70i9��[�`B��Ox]3��S+1���,,�W���K���'f�'z�N��;�����o�ʜ80jzt�0vط�U����!!��X���^����ş����>�~��,�����w��"B����m���?���2���u��u��4;x���h��+݌�YOc%�;��OSI�x�?}�6�G�2�L/�O�s�>��uu���]�a��n�}pt����P>��K?l�Ai�f�u�bL��2XLۇ�9�9�a��>��c�y��-wʤBN�o�1�0u�c�'�&?���1_H��;�xC"��8ߏ�7h8�'���o���a6o-���Y� �=n���Xk��B��qz��V{ݫ�������;��t�e�T���*B�����?xT��D"����s�s���Xv ��iF�CW-`ֿCҿVnI5H4��յՂ��c"5Y�=�r��|�x�Je��T)�t�T1&�k#vw:���:�s���f�zs{w�/V4u��r���s��Z�a4G��
���S�9\_L�����b�?����C�wg*q�����7�?��ľX�6m��k��S �Dn�(�	��g���J��qI8}�q#�)R��t['�5�Q��m���
"�\�6�r��~�NF��
�-��AL��{꥙� �K�wѧ4q8����"�iC$Ǚ%juY�>)))#����}����qr���@r|�����!���4���r��b��g�3Hag����	�*��ғ�bC�;g^I���GS[�jjjm�{�:�O�+g>�<�H��'��~'C�䭭}��w<W
UHHK����.H:���44Sǡlmm]&E~:�����M�4!wL!�ddg�������$Á� ��~jèU'� �:�G`���	2��O�>9M	�*����2��ax��~��x����M�8kܓP(y����p1m�7"FM��G���.3�����-���ߢ���,Mf�fG4f�rߛĴ�����)���͆�/x>F@@�����\����.,|<[� ����������
%K�(K���<0������ޟj`VωIH���:��7�ӭw��Ѹ/�:G�*���rs��%�ɰ���z�!L�qm}}�z�޸��K˙�D�������KJ�à�sB
�=vQ��J��р�E�3/��Y٣ᘏ���3����r�-�O����Ώ�kϗ��P�(�Lj��υ.F�b����yk���A�k�뙚U���S����b�����[Q�!ZA���G������R�@��3�_�� �1�9�ʓu��Ņ��&�uV�-3�D.��v�́t��(��ֵ?���g��_�4¼H#����w�:Ӎ����rrs���B%t\�Evvv����떑���RH�s�hy�=Nl�����2B���UW�p\䑢�ڵ�����}N���a�^R

	eO��W�]w6������=�p�|/��^�lC�(��B{��U�R������K )*���.kM��l?���XS���A��--d��$T��<V���F�-��bk�=hK|#|>mn�,��v�'�/D��qoo��lR?{j�ܴ*�trrJ;���nց�RhZcO��%l�l��Ĥ�vvx��ȕ ݐ6m}}=��'��-�����'�B"[���O�|d�����3�oǖ����߿�G�|���u;���KIK/���w���͹/��b�e����K�V@�k��8�p����l�7&,8�H�$c
㺂Ȓ n�����|o��]������ajvv��s�/l����|�)<���L��Z6�Mj�h�3R홱%+���G���q�%ڏ�R��<A���~�:\���Z��۷��P��2��VFa�z;Y	пk��>^�:��Y����W�!I^��������GR��'cq4��]OuLLL���<O�@�kM�0��a�aa�|�g�5��ϒ#��h/���D����)S?==��i��~>��ګ����=]�ǝȂ�r8CZG'q�*Vq����G}���A�6z��Ϗ�[`�+Ɉ��7}��������Gs8Y��JI��!Ï�����X�IV�Q��ܴF���لN�YZ�$�-�ʅ]���e����C��I�x��.��UzV"�'�Dn!L��YnO@�����ev&%�8����rR~�����V��ZmE�BT��w��kt��cS\�)����, w������L���G��ۯ��M������>�R�I�����q�>UUq��<�۝.G��c��TB	����B�k��������8[�\}_�rI�2v��뫨`�{��=�pq�}�?xh7+w�����4ɟ�o����������&f`:@^����+|dk:���x�p��wf�8�V$2Z\T��:�����٨�ze��PS����ٴ�������%�tpٿB����۬��
	�^�6�l����3`M�Y����*vq`��˫���g4^�M����1
=�p��I���������cf�@#�g�6�<�O� �O �G���P�p����@B���9�\�e�5��Ԕ8ʵ���.lD[�7�;�N�5w��}Gy H��J�p�@�]@l���(뱶�>MV�!pF����V��?���(	n��)�c2�����͒���o��{|&Y����/�bQ\������	�Qg�h�d� � B���F�ELǾ����y�JE+�N���&Q�WBu������ם����?@(�p'� |�C�oOF�L���j|�av� ��=�#�o(P��4#}oΏȐ��\�t�h����$ )heǞ�!-R�R��HK�'�&�F3�����pO�������~��G�
�PP��'�p����5�z|RD�y�B�2��0��f����H1���������BB���	�q�$��/w��O��O����Q�D�-(�@U2�kkhh��,,�%u�@��'�d��i�2h�|>. +[�5!|,�($Ю���pXЦ�!��!t7�����t������ j:�T�v���%��>I4�Sjd,Ԗͩr}�h�h�35��$��'o3zޖ�T�����&�<)�j�L
ȋ>�΄3yɭ�#-�΍��<��(��$B�����i6Ixm��x��F��D�+�hGA��dX,�c9@�sQ���}i�=.3������*#��>�mؾ�g�O�=$�HȂ2��.�Ӌ���V86B��`�C���}��s<W@� :�V�N�Zm߃�$71���� j�D�8ߝM����WWWcGuI<'�p�f��ύt���/��-�� >��L]hT�2�-/	�^"^���n��Dϩ:u�ҳ�Ca?t�p9=?�O�X	7'�#�����CCMM����Q�vp@�������U� ����geg?z�䉣�5��J�a�@�x 9��LP<>�4� Zr<�Ģ���3�R��1Hq�����q4DDDKy�a�T���ttti�}������			���k�0���&o�ݯ:\T�H}kC�g���ĸ�@�Odh���4���qz�+gF���]���G��:/��2�蕼�y��B�	V�0(˅4���Ẋ��������`df^ٽ�}������jh�e9����*���?�|>*''���yBKg9�!c���(��h�;�c�~�����i[ޯo�E��"##�0�n_.����R�u �q�E8�z���Ȯ�t8������Y�)�����8&I�%<
rӑ��� �Z�}Q��	�ם���_P�b�|�kcVWW� 1����vO�NL �`�oi��;כ��.;�C�
�92���o����,���l}[��+��
��Z�9��N�8�����w8�,p�����{@��W��R)��9���0�Y��CB���G��@�S��,��;½�|fVNę�0�{� �i|+d�����yFF�V,�KɁ���0h6���L��g�?���>v���|$���.���KG��WE����X��Jȧ��		e!�S �%G{�Tp�ȿ��oR9�Uϝ���C^�b��QPdfC���!�:�t��ccc�n��ݙJH]��l(��ՉS��#�Cawޞ?]�A�-q�]t����b�o����.vgK��
O@�[]�t�����IB��)�71�2��Q�lUJjj��Q-�t��(�Y��E]߽ˮ�M�-��&#�q~�O�.+H�0`ٜ��2�P�n`^-7��$;U��ij�b�kA���Uk���X��6�p�h��ugF|�Ξ&&T0R�6B��ǂ���F�/@���߷���b�x�^YY���1]�o�h�`�d�6��(����c���NЁ#�����_��d8��B������S�]�ؔA���Yx�����		]�P��<� �q��L�;���J]�%4���ݠ��+�QP`5�D��D����? 
�������e}�WB�����g�^�ܠ��̞���iU�n�Gm�)� �(�ˤ9���'//��MF��.+�$Ez0�5V�@��灈�
�GIIMU��zC%�+̜��a1gS'�+���i(��?4!�q�� d!�CJ///~�R�����~�����������S��;��������H�l���{tt�ʜ 7������7n'	�舸�$@zi"�_&�N��㣯t����}�\�a<�*#�j�� X6хW���V*U�4� Ã��CNxYXX<_����AaceuHD�M݆b��\O
�����c/[+4/��ϲr���3�� ��|��Ir�j�&HG)0v��s[h�aNNP���s�ǫi�і#��4ff4�M888xxi� :s�Y$JnS$���ÓV��Յ��gi`@
�����	����l����r"d@*�=���@9� Q������H���W\[��l9�~����@>w�G��_456�S���0�ɡ�>���ɁA���٘>���r�&z3���E��`l�C�o��tMV�߇{����O����lQT��"m�vb��k�M��Z1���(��`c^��O�)I��x{{h��L���b^��8�!���򧤤�F�"&���S\__�cEH%%m�
�|l��������s���BE6����Q�޷��� GĊl��5@������9��Ȧ���TⰢ�;cK̍V�oʙ?��K��e�6 ��5�j= eb��kg� E���&��2~*DDH�		�|0t"�А��5џ�M_@��F6�z�����		+i�1:L�<��|--ݠe[�Y����݊����������?ha�Y�V� G���U@9"d@m����D��C�߶�\O�xސ,ǈO�]()�-��G�2�lE[V�gw�T!��/Y��z�{���G��CMO�f��F>�g�� 7H��贮+�Ȅ�8�s9.I([r`D缭փ��s�؏� m���ưe�c8�j ������NO뺡󂬗;���	��́z�['X*""��g�V�7 �ĥ���lT.�?�4{ LPPf���\�CҴnJ!m\\�n�6���ϛ}�[��n��!�15�6k�e�"M�_.~�, ě���+3ib�gL��N�aPN���7#Q23�*2���v'-ɭW����R��ʦ�&�v5��@�q �߂DfZ�7:9�����^���_�ek�f��5C��ԂD%���?Pn�5���I�e����#�b��qR��*��}�ǂ	�8�&�k���LCO�:[�ًJ\�ޡ��������U?�@ A'd�[�;�z[�n�۱�
B^�E��%
��$������ߋ����F���h�&����mu�7�WA���ϟ?S��z���b�V���cu�Y4 6����>m�a(-�ub�E��x\�'&&t+�<!����7�J�[wHቒQ�L ?�W���׵<Ϩ��`�R�$'�z:����B,�ᘵ�':::�Ga�|�������Ǟ��v���ms�5�����~̴�*��5�C�0�􆇃�Ӏܣ����d��S�]�)DIsϕ�^ԉDh�T�r��(==}�����Z��d�8%Q-}�vq�X�B���}��^@l�xğ K@�����BLi}��Cy�֫&��Wkx�b]ƌ1������@���R��w��d���W�64���焄�y:n�'41�}��r@5`��0���eCV�:g5g����ޟXɅ�Tgh8������G82*J6���ƦX�o�@��0_�tk,�q+�.�^Fc"%E愕_,��_���[\�fr,�ꕜE�z���7'����!�E���	q�7���t�48??����d��\�6�Y�	�����UUU�n4�
���񥅕� L���N%$|\�-����T�k[��7ȞQ�����ς��6!p�p_%�in&�$;.N�����MR�i�U�&n��"��N��]��|d�:9��!Z�k������ݻw�"��i��B����w�-� S�?Q���k��k�`E�]Gs�����F��dI@�bb���<���nv��%����n �������v��'��f���?��[�d��+g���:e���E��޾��Y��pp(�)�.>�������e`�Ԙ773���O|����m��W���B�:#>�z%2RR���O�=�l�E$���o����G�Ѥ��:�͎���0�o�Ɵ*I{�:�m�+�_�psts �V�+<k{�c����lk�g���C�L���^�ax���o�		�N\E��߿c0'DF�D�5___�,�� �r��_I;�^�H�����YUU�E�Qb>˯�wY��&����$���f���8�3��K_׾8W�w�v1TpG*��!?.������~>�_�s�Ż?\|���>H_P��{)�9���,,�~����wa�С.�<r��<l	��@� (0 ���1驱����=�hF�|u�]{nb�ɹe�V+�
��Y����6+n���[�pL�y�Jf{k��qXu�N���q�\|�V�<�˗/9�0 ���݄`;��_�� ���r�o���b��K��������b~�vvv ؄�S�[X���� Ϙ�+����o&0�(�Wf� -~��-��Hbr���4�ػ���x��*��d�#o;�a �Bs\ #�j�uk�, �����& �|RrUИ�FzN��0(��, ̍x��T�YQ]f�b��QS��F(��Ҕ7��g-8����0Ã��@3�6fm$9%(r��մ��݉X���֪xF:��`5�+��N��:
����_' ��WPP��{qg�ޅ���B�?��'F�L��Ё����j��X $�P�Ѯ�B�Й�*þ���������頳WKm�܄����O��f��T�#�I���n@�R32�װb
s�^G�����薫3y���i�"�J'�H���O��_�V^OTt�8��b�����o�@Tg�T@⚳@���*�xxe��]��E����%��O��cc��!�N!A� �CU%�?ϴ�%�CǷ�����=1�KMJ0�C�?U�Ry�Y��+�f�%���֏�� H���A�^�ϭ�L&@��̰���m���d�� 9P���C�l��[���ٝ%�S<}*�zM�l̷��ͭ�#k|�����u��_���666��+��fs<W���/��c
�˛��>������d�%��g6�~�~^S��(����@i)�:��vp`'&&��&$#�o̬���z��Q;d2��o+n�o��=��>���I��}�2�g�**ßk��#�������ʏ����ӧ���]��؈P�-]r�`�L�O �P�ũ;�_��2��������}H��N�%����(S ��{���~
���A��ҲhN�ҌA�L�|���8���hy��S0Y�Z��`o_�[dH,��q�YW��uE�����&����>/n%]����jf�&���x}������:.�f��oѿ����R�ZG}�3K�ү�4�'������ܩ�0� ���z_8��+���U��x���˴y���`o�u�O�b�&Z�Ķ·�W0ld*�q�zT����x�k�b�{P����j����8�j�!P|��q�=TXf���rA��*��p�i����g4�Z9gK����&Wi��`���&4�H�g�F�/�k@�m�	~B%�4bb=1�?��B~�i��m�]5|����\}�* �ibz,Z*b����E����뇱����憆��M�bI�Q���C.%7	�^"�q�����ђ|�g�]�P+�oS���������IO���L��3�����)�JF���U����#/G�xI���\L-���䎮�i7O�jFH�0�#8��PᆞO���Ѧ�;�R����_Fk�rW�=����E ��D��h0�t���ý������7�E��<�_��:	��t-F�>7C�m�Z��jA�;���R�L�cT�����w64ד �6ѭPԘT���988c*^^m�B(�ʓ�#M��"s�Q�:�ڃ�m+�n��ł��k���ݔ��A�y���e&!%�S?0��WX�R_�il�TK��Z�+��[K���}Hpٕ�|�]�ϯ�]����"כ�u�;�bl�N�oZŇ �ߐ�|%2���1t�]NMO�GB'��*12�2���s��o��l��A��ښ� Ӑ������������rK����Q��Q �1�aaaL�D}��S�憶q?&!����=AF �=m-�D��F	���ԗ���{g3��%��%����LF�n���.���Hww*62���nO20"~ �On|j߸���L�w=����aS�"/�r�bhH����q���x�� �w�IGy�ߣg��C�T��
��l�X��H�:�ez[I�x'�aG�I�j�L�Ӹ�𨩥�^��$ccc�ü�J�<�[t�Q��po1_f�`_�Nට���r��t�M",K@$��⫻���3j��><�z�x��d�����S����ם�i��KRT��'���[Zm�ya�0/������u��;y����i����
����~W�89���&80�drddda�B=*�5��l���_��a���s���˦���W
X�q�PV.�V��͸q#B�Q�k�� ����KjiM$��4�9����1t����INJz_m3v�8�D����7��\ۅ[��Y�GI �}������W���I1m�����q/fǚ�0���2-�ttL6���+��f ��֚��ob}3�����BB��;aX� �j2g=��B�҄��8\BB#fQ�HҎ{Zl2#������`����{࣑"#�X����`����~�Xb���!M�"���A�ؗ��::j�lTT��^0XPO��P�2�����~�_��A"���z{����.\�&ȯ���q�5E+�ӷJ&���@ǫ���]#ޛ!��ƅ3��z<����t_��:��О�\`�������S�E:���2�'�xx���{}=�w�:/9�@�y���+�,�0_kX��ɉwp*m�����36%����A
*��ȣ$Ez���K�򞌨����0�/͵���Fq}�_��,�[@Dt�^T�x?69��\�du*�!UR-b����x��e�ӕ�wvԌ����Q�O����o�)�"�H�X\R��%P���6wJ[>��dMD�;ЏGӘN���-9��} i�}곐���h7FD,��ǣ��?�(b�b�w���f�oiL��l�e��������9�����!t�S��*�')0�0 8����i� �c9�O��n�F�C��tk\Կ�bv�t��r�U�����9�n���ng�>Y����\�������@� x��$ޯ������Lc #��2�Hgb�h����X6�����@�	z��ό����nw�!vI��9�)k=�_����-��-�(�&o��+��4yrA�=O�^M`R���!��u�2�.�x�yJ�o�m�s���@���<��6P�@�����kf/�#��ߣ�4�9�D���+�^z��ѥ��� v˕%%%
}?t�;K�N��3�s s�O;�] $.|m��Qu�UPZ:lc#&�u�;�H���k?�$
��cԴ��#�m����=��W@� ��U,�sx�\����2;{D��Ä�Ö> �)�1���`��UgN �f�R��x{���~�M��޹��r��ʅT;g^u��n�N`$Tq]�n�/���[d}��i,�d��=5���1�qVTy|�T���_��y]�Z��}x���Y1��y���W��a(1�U���l�rpR��K��X�vp�)������m��1�'~�c�񤦯��-�F�C�Q�ٙ��@2B�8\�.F�r8ȫN� G��#�$��M�K<����=��rM�ߤ�9A����"�k<b�F�5���.)ybhh�{PT�3S��) ���v���9dvbC�-��F|���s2�k/͝�S�j�ÎD��ᦱ<�UB�:��h9�a��j<Y��x:�������)oh��|�Uggg�MB�k-�(ٕ���@`�.�r��|}}w��/dЪ��+�Ѵ��[{'�Q9cK.��o��uvVVk)�����7�B�ȈT��t����i�B�33���?���Bb�7�j�s�=XЎW��H�ha͒h,�?P���ֲ�6�24�C�)�ޑ����&���L�����M�Ƒ���5�W^��U���}Y`�S2t�LYw2�ё����R2�v�`g{����_�>>��Wth�����e�T�w�Bi��h��Vǧ�|�y��B�*g0���J�їn��h2w%sYfM����!}a}TP@�4�Xc�34=3����*8:=�;�nN����	�u��4��K�Ĵy��{PFJJ�ׯ���V���&6���
gS����r���[�j�`���pO��.�S,7Bs���!�[�%X��~�P��J�I�,��n��/ii��,�<��y}{zĺ���P}�r@
�������)���w��Z����������[
��םKGO���vi�_�h��j�<�l
��t�� O�9�I
��f�1,\�%�2!t�j�{.�U5){a`@_�~E��",z���������𘳯�Y �G]���0S�R�J�1*�o]��ݩ4/�%���[��q`C�8�T�2X#}${��t �c��?��pssgegSQ�����B	2+�x�jV]�c,r�����ݯ7�f5��ѻ;�"ޖ��
ӫ��_2��z����ƭ^�KC�y�%�"�6��ǩ����s����z0z_��P�8F���tL/�D�S��|��MUC#�")#��R�%�|�]�H//���Y���7��$�]tkl����������qm�t+��h�SD�����%�uvu)]�K:;;C9��qޞT�9�\�B�����_�|��!x~'���G#������Z^~���M���,(���|�
�b]�P�׹�H�[xd`�#R1��\^�k�]�+���UQ��+�xK'G�n`�����⪁��]�԰�;r�#%%%9D[4��Ԑ���&��֒ ��Z�76���+�3Vl�vq�JXubZ��� ����5H�����Κ��H�	��l��3�Q��*)EO��:�-,(󠠠���Hdr�a���c�-����#��� ���Uv�9:r0>�+..���MJ�����+��ׯ���FG��|E����JF��$LM����E�jkkW���Ӻy�g�ܠ��<�ƪ���7��q\�DXbѝ�ﶹ �[[�_��dt��E&��/��͠��e� �&y�rѾ���"f�?q�7�&M���8�#uP�n� �E&=�5A$��j
7Y�����V
<���?0���sZ�%�?}�t����_�����C��54m�9!!��:�;s��4AT�ә�Ξ�ܦ�9k�l�pF��x������������ظ�A�(T���-�Z;b�ޟ?�PPE@��� �� t~-�B�:�s�]�b|�.6�OJ	����2��Zw���u��"�B�㵗-��xB�k(y�L999�����ά����0`o���G&��ΏKK�HVDNVkk�8==�:��?Em/Q�e>���rG�H��$m�y�_�9�]��r|����s��ҷ���ͽ=i'��443'�q(333P%��:3��~.�b����7
��������	��|�}�N��`:������<@ڞ9�Xl\]��,@
$��~l��J�uY��NAދ���j���6��A2n��s6���b��[��{�\+��gl3���TU��f���E�'&�l�TTd���:�^�$�Sz���_������>J{0h\�� 3O�XĊ�n��]7����(�P�O������J4!��x�t
_L��Tk0�(s\�A_�q��/&z�I	Q�z1f*Zn_0�>��(ς��å���}�};����e9��'�G _��6X�swu-C\���f���;�pw�;<6���+ُ�Gu�SS=�m��E�I����D���"#ш��C,AN�A���;�y�#�ƞ2�~�|�~�T��r�!��>�EÒMʎTгD���\�����NrI��^II!v���2�[q��t1ODno�pC�����4V�E,_����i�'&B�9�ҕI]Q�����4�͛V�4��N��F94_!��A�
��y���:�	�iv��iZ-���̺Р#=���Y-��`�b;�LI7X�K��_���C.����(U��VQY��3(BO�m��8j���K�:v}���e,���1����ՠ(��&J-�����iY.}&���r�Q"�W6������[��f����_IC��{��=���w�W��-f�����=����K��n�����{���?C����	:��ɩ\G��Mu�:R1??t��E���g�z��3�\H1ç���/��Nl�4!�p�����dօ��
�&�[ ݵ��O~x�B��<���x���N�Z��u� ���Ԩ0 D```�.;�A�M���E�^U�����I��^;/l�P��pSdK�a�L=TF�J�	?���tpx��8��	��;Q[�������Q�\�M�O޵���PS�s_��yM-1�z6RQ�(B��>lQ��S��=1�/x�a��� Gˏ��̡)ޟ^�Fn�h�CW�Ʒ���z�>Z��E�i�ǻc8�2�a�'�bVi)���^�U��	pG�´�_���[�!�/3!X����::���N�KV4'(�HV�ZR"� P�`�Adt$:-.!a�ɦ.�m�$tB�i2t��\%H7���>�ؼ�?�QA'Ï���~�Ĺ/:0�>+[��-f�CT� �pZ9Czxo�9��v٣�˧65�/��'D���k����dG�p���Y�~�I<�
D��t��!ظ���e�[� �С����
�d���L�y=P�)������tYe�X��EA,M���������k���׊f��#�����#cc��琍e%���9��������k�n���F.! ��-%]�!p�)i���"��H�tK}s����u��sf�<1�g�I�����p5:U㖼��^��(��_�~�UM�]`���"�355���dė/*]�� ���O��aY^�]y5PYZ��hv���r�{-�O�N��襎����C��*ދ���
��,��K;����-Ye�����/G����r���鍓��zAJC#�f�J��
�;g�I��Ն��h˟���9��C*L���YB���kP@P�}�f8᧙��b�0RM��u����ʗ'@#��9(**���o	�WTp&�l�����}s�t�2VP�W�?k��yK��0��;�ؖ�ZQt���/�Wz�@,�r�}�B�_pIIQC�	wqE�eU��rφ�[�<<=C�ɡ�L�h�yн칳3O�{"BX�TH��Fz��P�D���
���_�`�7X���_��~�K�8�4MMI���X���U�H��4`?�8\!��	��(+�����51�����"1	I�:FI�<����l�>�� )�N6�.�\� �u�������ɫ��W��2��ߊ����P�W,��󱘚�w2z=�u�<��*�P�z51����B��{ ��9JN���ʺ�����5�e�d1���Z7n�UXK�� �!?�67�y	�f)T���	�2f+77u��>��Qr�>�P�` �{xE��4ld#��6�����z�����t{&�շ<�8k��R�͞����9`�ґ��'�b��`�� ?�-Y�s��U��,�o8�΋$@ђ�$���� �P���+���=�Bn4�V#��xef���l���F�Y�Ğ?y��JJ
*E��/�_��yd�J>(��%t����/���\�:Ɏ����1���H����� $�eq-��>H����r0+WX�����g���iY�)�d�eaa�O@���kH!�������n���f'(���� 'J�5�aT,
�UK+0�����Ӕ�j=�iZ��������BR����ٶ�m�i��S$��1*F̴E�@��=K��Ҳ]�EK��&�ҏ�kzc\a��;5��f��74ނaC`����Xn���zd>�?�T��H�"}->D-u�N�ʊIL\\�>��+����݌E`ވd�,,1����*u�7��.8?�@�Vt���e����^�.Yt��Ȝսi�%�H.b9�����.�?�DlllCccg��O�<	G�RaUK��X1茈���A}X�����p����}��*���O�G,;�Yh�'�m��Q�X2?�Z�V	Z�G�p�����\���E%�̌��<�߾��&����D� ��!Ζ�#�k� �@�8��Fj��%k5f �~.��� \�/������]Ͼ]O��*>�3Ʒ����k��OX����s�r�Lْe��ѣ��׶X��_^�Gٞ��&��G�>��:M.,���(�9w���	�!���a@��?0�o\�Ps�Yc���gt�.x{�����م�P����~8����@7��i�rdl,\�����6?�/��2@5�tuukz�o�m�=��a�cm�/eś���B:eA�BZ4333��-YI�~dÍ��!��L�;&..X�Y��P|)5��2$�I	@�
3tI�Ym�	k-`z��|��H^�E�}ySPR�=��d��������c����������c!h��b���'�B_T��䃝UE��+�R��z�|�ӝ���>%����7v^)nݷ�C{(�s��������dzI!��pIV<϶рӸ���ܝ��{ӭU�@Z��"N�h�f���I��$}�65uW�ʺ^��D��qM1�-�7o��v �'���阮�a��N{c���;�e�)c��w�(@�̼4�us�+�ܳ�I� 226nP	�#n�/�����V��Zss�O�Φp�a�z�4@�B2�Cr�n=�����jo�d�)V����0
��)*--,,��ZJDn$eif���ðw��RNE744��x_B{Ҩ|�����e����E[g秆���h�����P?�b>���J��(hS���<����Pa�$�IzI��D�}��������_�p�A z�''MiH�8sDD���0(�??�^NN�Q,>��uE=r�}??q���a���j��E��x���� &�p��&�ɛ�����[�B`񹸸� }��_#'v��ÇQ--"@-M�Q�}o�'�6rW^�W�P���n�/����^�n�w��`��9w�ųVk#�eÜ���+#
+W���W��Ϸa���o4�5���M�)A�:��gC.6W�KV���8�[H$Nk��\�.�K�Tj*r�Z��5�-*t�:���޸̂�$k���C] �5444#�t����_i!:�`+})%��i�Z�Z��T!x�VSx����f�V�����S_�0�[ܦ�:�??9ʨ������oMM�ݪ	�P|z�������8g��e砱����M�������q�K�}�Ny,��� �U)Ӟ�<���S�S��Q"æ��S��m�����r3��e��p趉�:B�&G�F�8���B��ErT9��{��4�U>��f���ݻw��$�kiK���,�ǒ���0����?;2՞2'�/u ����܆��h@�-�If�sf��U𥹹�����	 �x�F�s7����#�!aT�T	�k��PXK��&_�݂�K��k0Y�N�����0}R?P�)A��/E����^��W���	[Ђ��S�F�gŭ�QC�֖{�O��ô���;`a����͕-���蠖i����w�-)i��f�I����OB�ٍ:쩐���o٪62;��J�c���2�"驩�J����tttP��!��~�'A�et�g����Nq�6�|Lm]�<ݯ����J�rϹz�i�Ώ1���M��M|}*���S�"I�iד��ErЕDx`����S��� b�MO3p�Gs˺�����v�N<>xF/@�z�����
�+�#����x�&�_�=�E)�[����g,�sr0��ӆ-��$�x�6=}��D������W�bB��X�Cjhn�z�&S��R̃us]�0�������Q~� ��t��ϐ%tBt<E�;�tJQ7���4�$���������g쩚!���V9���.nn�Ϝ�`t�M)��d"��Ɯ�}�]�\��ED~����@7��>�p�\��E�����<Sr~A����e Ƥ�G�������홀��3����y`t�]u��K��S�r~�����rl؇���Ұ�WT4�V�]�^�$� �|��&<�X����l�Je�ς�=�ۂ��2^b9��e�EpGFFj�8�ْ`MdQru+gf�o7m�����%]�]��fZ�N�`c�hDF��7�c�U�0��L��_�=�z�;��v55��P�XS��+ί���Y�^�MHX�5���y�~���o�B����&��+�xZ=��)�>�T�� ��r��[�PgG�tt��o	˗�Ap��Ąe�du�^�}�{��x��T�
NN[����ksH��a���D�{=ލ����i[�p��A��'n�*V�vg5|�[���E`�L(�6Ws��}�76�U���wu�^�ZMfU/���u�_�9���������؍ F����tt-�Pĭ�h������
�"D՚���6x�3�o~�c����j�[c H�yXN�H���
��X���T�~���Q N���S�.���-� /v��F8�_Z��9���W��^�E��
?~����IӉ���|�̔�{$��.@�M�P:xi]�F���m`�>t�I��iE�.@��r.3�����/ے"Y��
��Wj

���n���&�1�î�s�e3Tpwxu�����WH���ʳ����/)))T�'-^�����dT��ײ��̛�kkj��[u�חp������~�AWOw��S����ZK�H�V<�c�jaq:6�����`V�%����fx\�|l�I���M�P��X�܄{1!���6�L�;9��"<wdn�x<S�C�v|�ܹ��,�j9Y���}1�>@���Еh��q�_����V��OL뇡��O>�7h��R�\����js�8�*�2�@�=
���@�_�!�YC��~.��Q!:k@l���+d���9	�/���UtBa�v�P̚�O� Q ��-X����qf�`�Ϗ�>�^>��ppšvd�Ǳ�����i�*�uI-`C����~���z����U �I�������Qa���{���W/�ii�8�A<�x��܁�P4����0X0��N�pǔ��攈(;�Ό�/Cg3��\�cQ���ڽOEN�	�j�ӟ�
���2ģ޻�u5-�~*�,LϜJvJܾ�O�#��e*k�
gft>Lg򫪨D��&��'��C ��d_V]�`@.��DCr�+������A}�M��l��������n*܈���7K	���~gz��Q E��prZl�(�������Hٙ����}P<�$Y����a�)疠�����-�k
�]�f*m_�Zq&��q�Ȼs{GxB����Ůg�[�w�BuV�@�)} q����'�
5N�ϡ������&���kZ���FzhN���i;�{��3�i�����h%[>�bH2���;z����h
�+�T�z�%�������#���I_b-���b�qG����o���,��N��TT�|t,~ݢz����;��Ö|�;�G�{�ZZ�����h�x���P��9uC���;�� ��fz���>�H������!V�p��<*��N͜CFvv��c��ķo)�-��_����}���Cu��y�ٙ�$���� �� �%�'��Z����>���]��ô���������缽��k&�ϊ̲:n�[!ʻ@�:��')���sp4³ֺ�;��{��X���uV�����l�Z�۳������A������*�x9b��=�YS�6���C����#�mƩp����_��?9I��N�0q�\=��@R
�/����z���t�Qs@Wn,:���1�<#��0}�������m�e2�����څ���\��9�z��4����7��A9Kfn��Br�ۅN6�;�Vcx
>~����:��=��S�P71�==PK���8j���e��KIF���LY�7�����p�ќ��x���i��ΞZ���ȠR�N��Q���F�t��L���j���Xx{�(j,�<h�����x*��F�9j���uL����J��k�x���#�l5�P��z�&��$���N��y�������e]�Q�X��ۇ��e�:�)��=o�D
]�r�s�˴1�= �$0���w��&�ޣ1�.�5��ۯ#<��5E��?6�˜��vu%P-�W$ؘ���L�|uy9�P�sR���#�1f�� �J�!��}�A��פ�:��Z�>����
8
�a��O��������<���V-]۟�}�VRR"�(Y�bY�\�b�����d�R�Z�<vg姙0�(JOK��a�]���~[\��z���з=��q�n!:9o�8���ׯh��D�M�8-�Z�?|x3���:*d���-�8�k���O�	��^��D�Cw�y��aY�4�WW���$+W��e%f�����Ee��ͺ������n�x������v9z��/���.#��׿��ĕ|L:~�㺏١KI�h,�IM�~�����mc���]3Kn�o�β���|y?Wy��f�,(������j-�e?`�jJ��r<����wa$���*s�`zg��TGECs�80���Q�=R*R��K)�ki�;z�o�M�/�Ԗ,NBB��GYB�������uW."�ڦr쩫+}J��kJ��ѣɥ���1B��3\�,���	ئ�G�@%� �{ޝ�t|ǘ>rxZ$Y�R��i>,R$���ߔrU\��F�1���i;����l����!��^�F��#�����#��h �����P\��a��ݳ�D'ѱ >0�VKKJ���<_��4\��N/V���wťǂ	�:Ⱦ��I�&q��u������σ�����|�fv'5t����� �RRO�������4>膳נ.�Vij�O��t5�z3��УR'�0C��yfjj����vK>};����M��Ö���C�Ԁ�KJ�:|��	`G,��N��9���;�R�u�-���y�M�_]2�v���S��Ӈ���(�<�f�T�b��J���?��H��D���Z�H��"��{�^'���fh��8�t?�����3���/�	Xd�t�_��B��۾���A��dKAh�D��&j`hXtH)�����PCW�猋�55o�qE��S�Vg%&��P�yC��]�����~����Jn`� �x��X̬�3ml|�A��DS5l��-L���o�7�}��' ����i�Lf��utҎ=c�X98�E�W^|�i).f
|0�����^��*��kER�|z���� t�/z�"n�l������?�0�΅�r���i�(���;\E���Ŏ�#�l���M�l���#��·+4 �]DR��>_�:f��[��
�Y�"q��ޝnHxV�7��&��a�z�=sC�~�{c�)"?�8��<���v����q{'�p�� DDD��V�
���N*...��<v�ɹ9�j ���=�5zV�OZ_r�:Z�&*Z.ޛ��5�yțf������ �I8���x<<r�$PD�c��]����]�����3��o'(���TT���w/�uK�+�[h*su�ć�&K�(��0���|0{C��i�E���8T���������tS}�:�ď��3�*��q=<<�F�v`�)$/�=G1ɘJ��{��8l�l0W�6�{���~������&�(��ҙW���z�� QNq�ш��Z��U�}��$�����E�˪u�Td�}������.i��q���������3����_��'c��$y�#�Ҟ����ͤ:b�b�j��P�� �_��;|���#�����6D�鯬�K�D���O���L��]�M�F���Y�������CA?�̴ײ����KN�!����hV�?$�z��FUpXu��! ���$E�e�}� 	A&�W�[6��(�!I:�i�sb�w��_p}2��@u잙����� 2¿J)��k;m��\�~-U#s<�'�_�����3��	:����������r�W����l��~9?+�j���(d��X?�]�(�S�o΋-�(/L�J#�Pa�s抑l(mEǋ]�w^3}@��J�G�}L�O;�Ah -Qi؜t�
�t%f�r1a�z���KhUa��C���:ւj���&ў�!��6:]�??����:昡c5���T�h��9	��.�'+L�x(nh��Ҝ�E�:�o)	���ekʒ�l$$� p���R����������pc��E��w-D�k1⎍�E�ʁ���[�w��}�,�3�eX��A������Q'�2&�&���iw�Q�@
|g�K[[�I���Tz�Z>>cbbؖ��gz���I�;�����òÝ��ɬ,Yb�5�T��6�'�#�r��o���b�mf��AԖ�܌�|bq1 ח�1���ܴ�G���[:����(Q�+�{;�Q׉��Rl�B�߾}cl̰ G%�y �v�ݐE'���B[gԤZ(����5UY��B�=p�'i�
���M�xf^���߯�E�h��9>F��ϟ���٪,i���c�-׺�nx�M/qN�Hn/:��X��MJ?_�%�o��͂.M���X^ ��K608�va�v$����>�>K��#�4,,,Q2:�;h�qpp�����Ġ��d���~%��+Q�"����h������IH��c����Z�H �d׈��^��A�,��Z����s=V��O��4#u���w1V�������/#ؔ���o+f��e
'ѩ(�|�44���33�A$x�<��Z*���˩�b��I��3a�S3��G�|Y6��y�V��2�e�y#j��VA;�݉���Z����o�E3��]]��{����C���KC$�t�v�AD)x�Z���łQԫ�Qdl>��j	?���J��0I�9=���L`�\�"��ȴ�H�/lЕ��sLI�%���/�2c��-�Ik�8��ٓ��^�b۵�/�DAf�/UC�����Ęϗ�m]��)�����ry�{6@�A7*]��@}ɑ_���z�4R�bn�����^f��ѡ��|i�L[��i�;^�xArr���~��V�~�v�9�?������uJ�bؐ��T�ޞ���k}�K5#��쮇iv7�Q�٠z�������%V�UA�D�듻%EE�zzzB��q#.�g�83U�Ա�_SZ^E�V���Sp�����?1�>uÝ�� ������V��}@i+�D�q���c]�qz}�sܞ��Z�mS��%�w��D�l��.d~gbgo)5���k�b؇8������-a����,Clu�D('�{V*���,�j��x�j)��!��ϵ��aЭ�`�F �r7�pC����������?F~ʀ��V�g�'u���?Y�qkw7L�|`y��<kM�ڕx�=$����q
"9c��S�ښ�O�,���2ZZD!=f?�IJ�n�����'�c ���3�������eK�	>��b�4������kE�:ߏ�sP����$�������Ch%u�V{�W����Bf~��l4�{��]�C�!B	,�#�4�NJ/����1��u,�W�?
��L��޿x<���gL`�����i)G�V�\]QA�/Q'f5��w�A^ �9��RW ��^�j�#�U�D�V�ׂ5��C�y0�D��{��4������Ъ�=��i�p�V��g���fٓ!~Iɜ�[�a^�P& ����R'JT�t������%B��;�'a�!��j��[��.��Z��~��s�\�r͗�."!ݷ;��frQ]Ŧu���iI�PBe���\�ɟ��,|��x�)PѤ��ĽaXd'�R���W���LL~&�m��v#��+avЈN.#@!F��ٝ���P�ڜ��Q�	 �I ����V1�QcY=�,�s��|��	s�{�%D||�����A�~aGGG	w{^�Oh�?E�!x�}}��9���0ɟו���kO}y!�&�� �&+{�}E6��|}-�ks���3V�;�\Ê�v �����[gth̈́�444��;�Q���nRM�qķ�������UAr�Ohy���ѷ���w�>{3`�!u���ݹY[�:]�$����a�Zr�u�y�D�w=N�?s�,ہճ�� �6q�YA��i��{m���Ǐ���,�8�3�w�$����\�j���,+Ø�%����T2Я}�B��#������GL�\�V�r��2��x��g��@���5�녲,K�Ŭl«������BYRHːebggo�����jd�pJ�۷��>���_aa�K�T�e���[O������� ��},����*\ =.�Ѕ�}��I3�M����s&�X�Ԕ��D���x��.�[���ѥk�\�=Q`;x�C��.K߮IG�p�!��R�D�k��� ��\Rg�����|UZy��zrr��P�Ls�+	�	!o�H�[�3������&�)0��E���OOO�g��{�N�����!W{�xH�RE��bb�Y�9Z�Iq#\�Մ2K�d˴C�D�fX�%jo�L�������8�\�d eB��,���	;-(����]={�EI�w;���#a'��l kR2��,�Sc���RBqi��t E�8/u�4���umy��������|۽�vR�'�y����t�''���;� bdk�˫���-b�i�{�Xf�+(�/����92�
n�z���Ag��BEEu�5��*z����1vh���ы�h����>7IkI0��@�,�|�j���-���A��T�YS��Ю\5h�����V���qj6�(�v�Yc�@AII8�H^��u�Է���!x�*Ic%;d�ux���������?�p�*�ɽ���5Y*�P�c����߯��r@T�I !-'�n%�b�Yki@477Cg%�ޤ�� TkeuM���2B��v�tv�$k%�9X���[�B!{��"���G<�㸷�b�x啹�x��8?����LKKk�=G�5��'�a�2��.���_ٹdQrЖfYY��q�SrS?𬭭��ۼ���. ��P"���0:�[t��Q_����j�WHH���.�?4��777Ho����>�z����F<��'�yL��}й����й+*K��ǩQ#х�l` V�=]����w�����


�RR���+T��@+$�~mus����/���P��*Z�(�6�����F�I����!+�@�����w3�e٠ە��?g�[���J�s}����u���-k�8(�@
��R���>�8;�lhj��^}^8	e9�ۨ�?6�4��G��Q��+4�J����s�����yE�=''��^�R���q�M���$���e����֧z3��''E������~��*[{{&^Q����DL[�.�o��7%���+�����<��6ߌg�둴��!+J�u%�kbD��[����	WdLRm)/�*���$=Z�	�[�h#-�du�Q��.�N�jD�q{��>:T7��[�A<{&{��;�AĤ���J:���qfmc�OEg�?�s�*g������DF5έ��ʨ�9(�E=�⥺�5��������1����]9ey߿߫�^̃`�&Ib��b<W�߭��\��g����vj~d3���=����l� ���]Y0�׀�^�0`�S ���y�[t,���3|0�����MܵD�n:�����-�2].Vb�|i�?��3�DZP�cŗi�! �q�Chs��f_&��\�Vg������d�V#Hpux�*N������;��xr�/K��Frgg付��Eȝ}��B]��6;���8?56�ጡs�h.��;AG��p�6"�b�N��y�"#��ͫ��޹\ʑ�/h�\����=�;��Ry<���;;b�*+���d����v�k8c��.5/��r�za��*��4��,��w>\mmH0��k~D?��<������ qy��>=���M��$�����w4����צ�h9�뮿~�d���@��BU-��Y�1WVbZ���g$�,�z,j�0T�������A����"B�ⱝ4�O ��gۄ�ȱ-|}�v�`�l̫��e���B�˰uߞV_��Q"�$�S�Z���0��-�_���C'��*>|xZ7�'� &�K,��N��s��z�kZG6z��K��!��.�>���n��!� �X*�D�GF��^���1�C�s����b_��5�c�&b�����Ku���i(���_.�'^�W_�-�8(H����=:�3�Wк�h0��U�ѻ�v��hit˺y�>v��! ��4�Ö��m�`n$��D���B���bƭnLo��q��߷��.��� 7�t/��%��*�h�`�kI�I���gj��H����*u�LsWM�P/�w��	�5׺�Y��5��XZ޼4�#�qbRa�:Z�;=�j�h�]�7���K�J�=�}�L=�G�r�ٔ�:�L����kj���#3^؉���iD�
)�Y85��M��
��yt��]	�u��˂9�n�پ��A� �S��2�:s}̄*'���D)��ۃ��y��*վ7Z�8���Y�gT/�Q�Sp0�6ġ=�����||�_X\��/�����i��X�L�`o�����K�5�~x�
����R��3���ggq�A��A�WTT|���n#E���$��M��>{=�w�9a�ZJ$����V���l5Λӳ� �ۭ쩘qqq�ʠ���4MN�t�R�<�|2ߘN�]M�9���v�_��mβ��EƐ��̢�y;�8���K %��W���M�y��t=��!bQ�uӡ���eE ����F�{Q	�����\?��ϡ�+]��c�ݏ�S��@��C��K; �����]��E �[�r%���3;N��Db��-����lM�c?������uVn�����,.~ہ/�z�K�ȃүlm�o�V����?�@����;�2%�]�7����P�����:{��G�xF�-����3�e���X	��+� ex�̧6R�UA����ļ�K�<ENLF�6A_j��Ŀ{G�Ņ�z6fnN�eq/��Q?�}����J/�	Yt䝳�f=��-Α����^�����B�w��%�����E�q.�(��;�]��,�e��>y�g �*���:4�`8�,jh>+�ߝ����ڑ��zi�*�Z�w�/+}p#^.�<�DcNT���sMTD�N�⚌�+� <q�k,(..��5�Aŧǝ�6Et\�q��=�o���cyV�:59=-�������=m-��/�kh�.R�d�
�^�ӎ�$�|�%Fꂖc_�Ȇ�R��~�������E'�i~Z8#d�<����xUۂ�y:O4u6/f��R�k�阘ɱ��3�32>=���q��0��f�釪�_���,��7������Ap4W754��`Z��v]>�G�#7�c�:�+��z�'J��rߊ�u��P'^������`����֦913�Q�G��c"���:�/E���%�gH��\�ұ���r��ʡ����ޞ�B+g?ά`8�ȱQ�L��g���icƯ�G�ᣣ,z�5ϛ7��k9q��>�����4<�𿫨����� 3����-�z��e�dnK57�r����p��M�[`��<��Qb��m�ʆE���@	��Ę=+.W_ Q���iR?H�L��[��N����-�`�!Sġ�w�=FNM=���O{z��߻On�:���||7�nM3��0��]RIH�8[�OD��%''����MX֚�Zg���i_(X���%�IE�!��"��@'J�]�cQ��1����+�'��Ȗ8��C63�% ���&X�࣡��`�J��1���i:���j`��Yֿ��n^���$��c��U�;#����㬞hX�r1F�j�=�Չ�����=��#���Kd%_��&���:��#���3g�70t{�c�=����9����L�_�ˇ�Oi�F�\��]�/���	{j_z�p�&y�T�������}��1�P�{)�����ԁ0��|��i��)�Ğ>�s�uo��m~�(�'eﲲ���3�Kb�A鹶�@�X�ɔO[E�]n����]?���PP�������/�~Z;4��D����������E��H[w:���Y{�|(>�(�JR0�z��Oh��ϯVίb(���Wl�<6��z `a�6%�8U��������Ķ�6��BB�ѫa�]ɸ���bZ\��'�Z:1��+]�g�#uM���gwHF1�aC�'
'Y��(��toe�Z��Ó�؞|��
�4�c�\�ʩ5w���@���m�A���?��T�\cP����v�\��Տu	r�����qc�ٴ9�'C�)�e��E�/��_����7ŗzl��3�g���/7ғ���¾�r{��3�������c���*.X��B����%� �Нk�����Cg�u�`�ն�(֯�����-�䖺��n���&H���S0�8��u�{q+���-������A���{��"}wL/�����Н�!m����s�j����.��5Bk؀NJ"�3�����/)S��\qk]vk�ih`�>����q9�3����_��t�Чubb���P^������I*����!h�b�����W�ʖ1���𠢢jq�P����n�V����!;�Ll�u1¤�F� w_X$*�}bŠ���E�걑nX@���(u57+��������>K��:h�2����,��'���V�Z�265��:�˴ш;<���s�&�j"K���K��aa��5�u��BW�6;x�*u��u�b�����޿]!�	�\��ɿ�)��)_9��}�i7�*�z��^���GLӋ^2LJ�C���*	RR�&&u0
�QM�c	N�Ύ��$���ń��O���|�UY��f>Y�".<�K�[���8��	�47d�Vs"'nW�W��,	ί�/���ȴu�������i
��ؘ����2-�����
9{{{��gVvv���?TW/�.8	W�t�C|Pd�i�8�����FA
��1{h�5?�*<�������\�x$���sw���b�Jsp,۾i;��Ǻg�H:P�[��Φ+eDk݁����~@��g5���lX�0Nt�诊������7=�5�ž_8���>��Gmn��7��cv���P�/�L��P�.w �9/L��i��.���^��p�ڇ�ʰi;�"o`��bܤ1=��}N�/==u��1�`zzz�z{����I7p1m-������@��Ǒ���1��i��Ɔ��/9p-�����e;y>�B˺�1�a�����ۍ���.//�W?�M`i�Q�����[I�TgO}�\�Ph�O��髟��=��E�{8���D�ߙ����X��p�O�hk�����O��;D<-��h��Q(l� NP�������E?`Y��G����B����8k�8�������V�^566*�?�;�z���o�}������� E�.h]�i�h����..5��|;��p)���GG��L˴���7�'c����n�ki%��O.ӭ*��rB���b�����U�����9�y�$�q+q�?��:��j�iV�����V
^����|F�G�)0�RKdL�B>�<<��r I��_=u��e%�<? �x���!���4^w!�'2|���hu�|��jƗy1wbƋ��П��V�BY\���|�J\�;	�ڽ�����q�?(ʒ�.�k�G�L��ǕŚ@J�A{��]N�6v�K��=R�;.[΢�K)����a %ب�M_�U|��ӿʑ�1ѯz���������{�ߎ� P�}d$� *����9/�� p����.����䌅��v�E�N��p���Y� 8�Ԍ�(($D��D�Zz��i�z)/� �F��R�Ƕf�=&�^�] 6��DQr�1!��pv�,�Q�r���T�8'A;·���<�@����t��ÖQ4�S�¦��l�#`�.6�BT��|7-G���?��j:���2 0���$��f�i�5ٰQ���g�p�<��~�Z"^J�X;�F�@!��HC�Ό�[�ߧSnfO}%�NXƼU�qJP/�>��vcr�VpN%L���������$�$*2n��'>�WR�)S���I��G�q���߄�Rq��aX��9T�?� E�c�ﾻ*u38$���%U��ܮH���ݓ6��B�{�1�Y�k�5Y��n��!pS�Kx��% �w/��A'��\�:7�ї��҉/*��T"d�h���מ�SSI5x� V5�1�ZGZG��2*Q� �8G�^L��n��z*��M�0GB�kߗ�*u�I���Ǉ�@������\�9/ܨ���Co���2�	�0{����&بP�!~~~���l�_��Ϻg{��B!�.����v��@����,S1n���3�F�1'W,����A`���˫y�
M ������<�	�Q�p�>��_�) (xx�J���ӳ$@���>�;��G�������u�֋�/�	v=�<��1�Vk�Pr"�ɛI#3Ú
��c��A��{3�TV��]}��b�2�^`�`�^w:�S�!�Ȁ�b[ػw�*��%�����ұk��119�xv��aݳ�o��1����謔���u���td�ͮ3Tݴa� �W^Y�\q�;������j?/�i1i����.�ߘ���C��C��M/��e��FBe�%�]��wwK��;P<׋�vL4�;-�Z螜�LNN���Zuٚ�O�'2�&�2j��RǠ˒��+tԋųl#}�?YE3�*�"g��J���0��\w��d�QE�4�3-�<���㽎���� ���1��үQD,��I^�xD���7ww�����`����+�����y�Ǘ�� F��3G���&R����'�����<�����#}=�'jj	�)(ʱ����=�s�����~�8��/����`�,�����߿^������uN@�@z���������ަ��>L%�GɅ���H�a����=?&���� �Z
��A��M7���5$�"���M3�c�7�K�����Xճ#w׫w�������g�C9A�S9223�+q��)����e�SKvXy���y�R���X���Տu/�t�I��Nv�)7��w�5�ET6OLMi�߭�{���ق�@�^� ��z��n�Clˣ-v�j����D�Au�L���6TՒ!A�w�v�'08�&Pd���ԟ������z"e��W��������WH�+!��<0RS������#��T�Jl>���\�7�y�b\DH��(k2��R������\Y�p�,}��Xчp~1q��`���r*2܈Kz��;�?�[p����-C*�U����F�ѣ� ��,B}���]E����W6�����W8��:����˙V�U~�qz�CW$���8�R��p�A���F[3'��{xyAg()t��N#+�l�n�i�y�:	V�H\�?3�%�_X�tʲ��K��P��D�H��T���GX���zb���?A�|4ԋ��gh������ʆz�����R�V��;1:��E}�����c�L��{qR����@�o(71�7$]g_0>h�I\T-^��2�����NU��˺�˄�>��X��ve؊} vk��ս��v���׃���v�^������H����2��t���Idxz�+˙���V�إL��#�9�+b@0�&m���Y2�����õ������"Ͳ��e���/kɻ�%��|||F����;M g�Zg��Ć����bP� �������Օ 7�g{纎��ɉ�h�W[�ZPPu!=|�Ӗ �<�j7�;1�8fƵëU�+0�@ �A�������&����,B����A��bT@`��Z�����
���<G�5�ji�]�k�Te�XI	si���b���o���;���>_�|���X�P>-!�H��Z:0 @�� t�n�V�4�I_�_��HveH��"< �e.ff��2y�31�˗ek���"#�]�ܸٛ� ~�V��O�Bg'�.n5oX/-L�}����P�2+��44d���_����y���McR-��]�p1h�B�Q@@ /9����� 5zC!���W��iS�s��&ݠ�`2�3�Y�5��Rg�����yp��>x��It�; }`�^�i���< D	��>:JMG6P$y���s��@q�CV�ʖ~�6�,�*��!��|� ��Ə����R�刧�r�����V�M�_#8�!����:N���s���T��N�%O��I�r[����뀧�{���ȖDF�&;������{��%E�B�ɼdeuɸ��[�w������^^�zq���<���>�9��ያ(���9����	bv�����.���Y��ƴ���I�?ƨq����ˊR�,!�}ư���ntH���j��l�ЀO%o�|w��r��ࡊ�
�z P��
��%�r***3�TyU��X�$kR���d6o��pQA���.eP�]VvrϞ�B"�VUz����b�e{t���-̟,ݧd\LJƖL^�;��P�n��	\�;�S�	���_N?� kK�d���nãM�����*|4򶶶�k��J�H��n��DI��j�<i˻��UE�����{�\;'�'���۵KF<�S�8�U4�D4{�}um�_Z�����(oll��M�]RR�u���cecÙ��I��a�PV(ʬ��N	8a-_���`���Ι\1<�8��DO�#?I6�d�cMP�Y�|�Z��_v������ �����"`��
��w�[3�B�w���?���Zy%#��Ձ�m�}S��p	6��^������-�\*��e��W���~*��>��o3���?M���m �-3队��ɛ���c̓�����ۺ������'�\E{|��ŤC�<��`x]�Z�8�:�w�_>*<C��D�1l���dffC�f������!o��@�	�9C�=a���~��v��~��Nxa-����R��"�DU��-��X�Ȏ?�ݚB���CB[�f66���,d- t������������ä��3=0𜈄�P@l���۾� �]�())�'�g�e���+*F���ץ��-���gw�*�H-�|��8�{�oi ���m�h��M��:�3�o�pK�HS�7:��|BB �fU���BV�@�P�p�cT���z+$ �5���^O&ϔ �����|���&��R��n�I}���3T��b���k�2ψ��8FOLL�~k����`@�V��ŎS����p�W�ӳp�@'E@�M�*Zjl[PPPl�y�1-/{ls H��co"b�V�J4��+����Qr�?�7��Ӊ��#E��-}Quub�^^�Y�3g��i��F�Mm��J\zE�0Ktbcb�Ok��t�k�xJ�'�jV\V�����:�4�hċ��N�s���M1�EC��h��|��4ߗ4��:������Y���g�� ���r(��'��Ć����m1�]�`o�����E#��>�tĊ�[����ڀA D
�d�h=�`.H��+.��N���N�&w�ی>���LZ7�L�j�OW[��d]>�,Z���p~@�A�v�|С�Qj��������c�%�ۘ�o"i���㳭N'>|ll,�U�]⌯c�)~�ߍ���H$�R�L���ʀ�? ����c��_���zu�¿T�IV[�rp��@O�gW"[��\ӇƩ��M~I����W��>~�S���a32CZR2��"��Ġ����%+���m�u i�4��8�}�(J,}��C�°N*ᅟ[FǍ�O����*��%GwR��g�!����Px�T��C1[}*  �/*�����\��̗!;	J�)\k�쀑�Y%wG E�!9���2&&�
_ܵ�{H)��^�x���ː4�Z�p63�pF����S��CCG���.o��70`�l�71��u�?P��v|�Zv�r�v��p���f ��d���Ņ߮���fff�f�����-M�<ey������%a��� *���c!8ɺ�������W��&BW�%�OIMx�h���0�S�o����-��-��dM�4����p���t��I3�d�����| _���n�d}�9`G�S�Ȩ}y�%{ �~���/��?E�?A�1�Y<�L�����������Z
|TH��?*�V��*v������ӝVPk��&z�J����1ۮuF�1Cg,��U�N�_5B��a�W�OϮr#���
C��_e� �N�B�KD����Um�M�e��ck��)���悫hE��|�s��*	"^�2'���:%?�wH���H���3�ΐ��/�!�sgVzM�1w���6t���ʹ�P�sW��߿	�^a >ĉNQD��Bľ�Z%�W�G�kU��ځG�05���C�A� ����i�H;�M�l�0����C�]a�/\4����_���������P^� ���j�-9T.
!��J���?��e�.���z����5��
��|h	`�CR7�t>'��K�J�H�w2�Oؒ')�s%}����_��ڎ ��MMM'[|3QP������<Y��e}�rg	 �1�^-|Ipï��jf���F���6�%ե���c�[�[�{�9�`��Ƥ~���Qٜ��N�M��AUU�`��۠$��'���g��fvvx!��ؼ���ۂ:��P}ԗ�@;���$�F��;6�ݵsv��_a�����:���D��zM�C��\QW�T��s�Ez2�7���w��_>}ֶG���a���=Ӑ+��F���&ŹAnD����Z����(�ۻ(Q�ϒ�'*X���+ˋ[ޗt_w(��q��Ͳ�q<@���`(O=��w�僕��S�
�r=AP��G��,�z=�������3w++��^a(e��=(m���J0s܌C��E[�7�&*7<1ƛC����]wO(1���z�Q��X���\E�恢������<������h���F]�@-�N�;<P�g6�P�5��CE�ן���@�+��P�>����I����Ñ���Ҁ N�&�a������nWvΑ�sz���O��{�ePGf��9;99�w:����Cp��0�yĸ����J���G�^ӫ�,d���	hJ[[[U��o���CC.�����:Nx��#�6����OEi�Y�k?z8n�UU�`٤�w���C����Y>�?`W�����~� �c$��3D�v�>���\ʹ�E`�^[. �YZb�.�Rק��,R7��|P�G���qCՈ����1��S��[�7��HZx�<�ZN+m�]
���{�^����H��N��Ъ��j��6��W�ͪLU��Z}j�;������֞��Y�ė{�}�?~�}(���Çe�(Ct�U汹o���R��}뇟���&�)�C����X�Ǧb��w�:[*,*m���7�����Fh͘}��nYqoqn�����[���-O��_x{�iݭdg�m�c%�E��ҳga E�� #>�ֶ
,�K�)�?Gj�i���8��)`P���� *Т��;Vg��,G��M����=��;|am�p���N�L���,^����}�֥P4S!�U��"UP�Vw����d�����/SZ�PrI���=��uI"2K7�/7�mdO����.N�R�.YK����t�[��jc�{�H'�ڴ~{�S9>�I����pW���wxSK�m2^0�R�����/�y@�@����&�y��� ;��jj�������b��H���M��{
\T���ii@O�!�����986���f/�+++��z�Gc�$���\y�Dj���\WwMH�6�r�`MZ��lP���S��	����?B���+<;@LL��9r�G&�B��<��yk�wdd$�����M=��J�5��~�����<76602���Һwс���*R�3H�i^K���O��7���g��}����	�+>11,2���i���j�g!�K\�md�r.���}����?���,0�}es'�#/��k�$n�U�3��QN�e��IQ{�'}|� �9�+�-�c;��v��/�)2�j�2$6�fv9
/�G�C톨�s����t��Γ��L���cy���e2=��F���4<�t� z\T �>��$�}��a�X�|B��c%�K���0�k���������{�j����\\o��#b�?���T ��q�Xۢ��xSX�B�scY.vv�'O"����7"�766D��h.�G��P�a-��O8����m�>.�����iii@��Wp6�캙�sOb��&r�&(i�xA�^t�tX�|ǲ\�O@�uO�
F�s���4�z�M�^�v_	�w����Pў%�4�)�TK�>���$�Y?���Z�>47bZ`�!a��zr_�b���DzNO;���=״��=�����8E�e��P=�[��-,��SoG��1&(������#����/.n���#޷o��&�~~~P9��u��N�EA�hi)O3���<��켼'u��\������;�=@Z�j3��{8���{�gM�ڵlQ���9�<|
�VQk�~����o1���_ėu�� ��E��aqT�}���i�eGh<�E/�E�7�r|�g�ONj��hc�d�N������1��N�rr 6�BKS�ݹ�l���7느��B&-u#���4��w��ئ�Es��o�^�I����B�|[!19y�m�N��s�c~�W9�p�G&n�[��� &����<��M9�v���oO���\�s��`D�Zȴ@+���3���ӵ�P�٪G~/-#:���IC���dA����``@��.h����P�IIX{��w՜EbM�W1�c�VV���;�
�/> �Cԗ��6���KY//!�L#�o(U��q<..hV3�'����o��[��`�)���	"Z2��F<��k�c�¸�F\T�@zL�uTpiq|D��gYæ�����8ێ-K���,��0�RX����
��:����u�������VN��\�p(�)kk˖ᷚBg�r�������獫S�eH{Nr4�6S���;=�����t��OLN� _p.��a˄OO��{�n?UV�����`�Y,)#�����̇_PpY;��?�	�����o����z+�G��ɩ�����M���K���UD�����d�)������[��x�?�J�4<6)��� rz=;(u{��??L]h_B��L�9A�&Q	
	)��[e��W��nS���q/T�e���Y_�਱o�;�Q(FG�����U�r��Cu0
''n�8�	��Q懇�fVV�.��|D�/^<��|���[�8�"Dxxx<����~?	���
�t�j���"]�}`y�.��A�Nlt4�(1@= c_�� ��{���@/��:O�۷��x���X` 6�wuu�"����=��j�SA�(�뗯��b���|Cs���Bn�Y)��=k�Rőy1�>AA
-��p���~
2���
���y����Ƹ,""c�#�f������ͤOS7��	B,�>�m��.!++��~�y��Ox�� {�S�ih�4���ʏ4��N��ΩQ^��*J�k��C^?d�Jr����6���U�{���x���
��m����mz���D)�6�����8���9a\�M�Iٚ�99y�Ӕ0t k_=i��H��t��:�����ibvlGk��}I�{@eCi���P��:���3([��L��SY�Ϻ�Å��7�;{�����tL[�T`Y��O���q'''%v��+��R����7�2��rC�{+��2������������[�K��;#�Je�[��������ݎ*�7)�m���K��m�d8A-���	�� -c6q�5fF�*CC�a���-�$%@�L�:ls�ɰ�f1�ej$V�k���L&�#""�W�q���C��xD�kj,@Ȱ���tfH��v`����Λo��0�hx Zi;f2�����R����i(�2���-zV�Ηɜ3�P���-����5�jޫ�:����ۍ��ǰ,�p�G�Į���Q�w��$�T��hl�FF۞�j�]]���02�����Ƕ(�:��]��#je�� ���/҈���d޻�_J�8]-���)�	~?��g=���b���j�R��lPs��lK/�"�J��^^^P@#`��������ւ�rR�Ҏ��2��Z�A��1/���s�/�1�!y������]�g�bǮF��v-�o7�����&|��(��=��xgG��G�&�W�;v���%ϻ��é�����A'��s~k�������)�d�������n���*Gff�Z���s��W�.�&0+Bլs5�댈STV�<�ͅS���w&O]a����	3�\����`B�
.C�HH�r5q�V��?2��/�q�XT�����l�Z����?�7�J
�Y���.9��K�X^f�a�Jxcjbhxw8uh�=Z�c!�	�uW���x���C�'�_5�K��4�W�RgV&%�-��]f�nO!���X������ӡ����{f?E������Y~�J�Ė�l��z�B9:6��+h�0іێ�~wڷ��H��`����K�(�9h�GӠ3�2��*"���]_�a�w���8����;�|*�s,���[�=�㧍�����pt�G}����/^�9�+u�3.P`\UKZ�x<���りwf�\�m�5K篽�g�vC��]NP��f3:���>Ȅ�uk�������/v���E 6/�O�.1��ȡ�����O�?�_A�'E�P��R�[�\�����^����'$��fd4���l��a��3�Q���IU�R�tz��ۀ�N����c�4��
��9c��,dY��.{��~�)�e�}����3<��ke���_���ᾤxQ*݇;d�غ&~J��%N�=��7�˴8�}�w���u��NӖ�d�wO�Z�%����V��v	i���|-�,s�g	b6Ƹ�{��~'��F��Jv��X\B��Yf%�B�ΥQOY��?*C]���R^W�:	��R��ѧ]v���@�E������`��O������v��X���/��Ѿϯ.��gַ���<����g�Z�ڽ/[����`��߇����kh	�W ������������?�b�$���y���Ї����p�'����k647���.��n�خ��hI�B[��!�}�X4R����Ç��.������8E� �|���T��4.�>�
P8����S�0���׿~���	�r�� �Be7���x{���khh���Ƨ��@�����
�1�t�o;xRSV���	��"Y^�"���P�ָ�"�Z�]c&\\�搱110g!������?��@�҇\�� PC����@��}fVɬ�������A4h�������lu�<Vd�������Th��������ğKH�8�����{�6$�@(<�u�	l���8T���	f�h��ż��aT�U���qpl{���_����c�'"f�9G��s1a6^�f�9��BS�u7UUuuV}�cX΁* �C�T��\���u��im�	
+8ux����^Y�6-�����Թ[wRn�>t��O�Y�L�K���8�麪���x�*����|�Q�k^WW�o_��l]O�(��B�8���#e�^n�Ø��n��-��� �w&�L����i�ZJ�r���h�%}�R��<�.������Ղ�о���X
U4�Ѧ/pg:$5	>��8�<=	��_��1Bw���KK��8��(,*
ډ�&N"}ٿ�c�x�iJ�)�	�z6�fc��e�gPTXxy3�
��tΆ�g�2�8�S�����ܺ;�������A�o~���`���$wG�{GU�c��9��j��KAZ`|���nw���k�J��������ڲ�7���kX׀�y<�	�l}��қ¿5 ؊9�wY�g*1���}�}LG���f�����R�ޯ}S*o(z����S4s�|�,����D�0y־���1�� �q�e%P�?�	���=�I�ǌ��a�t��MW@�}%jܖ���ǚ�qS�%=�g55<Lq����<6�kj���WQQ�-6T[)W�����l�vl�ڀ�����#��-u q��A
&�@�J@���tx�k�Cg���A���~����>11!)�f�ѻ�*AV��[�N�wUX����el�_@`�\Y�<���)�N����3����G�}�AF<�Q�;����+y1���LP��f�b�}5��ȇ�A��7�4�
��'��F���^����N�> X�vqW-]�r��](�lb���i�Y�y����oY�{����>I���`�c@6�F���a���z�S���O�Nfߊ{˿����z4L7Y��E�H��z�Rs9�4�뛛m���B"ͫ3�o�Ն�����gz�z�[xa�z� ���E��&(o�6T~������tk(c�$	�G��\�����������FF<Ӏw
@p�c&9�j�8�y�@���Iu%���7<��葲��5z7S�~����A�uL��-��޼l�Y��qm��j�����lÚG\"�� Hggg�q��>zeb�����n��| kT�+�,f ���"%��+�R��3\��?]���b1YY�@����פ��!���J������v}�����a���]��s����*]	������q�u7����G ��+��l�f�r9�L���Oɏ|+**��TB-�|�ԍ;��~��G@�i�:��Н^��MP�SۘC96&�6�;�i�͆.�B�Kj�Rq����=��1�XqC��Z��h���w2�1���?�$yC�Ws��A�f?C�f��s?���U��a�d7�w괹y��`7k����!\��L8��l������g��)*�@�/���W��r�)�A�I�ξǩ		�4D71�uJ����j���zM�us]8��n�	�Rޓ+<~/&��d�$`[�WR�V�rs�վ�2���i��bgi�J:�Ѽ�}�uľq'Q�EIE�ȏ���"���OA�kqoT�$�dt�&\�wo��'=<�x���w�d��-\RE������E(����
������^tDJ�$�C�oP֪�񮈥��(��v Vяʴ�\�L�w�8޼ ���:K�(k��L�6�X�O�����"`�0�My�|@�iii/w&�о�����t�������P��Iq1m����o�C;�����?o��nØ�ynB9�@� �u�q��П�a�-��瓻BM���q�-���#��R��*�ʏ%�ܻ��̹��|�B�O�=�Ul�=�H���sH��#���qiii�N�$ǌg	�� Ul_�<#�i% ���)4�N,.Z�1�h-3���
����Y��	����N���/!�j�L���)|�}t(f�1A�I�D����PYw��Ǿ����� �ޢz����S���u�"t�r���q�X�F����3}==���)�	���X���ѩ�����"E�j�D0�Q�js���<+��V�u�~�2#���x��"���[�聿_�U�obH�|c��sc�_@����
��(��Y��%2���[�u;
��� ���4�����E��G8�<��	�p�^���S{�4�4�碂W�4��z��>�Ot#Z^`��}*82.���ɶ����K[��ۀ�d��Ц�Dݞ�&���Y�ʦ�����)i�wyI���sch��Qn���_�뇕m;�nW��^\R��[D���7/�4���	i�x����/,,�� m����rA=���-�R���o^#���J�Xx!S->jd�����))]8S��)]q��-*㉂B�.� ��B`o*�]�k���(o�{��}���Hg'�Z��>5uu$�嫞��z\TԬ�1�A��<P˯���C�C�6�-X�V�M%�r��������<���IP2T��9X��E(���y@W]]}�U��iL*�������V�U�*�% j''�k4<[�Y�	}�+d�K��c�?ZϠ_��|u�G��7μ]1�lgq��;zI�;kY��n�qc�8��(�"-=��댠S�9V2��>"F"�w��鮆��~��)���s�ۯ��===]��F'.|����M ��A�,���!��9�---������������A:<�k����[��9��rN=��H2����o���6�L	k-��ݠom�m��]XR�:?�F��m%��%-�%w`j�a�uֈ�xc�V!�?�˪�-3�uMM�ö�m�����%�t�Aɻ=<�5N��&�ۺEkΈ��u2v�d%�������r���U��]U����ؾ����&1E�?����?(?�� ��9�������B�^4�[�kb�|�6��e�}{@5\O�·���'],���ۼ�w��5�8�f���jW���XP�� �PLdr�u��B�*1!��!dz3�~��Ն�T�cy�%�]�ӛ��[[����]��fi�H��W�-$�C�~VΥ?U2��E��(��P-��Y	ܑg"����r������0n�$��B�%W�����T&	b
PR�ʉ����@"�ZgwX��XƂ..�����ikks�vw'�u�V%�ʿ=�޴
�/�cF}�M���X���)�A*�~H��,�{���YZo�	U��ׁ��ԧ����?s�������rl��c![�[�8г�eg�	������צ����	�:W�"ɀ|�۰�&��w�i�7�0H����@�]�7u�l~@YY444{,ۜ�6�w�]5�)<<L���05L�& ���l�������u��9�&y��(@6��bD{T )�HV��n'@���0ܹm�OeG�n{Cɛ������rs���-�ڷ+J�:�V�tmx*|ew�4'����N�ɽcrX6�L��/����� m�w8��;�hr�b�M�?#��%�"��V�r��> !_����tkILX8
�Re�.sR�F��$w����R[���Y�変��z���^3��L/H��a�6��Y�#�E��U� �3��3jo9G�ɡ8K0?Q����x���{o��0��zIQQ�JWOO
`x�%����Kٱ<�S�A��Q7����YBe��X[[�\[?:�=�G�*��]'�ƾ+��g�g��!p�
��55눡4�\xEX��k�g��C]E�_wK���9˝����e3�{&�5fii�y!��}����Y�/AMI��sԌ3|Ϯ3����R���[��Mh�h~!�A��ܼ8�l�Ǐ{��O.Źm�_�ξ���xM=ō�&�U�n��גּs�H(����O�>������
X�a�'��"jsM	�����G������F�>@p77tCQ/����J��Sc�ϰX�����X���456�t�m?���������2�9�j%%QM��98�N//�x�LGC�H$�d�6�C*ݹ�h4_����wh���~�L��*�Hz�W[��6z��xkb�cN:���d7S�F�w��6�ff������TSW��^>tO�������h/+��c+���Y�]��4�
�Odc;, װ��2;�3���!Џ�n�>�=(���Ⱦ &�j	]�w�����"�N޶d� J�ym�����Ĥ�}*�su|��R!7���x}�%#�}xJ@JSӮ~Fշ�Bz�m#�v�W��%��� r�c��#�O|�A�!f���>/�����|q�	�yxddʃ�:��2@�L
�<�H�އv�����٥Ζ�Zߍ"�G���Q����؝�Hs�`��iޛ�����A�<��+����7��st[�|W�W.>��� �5^�_�!��j�����1-���ۥ�TY��uG�V�������uXj�f��A�VV�m��������͛7G�8|VG�K������Q�A㡾(헐��so�7�i_�#�z����Ɠ'O��գ�����*���e#K@�L����6]@r ;^��]�A�r�{��Ԗ��5�Y�'`��P���k}�K��>��K�.�J�4��צN��blgoo�Fm(a����(B�x&�����1~]Դ8s���D�A_�3UU�p8�?n,��jR}�����w3���/D{k��K����@��]܈2dd�p"[�R��*(�~���j����Pή3>8�ژ��k�B��9�k�u��5�ޭ�*���\dֱ<������	���_tO-#���s�Օ=_^�*���|<�l~�qxX2\b:�v�,���-�Q��Q@�� �	�N�Oy�g�9�B{��,��f2At	0�uK���'$&�����=}�t��N%�o{��R�4vyMM�����	J�k+++Y997�bp,����4*��x��0�� 'ww`9�5n/Jv�e���H���R�ک�  ��rB"oޝ��,��7y67%i��V6N�G�]LȿD������`q.D/.��}G�~&B�ԥ#
��R���+�G�-3��\��H�"������m3i�ig����_��|;�!�c�v��E'����h_��_�ť�*�|�R�X�Ku����^ɬ����('55b�G��n:˦�c�xU
�1����`��o߾�$��cA=��m�����ض����P9��?Oнm��ʙUNB.e}��Y�
��=ܰ���s��jppp��]�ϼ����4�[�-�x�q;��v흗����a)��Sv��o�x@8�o|m�>BI,ypU�kgrq��)�Ǌ�@�>��si�&�eݾs�N���05�w�������Q4BCO�΀c�g��������*S�ܜQ��ۨ��;�Ʒ
�ɯ������I	��R|�|�xdX�� ��O�=#����3=V"#�8m�n���-���adlYZ�H�6���q�&V�9�6����}(c
c�a�P\Rr��g���`�PgF\�-BކС<uE_�̩:�Ҧ�?����<������I�S��  �Z\��Od>>��Qp�wUݱ(D� ��ۋ���7׉��	Q�p+�$��+�*��o+�ݺM�lll$�=��� NPj�!����OJm��S��Ւ��n��M�����eKfL���=	x�����)Cdddk�	L�*_��T�PP)w�ˍC���t���|�,x�}�
�?��"-O�gb�[��ֻ�����R���Չ��F
��V&C��r�+-cX`�l7�>uj�S@�Y�VoUFQ1J�pڄ��ŝ1����
��pZ�y��ׯ��;��4*��&n�8�C�G���j�4��],�������I6�ލ�mz#2w�1�z��H8S2w��up�ƭ�v:��@_R�^�e@*����&��>44�6a��b'�O�!J�_: �J$��/D��wW�ފ��( (O�>;{�	��%��ĮڿP��ϟi�Y�������`X�Ӥ����Au:�OHU�b��L�


�w;7<��z��?�Lr��	��ܫ8�&��f�nt32�44��:솉N�8�	���*��G)��n#�近�t&0�z����6c',���\L�=)������ �j=� �����TUQ �3(���%��_noo��q ��^'�|� ���x�,R!g�\p�b�j�|nv�<N�RlWs7��@2������@=�/���p�f����Kdfu���J������ʪA�m[��˄禰������f�~���\.�)����!H�g�r��>.V��+)��|��g�S�Ϻ�l=���f~P>�	~P��U�J�e���t�-�ݟ�/�{P^��:���������R��W��-�h��2�����O��>u��<'S7P�4� �9��8��TTT�\��I�',dY���rDo�����46�p>{ <�z�m�%W���i��s!��c�n��%�WDm�}O��Z��svjiۘ�\{�>�5qᐳ�J=��5'-N��hW�%X#Tm���o��RQ����:	�q��immEb׏�oWT�G���6�n/�� y�����`,�^��$n�H�0�K�muu�����-���Xs��<�WaŶ�6��}C�A-U$�<��-�D�Af2�N�tPv�����˅{����K��$%�5�3���+��L�IO<q���!0�v��*	گ��x��~�1��f�������?�ڍN5�?�����pm0���8MI`�g׿�[4򇴡=F��,X���ʄ�4���@ ��q��<�����
%C_F�
� ����k_[o�+��n�Du��mj�C-���+D��~�1�F����/��A���ڋ�S��װ�g�t�H7'+�q׽� ���GuF�������QdL뽝�G4ccb���H"�*܊��H�;na�ޅ�,:�z����Ɵ�n/�Ls���BK��|�8H�O�㥟�)W7tZ��LX�	`��޾��ڴG���o� jj���.�1`�����x��������k��b-*f��RiоP+�i0Z�k�:#����\� |��[�ÖX>�ţIς^�3��&ֶUp_m���^B2K�
����1@ȵ�)##����i.#��o�1m�k��r���~y��j(��tlΕy��$ �!�%*�t3�Ž��OY������k?���w������n^������K]��7�0t;;< 9��U�())A\&9�`ʟ��߾ڨ\rv��17�����R�����>�p���oPV�IX�S� ǀ���K��)�%������+Mww��E��6i��F��iO:P����:e&�3ɩ����� �a�����j.\� �`Ȣ��8_^T3kxl��
�8�Z����\������\E�u�2n����߉�?��"p,���Ë��s�&�DXX�?��e�"�ЬʠD���n����n�J�ʪ��ꃮ/����R�n&JA'(�����n<}�q�b��ؑ�Մ����gޡ��7��R{׷�;~���4@�S�X<d��m�/v�W�����ᓓ�A�#�B@�7�
����wS��W�˶.��W��.π�Jȋ�U<`���.����<U�K�_�7D,K�xƅ{���,)�ZF���߽#�#�0��	�=\������L����?*c@�����ʧ�EO��,�]*S`����������AI@3�+������Q*�Mn*B�{�ዋV��rL	?��۬��^]]��Su5l�"<��Lxt4~�ȟڲZu�,
�TS8�B���������{	�>����sI��D���ȕ��ݿ� �>����'���L�o	@���4���;���T�"�<���;�\��a��+֯�����75O�������zM�cT~�칞�h�#~T�+0+���3�>���/�%���%���`���ɉ��gx����h��'�>�(�3���@z�f�O��8�b�kk��%w�He��;wZ8:�:Rz�����8j'(�{�q<��낭X�H@��	�������F�aZ슆�&����ToQk9߿�|�ä���]9K˜9��i��Ix|������¯����=���I<	�jTMM�w�D�_�ͧ�;�����x)������J�L:

	A{���������ڟ�ݼa`h�id�q�Hӧ�:�@K��������_Q�Ga�\2�������Zyǫ��GE���}�"�%}{B���0@�����W/��H�2���l,�oy�5!��v��{�NAEuSbu�%�v%ɰ5�)A)�`��JʹR��7�_7^���
�߳��e���G=�9�(��YNT�0̠{w�^�������A[���H ���

g74L[R~��'"&v�t��{yrG�U��o��2�E�I�m�/��&*���f���q.m�k�� ��''aM|�M*����h0��ѣ����%ؐ���i%Ќ�%�It��r��G���������Z&�w�{Ϸ�H�]̇U�k��9���Wf[��t���k$W�9� -��G��aJFw������4䕕	N�t��x4hsP�p?���*v���OX�j���Arw�7U��"?fz�e����PA~��"�֑\Ј^�K���<kKAM큸u�x�U�� �f�Om��b�>�c,/�"��)~�Fc-���( (�qF���ݎ�WRQ���a% $�j�Ɛ��<�\]X�"���ۿW{!WR�أ7�L�8��gA�Y1V���%M?fv>�Hf�i�ُp g�.�␬���$pn`gg�ҖQD1f)*�@'�/\|>�����_�x�h�˕1��ѣG;1s�0)�����!�p:F2�mJb��EA�g�$�`����a��>ЉQmp��@�ល���cKKKR�[)eYYY��J�HHw��06���a@�՚�� ^���e���Ϙ �Ҭڠ��P_h?E<��TWW�\'�}Z���NVV,˻�\ݭv��t()���C
-m��hr�0����O���.�;�Z���jJ��pW�t7��1���؍�/��]���N;x���[#o݅�#�N�Y@�.,*��$"c3	R)c�C�e"o�<zerC��}�<S�k�O2���z���s;Ĕ\!�Í7��`Y�ww�gw�S;,^)���J�w�,��E�$���='(���%�Z���kw�-$?���3���bs|�h4���\T���N��"�7�H9�ɴ"ϾC4�js}��9��@�m�ҳE�r���+���:��=}@˵}SfI�y^�,���k��p�]i[�Ĥ/X�*������J�ѵܯ_}�����ɿx�B������NÐ*�q\� �`�F�;!�u `yCuV����d�<�o\&��|ֺ�۱O���"�-�n64H �i�k%�Mu��?�p�<�i�]=��eN
 �O2�6��M��.u���\o�6��W 7)~b�4'�� 1L�T�D�q½|	g����k[�;�5P��woOԄJCTUa� 95l/�pOOO�WML�x�jj���'�@Y	

�N���Lx��+��|�~ivu~d�r�ӣ�8]Kztt$����ʂ�<S�|�⡾�a�d�q��k���Ol��n� ��鰀�m�Jy�3��NQ{���:wySHH�<��S�:�׎�'��~����G@i�@p�ڠ��2��+p����`��' @���s�t��x���∐�?��
|�Dg�!!!!?.��kiiI�{���������###vvv{J�x��XI�I���Cy�]L�3��:�!�����{��w�^R���t�sHu�1@��n��c���6�o,�� �"�ʝ.ƺ-��7?a`ce� �y�;������L�I��E�7#���o�"�O{:;쟛#��.h ̅S��M>�Ԥ��]���]���O�:�(������ 
yU݊&y�r��H��ڌJ� ���c�7�^��\����n̿�n�y��s��]ZT�;Q��� ���ǘ��M���������B�N��2<f47���d�]>�]�b�|���3���"�MTK�X�ȫI�ɀb:��=��0o����P�i*�b8LJ��v���5+׃�Q�a�󫽩##�yHcmw2��� �e�U9ͽ{9��_�x��Ƅ��w��Srlw
S+("N.��O�d���5�7��gƋ�R��O����f�L�B����"�_?g1^�G��/O����z�}_�u�����FKK+��
��UUE���ӿ�	�e|���Բ]���/$�y��}1��5~�/ss;v�oÔ?� �V�5��	��(��F0�Ƴ�-���N�J9���1~�M �j׳ck�ʃ� �_9�|�k�0|�ޮ_È}�Z^����C�*kш=`8G����ݒ��"�����]V��@��,&".�Z�����PU=_����DD��P��.��R�S�[�������������Z�z/�̙���93{���\�(Q���Rz�c���0a77�����x�㎺48Ȁ$��T���IS�����o>Ck5O�vm��)-��(����g��.)eff��#���c���������2_����<��968� L�(�^�y���a*�k/��U���p��p��qqp^`!�������k\���;�z��84�ZT�C񇫐����f����%@	�\[ߴ��M�zz�f������+�����0<��d��Э���|�"*}�m���aRE1d�w�����nxr�k_�>��d�W���A䅯����傞������zK�|�dA�(�dA��oco{��!JZ� d��A&���%���e_�g ��jj�jj�NvP�����T��j��������/Z�:��ڔ�����'�ŅtXeMP`M�������AiU
�T
�Lv����oӲF��j�Ѭę���85���D��22`BWm����$��R�c�^KA[h�ϡ|��U~�]^����P���JR�t���8f�غj�)���X�ҩnW��3|�M��y����7��HfSQ�����o�z6l�44֠���6=��c;�I-P�U'�j2������|#�:wu��j_����f���@�W�x��΅����41;�A�s5� S�x��H�"+'��?r�R��z���u���<�?����=�A�|��gG@�e�&����N�Ƈh���?{��k?'�����v|U
Cϕ�+�"�����58�c�X��Fp�|A��:�a2D��ԏ��G��B��#�WNOO�%�����|�|KB�/���ȣa\�����[Zh�Y5�I�5���a��2c�E��e���rV����3�ű��|��bvb�h��&�����Z����	�'���ֿ�"�IwW�Ъ� @���	>|�| ��Y���\�a��c�'gҹ*.���֖bT�,ϩ��0��̀8X�S�o�����j�:=��?�iJc��#��X/�-��,�װ��[{s=�̈́z�
���������M�$�%�S�1Q�7���Ǐ��K
�>r��2���"�32e�������֌+p�������7�2	�y]����KuJ�J>T"@�(�>䨘��F$�����
O�W_u=�-���q^�A����"gg��ow��l�&RI�+TX�7��K�A������}& ����"�ST������%��b9S���������G�{~^Z�9>p�B�Q��	 ����D��9??�S�a��"�{�4����̈́�,�b��}GH8`�t�
����)7讛KLL<��W2JW����"%��$�vz���GW6U�m�������(��~�e:	99ƿ��-h?1y� %�&�� �R����'��2�Scȍ�팁�b!e	�4
B642ZYz�_����i
��%�~�7SyuQ��7���`�~���%�=�F������}�&���*`�9�|����|#� ��M�&��>)F��r��m;$p)̀���2��;8���p����R6&T��ZĦ�y�q�%�(�Ȉ��D��\�"E!�� �(iyy	��������Rε�V�d�72�����Ы�)&���Ã&f ���o�>��y;L��"]}KK4�z~�ۑ0I�_�̎��~ �$7�F�T��X5����ԃ��t�ྫ������+Zy��ď@�����U��5E���̐�[kJ�}��rn��	����R�h��%��{�U/]�.j���\�16].��w�S��;���X7�1U��.9-yp��� S�L�ͅ�6��-()�TP� l�Y��uȯ_,P���~C��7S��''�%-�
��^�n�[��T"
VPT�}i,����Y��sT������T ?�DyErB�-�ZȘ�P�.:�/_�u/E��� ������S�\���(%��s�o�ao��Bg�h��@�'��������9�/�6>���]I���<���s�إ���0y5�u�L�[��O�1r����lܫ����*s \�
#�n6��e�y�Ԫ�
� �,M����9>�˳mh�S�+[Q�2�E,+Z�&�SӞ���<��rss)S3��]��o��.m�\ _�W!-#�x*�+Ha��I�H��}`��	8�<K��	[�y�qe's6�Kt0Ґw�L�����LOlf&%�q��d�m�EHD��x��%%�?FIM�����������]��k:���>��"Q>�߀�by}�`h����UuT�M��DB�6��S2��V�np�\TTT�?����>�#k���y�����k}��X�w��!+_����i{S�/�����U�(`��Q� �h��(���b3��̀s�~�l骋�85��hp{�����?U�ix�\�����B�%1 �М�	1�9qȶ� V��k�� ��mlء]Q�����E퍀K{��/M��q������}A��﩮��C����A�Z%T����Z0"]ӰAC��aqn��ֺ�Ճ���#�2��S�r����i�;2�xM��H�v���[�TD ��������;-�
�T��L늃<`H;�.el��4l>u.P��!$�ҶC_t�"�����@�(���y�©q�!��W����=�N%C�������@�wcB0�ɉ�"�����MR[� ~�� ��O���;8��|��I��"����QK+sl��3�w�چh1U���$�7�!�gw�^ɵ:[�d"��{����p�F��x����0i�!�a�s��������n"��.�.]��.G%���q�����]�o'��ˇ�]���G�B۠�$=;&=����yX
\�!�U?̓���������Ѣ�oz����J,#�!Ĩ?4d������[5��d~��g����}�m��W�����7���C̊����NW�S�{����Ǝ֎����6UC"�kh�g~"�#��	�E.��͈�b�jу�1�MA׏���M�h��%�$]##���!�q�Q���;^�h�Y��Y��3�$M�#�A�"�)��j;�����^�_�vQ�|�~�p}-Qpy��}���K��]��T؝���ٴ�rneF^"�A��|ù����?��eWc�;��u�2����y��YYY��qy�=�0��[_7\__�Ui[\$?888:=���<�ݦ�
X�l�_��M�]��7[��7���0S�q��Q�x�{vF/����"2���k-##��G�
���q�a��P�X������xy�jL�������`�Y��;���aM�����w}"�A������r�{��+t
)�U���ھ�#t�,̙&��^���T/�HdU�Q:*���@��@���'��4Ʋ��Ӻ�#��f��/��n.��/�C&�+���¾}��������Q�-d�l�>�7��'�����	T���Ʒ�F��B�HB�p[���p�Ğ��Y��|x0V��%���G�V�Pj-aL��'��K� (�� �Z[Y]�lN�|v4YV�f(G��GQ4��1AR���V��\�h����6~If�wd��o�ޔt;�,FL�����.Վ���=��]��|��3�#�3c��z�%_��H������~����W�	8�~������f,X]���˒�G��WUS=Of[�	``U�klH������M��>ⶼ;�I�5�p,�M��|�-�}�@�^ʓ_;���n(RR�g#��a�O106��g��=�yd d]i2�cዶv��["0��R��B�O+*��7-�����^���#Q&�pUK��!s�l�a��	�Gy��M�×�����Y�?4���m�N{���I��@c>0p��ѓ�DErw�ȈNM��A��_.�o�~HIҮ��:��iVY�ת���g/ B�M7h~0	�q�M=�� ���	j��S6/�1v50�v�Na�ЦٿH'��e�8L���*�F�;v�Fhzw{9V]&����O��׽i�E��Gq�'��]+���K1���^":���婼�X�/��th�����J���aO2X�M[y7M�w�A����Hnw{i$��T��.v�[A��4�z��F�ƾ���x00��qu������GO��AV1��G)墉:���������pED6�Խ���ͅ�#��� �h�n~���"��ӡ���P�R�J����9��C03-�3,Sᄬ�Ń��@���%�)if��a�Mx��i���g��$Kf��9��PPYM19l��^�'r�7����E��g�_�!D�;k�U�R%��6z4��6��po�]�=L�aK��f��s��lwO$��Mƀ_�"��+�w��=v�5�n$��m&� �����F�����Q�������XP��]V��q֊��l��%��l�Bv �ڼ�Q�����U^������9zHQ�ϊԘ��
�ZZZ��˳I{gY��^v����3(�h�@�s��Ku/20����#�9�<uVh��a˭�[7o�sm���$`�bz�2MSǙ8>o��M91ߥ���uo�$h1���,��_���& H���ȥ���^YS&��rx{Vn`qc0$?��&�@�GY��w�c�u�r��^A��U��
[��F��t�e���^=c��R=����'�����x1��Kpq�Ia�[�iԾ�\F��sN;�l�G�d���V�u|�ɵ�4�tJ'�[Ģ�WT���m5���8�u�4C9^��E�Q����gj\v�*H�]�*-�� ��wFJd�㯔�>�f���9�u�I��3:�g���Ζ������ci~k%������b�T_�8�������K&��#I��&�,��{{�뛛?f�)��o9r��B>��<U��EE��xZ����dh����^�ٿ�Dw�xd�qrrr�&5M��MTĵ8���裀��D�9rwG5߄�]��3�_ul>N6W���_���Pݐ�v�=S��R�'�G�3e�Fi�������*�!Q��ki�h^�������~�Z[���c��(�K�p�C6���sb�%�E٬,ܨti���ʷ5���F�r�+����.&v1�7�mޡ|K�����"q�oo�U7lZtX��� �%En����1�t}C��k~~>53��6gw�G��y�ݪcʢ3v��O�zQ���&���x�x�
�.����B��;�����c��V�ӯTx��W��6.R��Jά��Ɣ]�ؾHu��'���W	�s�'cg,$R�NZ�3,�h0��s�-����w��/�+�J�q��p�'�y���z��%�0Z`���Z�,3ā昴7�������Oe�Tt7o��G��V�q�J���2���7���ee���ճ.7�_����� gs�E����7�?��#B���q��-��	vJ�z�ԭ�F��҃�������=B�2Fon�?5ge���HL4xU�F"�a�{�LO�؂���3�<#��C�W%,�K��G��.o�����f��+�fJ��2Sk���πw���x��'�t?���ON�)l�xR-�����~�nל��C���~�Oc���k������N�SsM��pI֋6�M��Vw+�X�G�|j�wvȒ�y���T��K���z��K�?90����_����lI����ʥ:&ߏQF��T�[�7ܡ�D�>�g�^�&&&4t��O1��}G�������>�te�X�臐�����|"�d�����%�w�İ�@o�L7q�/�S%����ْaY<�O�}������~���"��7�z����TD�	���j��H�hS,����ˮS���3��8��Vb�o�H����X��5�P�O��<��z���m���h���r�����}���t�q�$]�K�&mU�������8��fgF�B.��k\W�-�=>����al[���g��L�Ǉ�~������d^tБ�[����}3��Z�+��M׼�>����-����Gi��[�S�m�x�^H��>�4��|�{��S�\ht3:))8��������a� �[���Q%m�P��V.���H�ׅ���OR��bݒ��1t�Fo�<&z�;ߝ2:��<n+�����u.���Na��M����}�!�n���ۻZ\\,�,�
��K��ϯ�)
�B�W�&�����`�77w�ϴ�=��6GggoH��lk�o�*͘w�5Q���j�ˆ�����co}g��ϣ��c�Y���mB�ˠLb�p#��j���ձ�\����������Zggg�_�q�LW�={��o�}S��������5�����T��ɓ'��Ъ��9E7���(���FEGkt:��t�U�:�/JJJB�/����ޮ��̈�KHH��1k|]���^����'9W�O�/6�1j'����T�*�Q�U;��IƋ���?�g��B��㣖��B����h����X~`h�%�ǰ��7���[�w�2������!r:���$<Xj-��QZ����K����=���Bc�H��n��Z�P�|�[��F�5�_���zܰ��Lƥ�޿k�����**8����w�k��ag�s�|N�_����^��������~j�M��AF� }Ť�5Z��Ns���Н�ҋ�����y���XF[999A�oq<A�w��y:�wwo�����^;h*���6++��d�|��#�wȆ��r��|�i��t@����c� �7���w�ߊ4J��qC�n�梊��*�+�����v�`}KH �z~���e��kE��y�����C���%EΒ�����)���^$M~k5���sO$���췐T׋� ������m6��3bA�?��&z8y�_~���FRh���	����!�iq��6�r���P%���h;7���f�;���;���~q}}J`_�HHBzz�S=>�<�ӽx���ٝ,������������n�C�7�w���㵑&���k�;������P���r���Iϩ��B����ӭ�嶧�S��Ħ+��-@��%kW8Y�g���W�,g;c� ��m����DS���J����涶�3^���jT�̨N����Ϡ��{��HI�&��3A!!#���*���O��d�����@�@�K����!%~kYP�V��7������ݦ��?��(�[W'gg;�P�Qh�K��"6�Oj��'rh��X...Tn��'��Ç�SG�w(k;;A�v[���3��О�Ga���o��7αY	�(����W���ݠ�_�������+��t���-��!�uG��{���՟&@�!l�gb �p4���We�:P���\}��pw�nhl���_g��Q�]����k��Lڳ��O�m$�M>�?͞9~��Z���R�F���K��	5m�[nY��
���71A�����'�^� �ǰ_n��y��l���]�!N4~�?~�_��R���]��v'ԋ����a���б1��$ev[
�WІ�@�1�ab`Ў� 

�������T=Mo/���Γ�Z.��Y4�C�wFs՚�j�(o!�fp�����s�~XT�'|s�o�v#NJyqqA�����'W���7r �K�Ϗ���
��-��#�-��)�0^
ll}5r��{�m	�r��>�y� �L�xޘ��Z�`�T��T2���a�DH(�5��z��<���Fs�rR��	�Lֺ�|׸g���܈�X)}�%$�=n���8�H��x�W*tw�}� �D�-�uf5��|5&=��T�ǻ��Z�n���%i��5d|�j���� %r�<n���xxy��V�o�ٵ ԕ�y"�F#�1?����C�B��;"���x���̇����̗Z<$g�XXh�#��/��Y�n�c��|�H��B�n���u��9fcy��6��R�Ku�^78*�~��,�U��2?E��"%Sÿ���z���a�l����;a�#R;��&�H<�"(�� �e�ڑһJ�ɲa&6a @�JdH��d`�������3��ۛ������<����S�}̓O�y ����<<��xLr�����jھ�@l����0.��T��!�:"�5 L�|���]x��W^^����U%�pe�]J��Ze:"zB������02>G�}eO9i�W��J���z��tk��g�1�t2�66��"ȣ xI���W'�|�4�<��W5!n����GO�kfx||���J��ut��29�r)��xew�&�A��/���ƏY�����NW[�3<�"ۧ�g�!��I7��!	��Ƭ�	�>�(��QdV�ٔ 4"���!#"������M���o,?����i-�a���!��~�[D��=]��!����t��@S��ii���1[��� (���PL|G��&���Gy'^=��d��=�{�Oͮq@T�Z����~�!#���0:6&aF.�:��؋�3X	4��Vհ��p�î��{[ �o[	H�ss��^gj)�*U���Qv�S�G�H�e4x�O���7�2@?��	�V�V}�;@�k�@��= �d��2��7f���R��7����;���DFb�|
���OቩXY_BD�OFZ�E<�'�jj�w	A�������x���d����h<ł����O�|�n��$Ϫܞ�%jܟ@� FFI�P��1��沲Hqq�H��ع*����6~���`��E�^^�i����a|�}qP��!�X���ó~�ѷ"���M�� dT�U����*|��B�ו'222؝���������P���F`
O��Qakph�d���.�ᖟyK�4?��;��~v��^WW����']QYY(k�k�)�N�R{ *�ONpf����=�*�2��!�%���tT�P@�M�^�q_I���zG�Q4a8��Zi]s���lc"�+��3�&�G�1�*|�1SaD��Ml(1g0�N�f666�9�I�RF��W���t�T4��f$��QL�tt�K�"���~�E@#���{!w��FQ@z�}���Є�K/mj�@�֒0Q��-��^������x�& ���ʆ�e���hh4666Yo�]u|�PR��<��\K��������uɾo3T$MܳЩHW�btLL�i �L��ϓ^�$^��ùZ6���N? ���D�H�����)r�
��Ĺh]5��bGG��������6 �輝x�oX/���I��O��ދ��¦�	�խ-��G�mFF�$`�^�4�p@5��zc�C,�P� tD�ꕿ�}7���c,O��'��gѮ���������9��F�vy@{�9@�%=#��۸ۺ�������Iv�4e]B�V�W�>��<��@Nj��prqi؎[-48��	�?E@{��z��j#n�dql�̻w9�c�) ��5�����K���_1@2 �>���"#!ed�[���g�<��u<T�A�h��H=<x��L����c��U8��z/��ʊ,H խ�4�����+ռw����Jv�߿g�JNJ�i�<37'7�Wk�������Ll�Y ����w�U@��6:�'dK\�𻨌�@5�
*b��h�D@�_.�gff^�MoF4+<�r�u�L�4��Dv�B`7�Z[[~�Ɗw��`��@ᙁ�����"#k%#S�$22::�X -�*DLr<�����c��*|����C��̡s��|�=wWL|����|����t��S	t�W��3����0)���w9�5C�9��ob"L���3a�u�KIKŌ�'uhzD�Sp��*ъ�^%&��0��iu��L��ٍL��A
A��҅�~k0d����g=ی݀�rV@�g�d�u6�u�� &y՟��P��^H_��U�)�1f����RN Ê�'*���v�k�V���=S��듍�X�La]Ȼ���F����i'�LAQmt�RY�U�'�d��cq���W�U[R�J�ÓX��(7�]�%�n��bg�j������5�-�[@,P�Iqw�Jc1
Y��G�!��ss1@-����kJ~cݶ{�� L���� s�iWʔ�OE�Ĥ��'�N=S^�C�	�Jԇ���E5[]Y
b���E5n+֔h�n:<��|E��W�ߤ����y�=-8�y�P��r��Tx
.k�dEԧŨ�y�8��ȵT����X5�_e1��v���K�)18���}}!�<��(�*����|���I��dde�������Us�{�Pseok���?�~�G��VO���̧�1*+*�Sy�mJu[:'�}���
>d�+�p�,���m��'1���������'�AbPM[�~���N$��������2�|�J�4��v@ܼ�����b�ۖK-�Yd�cc1W��r]�Qa�{31(�x�s��3fs5�b�����U��"W:TmTUT�J��,�
՘F,ٙ��`�iD=n��?���(��K�y�H��SV5U���0-8��UԾ���呔I�|�N�N�)sP��a-�_1i^�jjhh�<Ҭ,U/�@��\h������&��8�S�Q��r.�҅"��t+��J�<���X�@����d=�;	(���#�H�W +$PC��8� K��XT`��k
#~��O�@���p���y�tީ�N��<�t�ݙJz��̙��0��o:���i99�?������)�S�fBz:�z��f7'��6D��SD���%O�J����[@
�+�L��-����~@>Y�wvv�O���U~���C��P��x�Z�d��E�Fix` R�ŬE��@J،��9�$ H�8ދ3��M���/Ml�i�+gK&pY��<�X ���Gcw���z��RKH�p(&�K�L�����>gkjj*6)�E9��E�
�,,��ZwF�>nW���o���=O����k�}��611��מ��� �$��\������}r��?�\���v���Q��ŵ�?�&����a��&�!�i��?K-3��@����p8���g��>�8-y m��9m��Ag���R�)���u������;��#�*�	YiiaO�C�>z� �������6�_a<F���8D*4 #����짹U����@�-J��y[Ɔ�>"������B���#��]����6|ōG[Y�W�>��%ҙ3L艩<��H�]A�h���SS�e;�F�P���:zg���+�w�FG�1BJ_��hڬ	6���μҷ�(��A��p{; ��2%/|`D&�'��� `�h`P��%��Og�3�n�����O<ov�4t=h��Vd���f�#��,HG����xnL�������Z�P�h�\����,�>ޗJh�X���Ӹ�6��=EP�mPG�����aR`�~�Q�,1wxG_<�h3�ׯ_���r�뉢��� Zg�m�45�q����x�[���(�|�2:�����w��q?�)����#�JT��d�=�����;bl "OPHH��B���D-���D>>�0ɒ N� x�W֋�3*X'����5J����� �,��W!�5�T8i�lr�p^�0�cv�C�8��љz��ɒN��٭�~��/��[A���g�1I�nwm�ڬu趶?S�r���F����-�̓�?=mm_o\��q��]�:^��A��t�WQ'j3��[M$����w���|��:�񳜁HΝw�������P�G+��/��|�KE�����^{���cV�M<O�<ys�|`h�ޖ���8<�.�f���n�����p� ��4Qt�p~���SH5-1����	�F�������� G).��#�����F�|T��<OxH��k��7���/)�+Z�Z�Ko!��qiʃ;@KC5Š�c Z���>~$v�<��
�jv���c�V~��[{w�T%TU\��ZWX�ݖ��Ŝ���)P	<�ׁ	���h���U{�j>�:c=��ҡ 4ΜYe`(�kG�ʾ_�V+�8a�f^��o�BF����4��D'��,�B�lx �9��{������,&E	xu��GzLHjALt�/ �.�K�n����R�.�2���[WG���:�P�oHQQQ���1��̟���	h�,��|_��}b^Ml�5����CȤ�tt�;^��,�D=9!�P�CT�$n*L�lj���6@՜�k X�00X�#���j��xV2O���A�tq{��ـn��Mi����q��V?���b����_�!/�����wIo���h\���|�n�*޻�⬛�K��Ͳ�|�=�}u��.�'K������5�H�������Iks֭{�����I�j���-6'?�:�z,sȠD���
������GΌ��tF�LO�DH���/�z�%???,���b���dU��3=Ao.$��5�oX8"H;pzOd�Z�:Ma�g�0TdJkl��}��E�(��>Ǌt�J��S	ź<�*�Ű�����?'==����(BwGO�z׳�VL%xK��܌ML�T,8�-*?��`_��<�bⷍ�#k��Jl��,���<˧<��p	����.,�tv*�����Ơ���zk�.m9[%s�����Z�,��h�d..��3�׸���y
�=op:L� �����/�����t��^��+�=,ljj�zu�_e6&ig���%T7ZƱ���Y�"��߶P��6��!�B�x��29����s���rB��-&����n��n���ׇ�~�8Nx��֪PR�v&�啔�j���T'�~��mf�#x�%�#@�{s��?����
		�p�|c"Y�$�?ט9ɉ���[��c
����͙�3xx"�FIٌ�xx�)������r�B+���<#q^�*���?������#�bhci�`~{�h(1��e� a�m �
�.Zn�1���%}g�M�`�ndl�2,f�]�$���߇=Uq2�'u�jJC�rC̊g��D�����&���`�X�Nu�b����ȔU`ӵ;�n �	���ȓO���l���ڋ�=Y�̰P�x{�z����&;gWW�q���Í���\τ���Fi� �$Ň����'����	X(>�����j�@�ajYS�ov{q����\��֓���3DD�����f
�P��@����7ѥ477�U���J�c� �癹C� �d-�T�k<,�ϗ٬I~% `�Yz���@�ȱy��nҷV�4����y Fs�� Z��Ѧ��PȳIB*�'�P�|��:bL2"���$���~��(��˨�Go�.��C`��bgk�Bh�~�{��z� �C�^�1���OX���m����r�]u���8f��<y���k��嶤�Z@�)|N%jFH���SXdda�Ԓ/����;;%8��]��z�|a��*h���)]�0�̈́�m��ى�
�������F�bCR����|�в;� SS`[�Syu 8���F�G#��_xNY�����<E\]�I�z#$D�.Z=o���@�ŝ��ǪaR�
Cdh���[���B�[+b��sw����Ā����qh6{��
D�oh�: 9Uk@���[�~J�c[X��F��;+��R�+4a���?���ð>ב�D{��d�?:���f0%���1T?n 3�.�KU�dD�n2D�/on��� 9֜�FDD}����@D-����_��X�.%h��Z!���������G�f/?�{��'�]z���������Mqqߙ�mbu�������!ϳ
ǹ"/..�@�r>���6��;V���!��8�C+h�ȯ�Ȩ(�3�O��@\+t_^N�0[����Sj���ߝ#;9=����Y_@-��]�Q���:��t]�5��EĪ�j<�d�q>����]�L�8��+���2 �Ē��@ �2�:jj�ȸt�`0b�:����@h�/��e��(�r�C�	ڨi2#��B?��sU���Rx��O�W�;���i�Y��/�\`��=H_�9�R�wA�G
��Yt���a$\e��I�r4o���k�!N}��A��2e���@��z�&!a����\�M��F���*�#.N,�_����>��,=�����p��[=8��,p\T�>NjY�4_.�v�n���daH�?�MY� �=]N�(:Z߯��� Y���h� �bw8����[	��W���4����xW:�с7���H��!������w�+�a�����Bp�z@J�.4pN`c2�,�r�Z(}��V~xc�P{���ݦ�������t��N.�[�����<�6��7s�����
�8H;��|R�._�H��_���tr?X2�s��c���Z�4��W��,����z�H\��fʰQd�Io��ZN�/����_&�p��WQQ��QG|�T�g��pm[N[M�f<00 ��u>SiBuI����K�x�OT������Bm*b�̦���4�:44K�ru�]so"�~���i� d~7� 8�Qh�).��bJ�,�T�^�D��q_����o�C��{)��&���q�?Ť�)���i@%����X+533���.�˪�U��p��&	S
� ���xS�P(sYN����Tn*B���p���� q1�����|UT�мA��33� ��Q.�7�D���46ŝ� �4���5@��"B�� �	 �ށ�	�ޡ!z�<C��pgݮOr{�_�Z-4ġ4ZL��ʓ��� ���ֺ�4���0����1i��(<����q��Y�A���%��9r�js��/�hY�^������db Q���eC:Sa��_��!���ƭ,�OB"����
::���KR�zh�a���g+&��?��7N�W��zq|'zxZ~���o,cn����^9�'�j8S�]ߦ�s,��p��'[��4�y��9��On��AS�iKu6��3!�l���9NGI)�o�o����B�1V�����Z���f;%�m�G���D�T�j t��MZrrјP����Ύ$�E�����|���Nn�n8Ϗ�)���c�A(���<C>��c�Z�qĥ�p8�ݕ+Ѯ�������z�#[1���'J!�7J, #�bWn-�m�i�:�B��?�2ۧ��bP	X�V 5�`r����veA�pR�7+�����y_�P���آ��=LP=hM����0	��%����,���w;�ۃ����cK QB럌�ίw`
ź#�T+��8��;���q{}�kԟ?�L�ll�]N��g9%2�\�Q�-�"x���J3�\]�����\���j&��?���g�j���b�wGP�J{<Y�
�ٛ���#=���o� �Y{Nnn����Ϸ���i���y���Q��%�Ĥ��s��@~񥃔��0��8���<�l`��5n^���?�泘-���2^��>��ɺL�)�.C��Pz)�	0  �R�g��uӅ�h��p�"�pjVVVr�'~JƥG�2U�%�/�>qsq��"d���5���kkk��נ��z�UfԮ^'ɭ��=��������ӣ�~����V0^X`��@�gr��S�\=$�h˶���5�͜֋)@�v�I^�j��k�#�א �����?6	0Gb���K=q 0��C�9~��/���W�O��k������ .<�	�V1�yn�7�^�~m[a���vkdU��P�'mm"g���i�+++�D33$窔�&�����𶁹�TR�,�����ws(]w�/9�t'��v|N9�O�G���+�'�^���B��4�@q�$q�1ى����+��+3���k͟��C�B  ����4\�iD���j��+
Ί���`*|&���66�`���}�������	q���Vn��/<2i�%�u�tAYNc�uAۇx��7���ߔ�>��m�b�����F�ɐ���h��e>r����j���JW[��ȥ��Q�P���(���Q�l�E/�^�K䠵1iB^
��aL�w�|�|*T��F��L��)�)�g��\�~x�;�����+%\k�jӻS�1 ���b��<�s��U�n�w�r���K��#S�۾�'��m���XlO�sQQ}��.�X����m���ld{=>��3�����\�f+1��p�*�����
����<���JGGg�|��#��aw��&�uЉ��S���onn��Q҇�o�EQQ��lG��]�͚�%�����N�Zt��Co,��gJ0�^��;�m�ʖ��+���1�@s~�XX�^����C�ԙ��Y���R�'/�%$$���XDR�Rȧ��; A���`��.�}�kC����ӡ�W��4{{/|#��S���iҁ ]����p��ϰ?���l{�pg47뭪��Ϻ%Q�6�/}[��-�C�5����R��z��p�,��ݧ�-�/��f�/�P�_ e�k�����\�z���Xw�4 ��<�ԟ��Y���xa�{�d���5����+���{L���4đ��������q��4~&�iG1�M��kz���B5�����J6_jj���Dl{1轘�O�^�ے��; щ�bO��&逷��ƼAd���ϸ�.�g�$��_�J�grn;#w��X��^����Aʗ)����QV�����hn���+�u��B�����	��I+�Q��Fd�A@��3��7�S%�t:@$��Y�	0����s^o&[�O��3V�$ W�����eD�3g�&08���;z�����֖���~"�$D�Aƭ�NWH�䅃�|�ԕ��dal����?��+����Ȱ^lJD���� ԰�w|���7���(�@����t��K\�s���:"(>>�g�b��l��,	ԘՇ-�����`T����ҟ�6��������x3W�7�#-�C7���Cyi/���+����M)�#�C�������$_��*(`T7������ja��Wl*X��}�"�Њn��h���W��Ł�f������J���۟�d�VA�nO�R����H�s��c������~�����u�3-�'حvp�+�Thli���`�E��ҧ�hs'v���y�kEnrrrP�Жl��2���;�}ꌬ�]�RG����44Ϟ"��r�߬X���;�k���Sw(���2��\	���C���O
��]�Ɋ�ͪ8hVw�

�_��i�t��J'�aD���@�&W8�e�����^�].yIm�_�Y˕��bc�@���� �d�V��������`x��_��S��k�k�H��m}���LL��f�zy��Xߝ���]�{��s_��?�ۮ�N�*�(("���DBA���-17��z��`9��4Yy{@���tt��B��H Kv�|_���W,�L�ٕ|�m'qp*C5_����ŌMF�9�2�=�in�D��Ƃ�t�`�򑋋���f$PW�~����x���xaL��O�5��F'L�����EH��5������Myh
Ϛ�{ �#?oD�e� P>o���ȻǼ�C��!�鵇��{�����;����{��B��eK�k���A�޲g��*�-eoٮkvmQB\.�k�Ȋk������T����y�s�u��9�y���>翯5��]GE�j�Ꙭ�T���M�B���Gl� '�G'
~Z_�/
"ᖇݵ�60z4{�!0�)��sס{ ��8������.����9(x/���a����� �|38x�/��Cu��������YE�BW�EB�D�v�@@R2՞xQ�W�����,!��*�:000]�k�*aOq�]�=���
��TY�`��-LKc���*7aiShp01p��1����8���@�"��b�����==�%
������A::qެ���9�U늇�	W�	�Q��]ZT�����F��0Z6k�--v'��4=3z�{J����q�Ak]���k!�ׁ� "!��M.I_�x��x����+��6-5`@f��D������cN��OLN^�ї%w]S�AZFF�2�<Xx�A���O���'O�g����������=���C>���~�g[�X�N��A���	�z�Zv�5������_g�q2�B�Ѐ��}oo;�خ�ޒ�0�����^�)�9olx���������	)��N2�������޶�=�"2����}���OCF#�G��T�W¿#A���n�����U�Ԑ����G'^f`q�C]w�X����ۄx��2�Ɨ �p�	p��k�	�\!��cwѢ��W���}�,Jl�%�!�I�IH��ߟ����~��QQq�9��_�$D�����Z|��C��ҨB���)'�i�N݈Rhd�_X(p3�����Բ��J����;w���$j��_��x�˰�<����`iP>F#�穠 e``�+Sr�\�4U�����*7��c�R�aǲSs*lFk���f�]���e��UH��i���o��;����^��h��ŌS���w4�����U ���mAf�����廐d���V��'��o���!7͆O�E<�ǳ���FC���K�>�H~���P#�՟K��������P�MR11��,�TU���g�%{��;'���w\��q�$�#��ϡ�Z�s����A��C�<��!�M�����?��NT�yM'�j�_+�H.�+~���kԕ����5Y�n�A�_��Rr~T6���݆.�����o��\�2C��[}3�J�s��߿Ia�����&��c1W�Wi�<2���`F�S3�N������d�L<޳h(1����俑#X�b-���;����..."? w��BJз`���}u���*�N�b|z����9��� V�>@��43sfqE���i'`3=4�&Su�e�W+[ۧ���j�~�`�Jާd�k����T�sVFf�b���hfm�Y�tJJ
��*{����K���k��.,����.`�	!��J���{̬��e;�$�VT�sנK���q�b����׻�ty۾D��F�E�a�2{�ɻ`B�����O_}�ޮ
V/��Ą��2;(W��������]qTU�'�LE��N���V�%p
��qʾz���^��O	��U-�ͅ�/^6�7:�1��mu����e�P=3���6��[���N��YJ
o#.(��Ǐ\�Pʪq�~~*�9|�*$����~�B�Of�P"����=�H��`7	�߾��	}�]�Z�f��&g�s�����_z�Z399y��)����9�R�V��l�9�[EF�U�R����ssq��|�N��|,�h�e�/�p���z�*�d{;�TQ�joeO�W��$l��P�&�@/���gfƼ{�$x0�ry��/<��04�9:9�ZK=��a���mW�F�J�~�MJ�2��@�FG�)YAAav[������G��gj��4�s���̘�6�|�"���EG�Q�]��8\4��A��/�x࿭�����s�#���Qc�(�QM�'��Z[�����1������,hv�	���K��x�s����w����A�P0�T�0zll��,i�_�	D�˧̋�%Zq�"�����퇧�9	�*�
dKt�c:�Y�{��nnq��W�M\]/�gdXWwEn�m3������>'�.����Fz~z�8�h��#�1Xw��ݚ����g�(����R�"t��	&�/�>���9�����l��b��~8/�s�a�F���`����[��c|�Lt,"
	��bZ���٩�8zB�=G�5��w	9G���4;���M��`n��a"������f�d�:z{i����lI(���Z�qXDB���$��S�*��|d95o���8<�$|�X�Ei0e�	O�ហ�CB������@�Q��P��e�5�M�N�,���Z�[�˕F���(�]y-��&�F&�<5(l�I�BZJ󜂅�d�=��/��������X�E��X�N��P�w�~��J���@?0.��� ��8~TjR�524Lߊ/�T�Nޟ��6��\je8�@޶�;����@�`�h�b!o�1�#l�� �/�w�����NTN�*�]�7���B�������W�9�:�+8w���#�P�Sn@��/�w�0�c5�8�J�J�������W�7�g�W[|��7���t��c~�wUv�ڏ��?�w�؇�8j�o��p����-FA��J�f����b|��/���|\�O���@�? �W��m���e^�_�@�;�b�G���'ֱݦ���0G7u�vTZ�a,U��`�.D3�c;������~�HG�ev�Il�D�l��
����0�w�%p2}�ۭ���2/J����$�nzDfi�F��y�z�<��ۥ$��E�݄���CЀ��˾n��3_�p�Wn�o�����t�/�������gb&J�WS�W��򒘁V��pV� 	f�W���/�0K�P�"SX����MDx )\L���kf�o���S����Y:42�ݼ$q�Zp �[<��z��J�{bQzh����)�X�*�����qӜ���d����Ғ���e�!����9��L'�Q�b��5Q�ȱ/����L2��A���:��?_��?>Lg����S2�������=~���t����� N�����#���.����� yi�N��I��>ۤzGM�5w�,7��II����O�>B�D�K-S�j��*QwF�,��@r���ם[���o�~�!�I^ggg��W- td|�m|�UHH��������G�G�)��g$$��_�}1�L�W��֙�E�A��Z^ �	���ٍ�$�C	0Z(�Ũ���kB�nl�����&J'666��×*�_�>!����-]\b�P�R���E�2���^Cv#�����MN368�xJ�<���"��U��n!Ϙ�OU3��	"\?p��h��E�m"~���j�<T�7Ď�%�����2Ggf��vR��iO��dY���Ѱ��P�uj����}��F�S��=C]1��d[	���3-Q��jC.��yg��=�;x֋����拂��0��^(ҽ)�5�������>qRb����������3WlU�@�.Ňߧ£!a�b+sC��9����Ӊ
�;��k]��I�+S��<���*��K�S.?�r�!�++0g͑���(�}�9�	*H�@��$��&D�E��
գ0{L]S��	�EfP<���-(�@�'C!{あZ"n/�lF3����IW��y��:���}���]��*�x�j&�o�1g��|=��%����n�(��*>�0�OJ��XMZ��U�OyXօ�+ޟǜ}K֌�R���ܸ��,�r����ڿ"?�z����6k����@��Ch=�A��C���^0g�C���?���V':���fF��$#W\]C������8_ђT2�Z�f����W���/�)�K���񩸰��w��^!-���~�rb\��Oʻ����̫�N��;��ك��:��B��K]YhuK?Z�/_��Eگx��-h������.�r���;��
���K��I��\���7s$�D#O�,�yW(1�$�-ż��c�f�p4��ᕿIl�'om;Gd�T!������#�+�	2Z�60Lrp��C���
��s�	�gP'F=Lc^�uXx�gf[V}�
_�I}�,>G�+5�"t�7�F���k�@� ���M�.֏�ȓQ���.�³M9����y�ٺ��ɂ �(��K��3��}<�|e�L�d�1&��/�T"�z��8��@����u�r n���4���'X�`�7T��VP�����GȒH�S W&��m��Q�w��I�A��6os7~����C͐@�:��~
.^GWr�S�%�4�๺�l�Μ�o�d�����5�"B��F�y�~o�C~�jF�9m�6�3sN��^�Z�Dܽ|5�4:1�%(��st�,7�|@Bo�)�R��a)*� !b
1ue�}�h�`�h���#��ʡ	j9HQt��bܦ����;;&I�3�VGP#���nT4�8�+30r�,�!"y,���0���8��85���JTq�Z�������K?j
2��#����N����:���e6:��܋�����ou�l�3;e<��8y-����,�;�Nz;aZ~�g; =Z5q
�M*a/ )�4��2������x8���N��)��\ﮩ@���5�$<�n-������L۸Z4u֤/Z+(����u�b�|�}�|-%�m��V���#!�t�t�im�}���x8e24 �L.u�Id�\+�2���
3�OdA��rZj�M�֢y�~t>0��T	�FQԢ���ٽ��B��n_z(��P��v׉���y�b��3H�T3QG�Nvp�w{�Y���Py��͙�b�����0��m>����epҠH�˵��GrЎF��Æ��TfٰA�!/#����5-q�lQ����K,��R(O��G��|�V���[VFe��Mh���,c3����"Ϲ3��j�O��)bW�e����.�j��!C&<���f}G;����}�@���F�ԱL��@{����e���Zv�1]4�=ތõ�6;2lY����FY����;k���[j��A�A.��6n,hO
k�X��[I��+ق��6�[�5-<=0��C|H�7���ҹ0��&0Թ����H��������쯺���G�K�,<=?�oB�(�M�s�[�q�S���8^�L6z��>]%&;H39�ٺ&�͗��á.{!=%{߿CmV�
�ю�_B�G�L���{���������,]]�ǾM�e:��ƣ����̭Q�5���k�>>#cߞ�#-*UM�&#���[T�rppH���=s{��F
�A]�K�K�Z�!CO���<����w�ik���H���3�m���k�nʋW#�����aoO�K�K��V9��L���YS�c$vA_�}��H׎�S��F�����?:zc�� S���E��k��_l̏��.d��J*u��r���N�����M��ݓy�����x���V�_Ȟ��?���5��[=���5Ԭ��,¿L���>y�e�!�����R�/�M��v�����<�����-��͛�Wi׾�άsŲ���[�
�-�~R�2(�3�8.{?�}���o�_�-����=ſz�1���n���"k�J���`h�����6�Ot�q���a�>�@+I=^���Y}��1�L+��������J�w.�IZ
7=Q�+�kh�hl֭)l��@1�FGGW��X8�f�U2Oe���4)-/�����е�'
0t�/����yR
���h8�SY2=#%���BSWO����C��J�����x�&f攌��I��f>'�MuOO����v�n�Ӽ{���� S�fqH����/z0��6m&	5@q[�����Ɓ�SQQ���=l>�TU�vuU %�eQ�2���q?Iؔ�-@-����.��326����X��;II���#ͱS��y�=�P����hchj�8Q�a�7SO�wہ}G5�i��ΘB�).~g[.ֲw(��MT�::�mmmY]f!������G薻�j�����a�K���,~����w���X���Q3|"�r
���->9�u�Ew	0z<L�F���hUq������h�^Z�T_��#��鎬
g�\W�d��kq�;f"��h8�2� ������
���G��{�s���)���G=ۇ�Ѫ��e^g�V�"����MC�6\tN�l��+>Y��r�~,|�����Բn����S�m�S�<ڣ���3|�]�'˼��O�G��@#����)o㤾E��\�H<��Ul����B�.���8���@�����\�ZڦR�A�MKN~� �Q,Q�٤F��~x�~r9ڋ�����ى����s{��+d04Y��&鬯���0����e�5�v������{;G���M����y���B�];�w�f�V�\��$%�c�@��_g`�qtq�拾�*��H=�Uڻ�闣g'\e�F%����
�0���s�a�k�;£����'+qS=��������St�������Ɠs��Ϩ�����^4;iC��ڌ��հ͐̼� �&�lsB�b�Y�Z��Q��:`(�1������f��i�m����h�΂�/R����)�tV��{�@S�e����j?��>��ǙG�٨ �o�\E�DB��-�������`���# T��B�e����lΐ$dl��r3�XS���y�0ws�������2N-_�\� (�Ru���H�~��|�y���ɼh����R�:Ph&aZ�����b�Jۺ��H`T�y����.WA��3 m8�����Y�L\]��~Q-���ⓛqS��_���C]0d �(�5;�gb��6��	[���F��5�J�f���$O�<Y�A9q�#y��1TqS�`���I@ R��fXT��xGn4�q_��L�m�6x'\㠻����0�ge�$�CU]�C���Q��{����=v�.o\�9&�@�}�?��5�ߩo�>IV��,gt���#�L���Kg5W�ӻ9�0.+�
�z؟ܞ� �2�q�T��}�l� P&
fv�� 8ݡ-
��Gu]��d<+}	݊h�C�)h�{�$h�@�(`4M�{D��r[Z�l3}�=zE�/K]Wx�+�����������cb�2	j�j��P��1l�{ͱ����'(J~�I�ԔsppB��Gr�+E�X�����
~yT�Ogf�׷߾U��z+����ܾ������;�^t�0,�vp�(v����Z�0�x<	�"�v�tWε�0���9������7+���b^@żT���ɻ6�Ȭ�>�ey���>B��žmz>L��Q�/�b����c<���
,��i�.�$�66.������p"���Z|ʕz��0���

��g��.�V�:ۄ���<��j���w[�w?���;3s���/��]���d7���՘�Enk�{��e*��B�E�ylum?�iGk+�3����v���{=[�w?L<^S]]]o���Au]�}\�ԧ��p|QB�������^���{EB���y�C�W�XJsx8���Ji�1���T��R?WGG����~59>�?q�p�a�f4��ȥ1ћ��el���+sss�bcYu$3l�x7��f��m�������;.�.���H����R�NG�6Fj�$�������[x�m�>��H�|�p���t+W�K�	j��CP���nWE�-�|�. ^�����N�3צ�or�=��LӜ��Y��+E�z^�V��z��6tgw!�W������J� �4�9at�>ށfP�(F䤅�	�WY�H��}n9L��LCO/��5��(}�%C:��g��8������1�*g��M���<$s�-Q!,7�o+�)�=�PK   �cW���/�� Z� /   images/d0383ef8-9bda-42d2-801d-b77fe86508e2.png��US� ��%�[pw� �5�;��ap� �	n��;���������}����˩���>�j*��(�(   ]^N�  �  �#!�'bh� �T�JI��KIQ��9[�:X �9i�jz�K�ct�B9�nyg`q�,�"	2�Rp����+p9$�)�-��_b)���k=�zCéy��0U�����M>���ô�Æ���;9 �I�Z>�`�^��\i�s`���1 ��Y�"��ҥ�[��#w�U׺�o�11�S� )����G.�+�9R�Z'v��.�@+�R52���x��t4N�X�i�1`{\$����S���4.G��?�b,Wg6������"�c����Y5�G���Ǝ�g�8��1�����̖�?G��kk*�K+��T~M�N�U�7�'�5.�<��>0^d�tx�V�J#��C��}�2��s��I�a}�o~1>sǞV��(~1IUQ������	j���c�����4�|}�t��v��t�X��`�p���r��{A=�%9���A�������k�
;����մ�����gH����*3�9fL�1@D�K9 N�s`)c?�9,�Q�	��l�cU.��!�/�<t	
_��va8�x"qBTֹ�h�3�䮛X]) S�������T�h��oO\�Ŏ��9�H?�d�a�L�&�xu��}dް�Xp�_>G��)��h�o�Mu�c$W�ZB���C`�9P��]�a���]D��f1�C̮��$��B����n)-�>5D�&��#�K쨑� �J��!�F.I��i"�������,�oF�~9B�%����8�C�Yu� Ef��`��-⹠�#9��.ow֑"' b��nյ�cBQ���}[P�D�$�
��h�%�֪u�C[Z��;s��Y�AQ�,��ٴ#�#:�g�Ѹ��B�&�tB~4�X��\�ߜ͙8�������~,�}Y�Fu�+L "���c=�|0a�E@9�v� fo���k�y�T[c�A[���rmd����޵�?��4+!ULA��<�/��EBWaEbE�;��-�L4���/DΔLC�jJ>,�O�[)r�aS�m���k%%$�����UZ�rE�����_���l����1��:+��F6�}�m��|*��h��eB��ͨ��˸�ͷDI�Oۚ�]sZ�MG��_�'J� KMP�ܓ�9�7�7Q藤F��ָ�^���ߘ��Z9�ѕ���j��'��b�1�r{��M�MM�M�B�N
�s�%���*�uY�YE�Mk�������b����He�6�fN�N<}�}C�Y�0��y�xÈi�㉽x��x�x�y�m��Ŗ$���O-�W7+��Z�E{F{ z%��N��.@�7�i�>�
0�ա����ht2��&�l���{A��E4+�,O�9��M��K��s�ڴ�;�������V�N]	�
1:9�'t���u����8kV�J~_S%k�2Bg��wSs�OKū����<3M��d���	��ꑳ���<���Rx��dsu+��O--�zMgY�?��4D�D��֙�+���Yfd�F��o�G��֩ʑS����-���!g(g�������K5�W2m�&�.P��Ѕۙ�/�)����������ƶȑ�~�v��_��i�#�p�s�M�����*��y��Ʌ����f�W.mN��v~d0�Eb�F�����u������k��#�+��iv��j�J��C@����ˆ ����z���'7�2P=0-P��5���-6&>u�	�ktq�_���eFޗ�������eT�TsIK�Wg��6�Y"�"e��anR��b��(/�l ��������H/�Yj���q��8�T��~��`�d���0��$��l ��V>�Y�w�w�Ֆ�m�����:&��cpx7�e���|B�
aY��칺�������'dNdD��+Iޮdi�݄!3�����o۬+Ԅ��Ha����V�3��)�����%?�Т~)�9]�[8Y��-�}����#�"B&����q�+u:H�d�.)���q�X��eAO_��ZEm0p;���0��{���}�� ����v�BQ3=*��Į���X"/:31;�8��~�n����7��6�{(ͱ
Mr2�9&^��&�x��o�4Tm˺�8�~�B��L]Bm����¾*H��Ṿq�����ӗ��o�s���OO!�ê��K^N.�:{P���]�2�o���~?��@7���K,':kb[��Xj�2t�t�H�W������Ӽ��+���_2@���Lk���ĕ���U����8ue#ť�� ���˯����v�vUK��i�u�S��'��'b3�Sy��]h�E��ʃ�b��`����1��4h��׃]l�Y��v}MF��^!���Dyp�q�_z[:$�����������sY�JU.�%»�jre������a�4}��������Y����0;�I����\8htu�<C�ȵ��ө��r.$�q�'w:W��Щiã{u���t���������w��)���Q��w1�K�}+қ�q��X�yCaF�&R*������f���������|����K�'�{
�g�|��4�#��֠@�٠��X�g�����	:ֵ	ߖ�vVvޗ�-����;?r�:[���/����O�O�}�Ke	3���2A��v��wW��D��~��A)H�����? ������ge�pY����W���yX6��<XJ.
��3���.��u:�IF�����^��w]P�CjAg� ū�����2�=u�~�^��?����  �����m|���v���q�?~��������������c\8�@���W��Tfz���I��>f���tn�X�7�sO����훠�e���APn�u��[�sT\3�s��e��s��R����o>x����?��?��?���A-��uz�I-8V�����M��U�*��/!�7/��?�B����Bsڇ*kB��S�����Bwo	�gG���6�R������C0L����/����8?��v����2��fjU�s���b���}YU�������_��3��I��`�0����fnE�,C���M�{Y�<#RSM~�����B�|��O�m�������bu����c;���x���>�[N�V���׃G볯���榰ѳOUsZ�>+���i����zn�4��F���fͮ��U��c�[7����S���y����M���RGQH���d�̱,�Ie�������ᶵ����szm������������%�����������c���A����}O���ŏ�KϚƫ��'����Z�U�p��j�P[c{s��1�y37U
>�G0Q^P�^�?�>X�(�>��V�֕h��*��!�&폹����O��ſ�K�k��tT��|����;��Ck��e<�Ҵu�A�SlF���-�����'�d$/�l���=�Z���ׁ�p�/Ϫ��ju���(jۯ/���έ��0(p� ���@��$!;�P"����^G�#w@I:gV?6!��"���_0rBFKK�`�R�e��h��+����O�p���D6$J���*�Yb�.L�vq���@X9��U��)h(bo��&�7�.���h���o��g'I �����W~�	���p������n�^�ˎ����xȅ�o;�GO��8�k��8�u"B�rC��]�o��t�A^�ܓ���e==�sXD̦�˭�G�q�o��Y`�����(��an�JiBi�~�n���-l�J1Z��'��шp�t;�@��m �R-E~Ҋ@������I]1��{2�Ñg���pB�(ٿa�+u����\�G�������_]�z*j�.ʙ�//����id|,~��X�/9�v*.����G��xױ�tC:��Qj��C���v��`Hq�Tc���8 �)�g�����X;��)9��������YzRl4N�֜&���x�t���_'���X1�!�ϟ�5gn�io�,�M�c[&b2�O W�ݬ_4��k��7�';f�s}���a�o�>�b��l�dnAW��WW�||��n7֢W��&Y�7[D�\t,�lf����ڻߺUI�H_��	M����k��͍�M;�R'��x� eV<�S1�V�׺����amE��tc[=o3&�OMIA-�s�$��,�W���?�$B^��o�5�*XH������ ��3��w�C-2
j��r#]��s�0�W�m hX�	F�'�}�]�M��U$0`+�
���l`Ϧ�W؃�	�#r�&k��En����_5�yfr�xx��Y��n����Luq5Zol,-�L� ��m����)m%�KuH��6*[_U^�F�Ñ�c�ֈ����r��E�s��s�R`�緍<w_@��ًd08�5��sp�@�V�� �8@)5����m0&�wJ6��{#��\�o�/}����9�ڝ;��n�{o���U]���(��)�d_[�&�҂��/�o�a	�m�0<�8�#��z�Y&���xW�{�ޒ�k��A����ԑ���d���R�=�����/p!v0Z�`�`�AGH-_"��H\F�pF��3��Q��d��}�ë���E�3�z�����̉�i���O�����A7� qVT��*���h�;���71�a��u����.ͽ9]'X7.Ҩ�,�sԱ!�]b�f���`v՝��Y�;~����xK��;2�@Dݠ��"�ډ'�[�Gdg�9�5#�QwZ:����#	g@���S0c=p��ƥ =�/��0�I�]]�@�/l�5-�~-,������%=aD���>3}*�#&�YYp��������X��GA�š,�1<r��K�n~a_Ȧhk�q}P���a	�^|��,�;����	j4+6z�r�~:��FG����>����}����yI'�Ŭ����}�[�rJ��4�Z���$�%.7*��P�H(T�r9	�Y�-���p����L;�&�-Ҫ0�.�5����ͯ�P���,'�>/�Opx�uHj���r����9��Žgh�-��*G|�������Rr�w�+��ɉ�����)�?���]5�1�F(�(�Tg}�$��/>�7t�'dx�|�_f#��~��ԅp�M1�����d#+E�f(ӬG�;[�@��@+?9��!�j�6��J֪�9_\��4Vl�TM�!ٗ+�[(�� �< �$����� ���@�[�.�њe~��}-�O_�`�&iN�|��x���� �+S�M��<>ᚙ�J9iF�;YY���0�F�J��.�e�Ss�t�L`����D؆z:hp
qZ[�����Yr���)��d2XI�TI�I��8815ƓY 	 �d+� u6l����s��ޞl�������%�~������f�@�~BRD�xw�\g�/�g�u���CӪ��m?Ӑb�1X���R׾�ݍ��YؼD��8�N e�����wtu9�	!  �fzT�֢nܕ�b2�\܃�kNGB�������	qu|�� ���):�����I�yX�a�͹����_�D{x%7�pV�,G�� �O�f���JɁ�o72��(��?��#�{*\��ϏHICZ7a`r��D�%�.���I#&�5}AуGgv�<����އ~������e�a]J�f���n�E{߇*��׉���(�����Bm�m����:AXs( �9Gv�-6g���7���q&�u�E�CqWk��Z=�pz��B�CHO�*wCm�s7��Gpn"X�[�F5���[�-;����pF�e�%gU��g[c"J��������Z�;���]�YN`Xr��	�l�^h�p�pt�ԧ�o����	�js{��πY��).�u�zv�o��P�I�~��=m�o���4X�:�o�T�[��W�B��Z��LΚ�ha0PS�Rp�I��7bv
��5�ʿ�@p�� ��r"��C�1�$44�)�涷Մ�ov~�?񈊞����`��/��U.��Ȅ�--Y񻄍��I2+�{rGF�K�W�G|�8���E[%��s�%T�6�(r�賟9�,_F޸X��<ja\�Ҁ��h�T *��@	�em�q8ԁb
�/�$����2�ef�O�O�>���"|�~�(�M[��緐��f��3�M���d!3��_���ȾfԌL����2�ly7'���u��� ������*�����68k�Q��]/�)�1pW[�i�/��ʻ�?2:.]wV�:�Y��H N�b;��Fh�t�м��5F?ZC
�_j>��� �6|��	��s���̄�i�j*V��q�H�:ʝF�nY����<�����+?[�|Ej����~�7�9��ax&"��<���k&4��v�x�����dO115#"2bn�w��u �t����{��8��l���:�yU �z?p�#aa���(K R:�VtLA쮤8�p�4�q`�ܺDm����`������J*=�xx�=��>��t66���B�94��N����w�S&|�9Y�]%��;�˯%�})vd�#�v��^�#��"��G�߳7ۣ��u����>����v,�����'�4��8���o�~�Px�G;�F5�[�K����z���4�K��b�Qc�:v�`58��x�rU~G��g�҂qdw�Nm�A����qX"4��`�W�m��� 8 (+{�T�%���&24�L,�J�J*\l_.���c��k�ڇW�J���'v��n����9��wN'�.08�H������{� �c�j���JQ�����V�Δv%�	m��,�=v��u-�py͟��R��/f�1���-K��W�@�Q1���㯜���4e
�gE�3�f-u�:���d�vڡM�����Ґ)�#&,#`Xu(he�@�qV��9��*�f�������!�%��}�<�gr6�E���6WA$�0ʁ��d��j��Jʮwk�a����0a�1L~�\�����`��Q� ĲA�n���G�����<Bp5��H�H
	 �r��U�v�z��8X�h^�,�m9��U=Q�0�ae��!d.��-[����	P+m(��ƶh`J��i\��m�x��ro��f6+�����ٺ�?~���|� Ks$����l���t��HP���3ݝy��^o�x�v��ǧ5��Bo<��oJҗ����< N��V�{�-V�M�6����1�5}?��$��rҖ�-���<�S��ݦ�~x��j�#�;��p�i��z��|p����V����
?,���Ԍ�N8a���uQGXD�NB�[h�x��ҞMV(������iSC1ҹ�?9dG�b��Z^��Q�?=�#�p�3��ȓ)��r8zn���1:��������K��\�^�<����U��y  ����A��{-�h�D��/��̐ڱ�N�o����CpT�H��܎Ћ��>�/E^]ܭj����.��S�x}l����i.nfj��Z_��U�'e�~;�����T�#M���А� `��"�#����b�UI�%Õr��+D��V
�[�o�� %�}�F���ź�KIӘE�FHl8��g�Q�W���I6
�mtyNӃ=�������5j��7tt-0��d����)����L�p����Z+�B�.5h���oPz�Q�Ų!�FyJ��ɦp�긣��ET*����
u�z8�	��m�3��:V-Bq��'|��4���}��R��-��nA�|[�Sd+cZ�YR��T�rT��b[]��Z�BXo�2��>�#5�)��pV�;Qs�S��t�ZEia!�Um|��I���{�g[�b���Z��t9{cZ���"�a���Cс�	 ����L(*:֝˹�����^B)}�+�G,�������V��߁�5�s�h�٤���'��"Ŝ=p�FA\V��Xw�/��[е�m�S�.�r�����pARq^rG^$[p���
�c����EG�O'G~�����;���r���T]�M��K9�hǻ�-��z��k�Fhq�˨*����~�KJ���7�_����$�-�	�K��	�F� ���&�4���Q�҉�{��쎟B�� ��Y׊��R
�o�����3�缝�e�ٲa�c��r\�u>y��~�#��㛻b��X=�B�-hol�5�u$�1vh�۝�������o��vT�Δfj��*y��@{T5M�O�O�鯰�r7w�JN��1���Ek�E��쯽��+�[{��)��$��+����h������0�f��I{���:�^<�J��L�~�Z���G�����(:�(׻���9�6�a��T��+��]���hϠ,�{� �<�p9$�Dˡ!�pzE�b�S�����z�&^�8�����o��N���߿�"�m�g!pCH��C�"�����&ЕylF@���2"�	���վ�y��<�	Ġ�&�?�;�Tm��t��c�;-UES��K�&��8� �@�;��#�N'���}�"R��CKV���h�"�6�����a�N%d�\x~�6�#��^n�tpR�z`:�a�C���n��X����f��N+��д��0��̀�� t4�b��eW�(�h=h�+�iX�`$"<n��[r� ~��[�^��Z�I�+�1:�kV���B�0��e��·�n^m~&r�G���
֥Ner\�s�W��Dl�p�|�!�fp߬Iq�z���Iw��a�2�!д3=���� a=Q93�Z4'sA=�e��0܊i~���Ȥ����np[>�rK�����a�J��M�|R*�E`� ~�ia��Jg�h�.� {Op� HٗA��a�C6Y%�`z`Q>��8��MM/����t���˞1�͎�l��u��گD���AI����z:h�J@؝�]�z�*^8:%ā�*$�`QN�k�_v�Cgr�ï����٤��{�6w� W%�ڬ��?fΟ:x�g��mW?�r�qf�i���i����%:}���ѝ��(0Q:�_�6:���y�%���������(��|;oo˪�V
�����ϒ�T��M+ϷԛS̥CtCP���}sޚ������I*��nu8>轧�}���#�?pX� \@B:G��w�:Y4�[��d^o�U��Y?�7�����u���I���y��ݽW�}����e�)R\�ꌹ,�\��"|q��S"?4������ڡ_㪂E�	Ot%N�[�� ��$-�V���B��=���ia�<sDv���Q�G���� `^Q:�Z��Pa+8�0`S��R����
��UH%&cИ�f)�ɴj�j�u��̿�f��E$��끲��\s�X���x-A#ղ6�7���F8]S�DWHt�;�� �ս-nk�)�Ԝ~^��%b�/|�!�Rt��D|1AF�z�~����PE[kk>O���`���Ւ؊��(#��u�l��ӓ��z��;*��6�(��Q� \�nX�u=��E���PZ��U����$m8�:���-x~�<����w� �ASض��x,&����ـ`�>`�fp%/��\蘊Ԟ�V����F�|�@u�4�d58�Ô�g٨mc�o��e,G��L�u>��<��V�P����t�I��8"�U�wj=�k��&�i����\����O�s.=>�����G1�K��2�Dq\ė�2$bv���I��`5��*�'���:�:��L>�� @�L.�=�"��y�4["��O!s�|��'X�� �A3������p�m����Ī��U���/�?w���W�����r!��\�뼐�H<��@u���\�qa�iD̶ڡc&,my���A��}
]�kA"y�̴Y%Y� ��5'�`�
x.9���s4yK�P�����L���N_��J���w�n��K����:Q����?�jP���Ѧ窭�X�Mnk~^����?��������]#cgYT\,�Т����ѱ��y���+�w��Sy=W���^d/�����ۏ�'E�3�g�O3�S�|	�3Ϻ��,�5:V%x�2xS@��!p	9ص���1H �M�J���Pe̔�V�e�'�9��9�,,��AJ�v���&#3��Qjy�E_�Չ�2>���`�F�����} y\�X��f���g�)VH���B�;|�mVm����͝�&��SlRc02�ez���-�J�9Vv�x�P/���6�R7�=H��쌊�gS|ggZ)���׺oe���g���!i ep�<'�o��[ ��`�j8��X"j0�2�!5�,[l��DB��^�r����%X�6o̒����л�A�-�y������Y�|zK�_o.�p�Ư2��d넧;��W#����*�H�$��je�e߲m�\���ص7�nߠ�w���
`��tS�w����Eτ������5�b��
~�w��5�i���Űb2P�w4�e�F �O.��LX#���� ����������6<�L�
�ow,A��B�#4��4�� cш+*3b|��O�h�i����	����c���o'�L �׸�݁.!��
�ώ�'ľ��k+����	�R�)�HP�JD�=?����������K�O���T�f�w�0�[��}녎rK�m���ūJ�%��l����:.�Ɏ~�}<�S���z�r޴�v���@W'ix��v�.���{޵_nA_RӾ�W���Ɩ��&O�����{a轿��Ä8���3i<���]��me�>�pP�Kq">�y%���_����wy�L�8�{�:޹��yu�ۧb�#4�x)����� P�Q)��Y��w�7��]���[�H��+���z���);�Ԯ�̚�#����J�%Sԇ��W�[�x<$&�j�a��#䁑���h�v"1�sQ[d÷�PC�^�P�n�BX��X�!��:��h;K��'ѷ֠��=�=�7\���}��wƤ�{��ʞ�G}s�����б�g3tF�_�V¦CE�!�-��`.����|Ū��P��\����ʱ���ĺa�#e�Jɗ}2a�L0�[p��C�Fr3���}UNLb���Φ��IgGg=�>9m�1���IРϮա�XK�D}�^"�=L5h`���� biWOhG��U��զ$�נl���_�6���A>�Yu/u�ꠓ��l��t������#�j���0VE����u&0��37�#�����Y cC]�-����t�9�I����}���W2�6�KB\�I��}:��R䇛S�#6RO�m�<�4)\E���͔9����ȏ�k���]���k��m�S�A�X�e�=>u/ 5�ah�i^*eAy�b��Yq��Uڿ�|����%@s�lD������;4F [=����E�1Y����J|�M��gEv�N�]����/�x	:�����W�X4���q��n𿍝�����Ӕ��:U�o���t�a�����?���7y�B��L�����I̢��]�q75s��X ���/��_O� �{M�Th��?�n�ݘ�߇�Od�z�_��-���7�b�H�� 0��=����i+x
�d����m$�aیe��hN:�H�h)��+��ʪt���ğ�fIȷo�ˤ�e����5�Պ6x��g�O�	&���V�;QM4�99
̨�Ϋ؈80c�.�U&Zt�wm�������;�bNJ!����f��Դ�� B�d��KD4�>�/١Z�*` X.Wզ�S��Ͼ�Xŉ,��i�a> �|.͹���ְ����Qʯ��,����+��gF��G��9Vb����e]&RY+l�<~CB�+bݮ�'���nǙ��ř�g�{�h��%"�&���\[J����I���.�D�M�gJ�IDৎ�L�"�G&��8B��-��\�P��b@S�.`wӊ�D�&�KHõ!%�ن]�*�c�����'-�lu+bww�E��U�V�!�-�A�EW"��&?{�x����Ռ	j�h�h���+���'$�F�r�QB+#�X���'@w����;�}w�6Afx�$��]8YY�a��QO�����P,vw�l�.�9R�b7'��K���Ӟ{���V�E�4�@� O����4=��3��)|��#O��cNN�-�"�fi9p�}b�>�i�y�g!�%�(|����3���=Z��ƥh��&�ɑ�.+KZߋ���
q��|���D���2�h"�ӣ{�_��F�~�����S0����<(S [a+%�����2��U�z�I���`�X�G�� ���1�:��L�\��^��>J	-@�i�
�U2_��y_٦�˚K� :���&)�J���������I��#:ԯۚ��>4����{F�Wm�?@�A�g��w��@+83E�Ɗ�0�&n�gG���	���6Vf�_��c�;��ho�T�Y���=t�z�ӡ���P�*��Ç1�Y|������)���T��,�-���F��͠�R�E��)+�D��x�*��}�v�|ߞU��\=�)���yÎ�w��k�{G��9N����6?����v�Q���AA���,�:�NB���,�L�]Pؘmg��4���TP�yc`?h�#e2��DS�r?��<�N�F�t���F-�:(��� u�t��jKT�����vw<s��/��߻�"��|���}��� ��҇�@/Q�9�3���z��P*� �ݧ�-�d��P�Z��a�R�])��0�}|��K�����H	��ƿu��<D6#~��*���#��Ū���
z�������R#u������^��LC#�U�S����~�����l��N!��Y�~x��>�Va_baa�?H��s��ǳccV�ЅȣǞ䩠{w���'��>܀#:�6��m��%�QS������[&Q�%��W�"�y�y��a��=T©�ѩ�`�e5X'���$� �>��Fq���0�ҳ�"op��58`��������*��2����Q�N=����t7	���\Ao��Q�
�(қ2�}	�"#oD6�_1,(���0Nv�� }=B[{��x,n�fb@JJxcn�m�ݰ�SG�f]A�g�E*�=����������p҈䵞��� L�+
A��L:�t�)��8e�B�� (��]fg��}�̔�hfzEmFuy��6�Ve�R�_1�,��OSsj�a�@lՇ,�o�5�g��S9kڂ]Y��0��B����X�>>�^��w�I����oJY�*�����6����N_�e��y޺��En�-��r>����n���̖E����U�D�w_��D�P|o� _D�nh_��y|���<5�Ji������!�7t-_O;;�e5(�@_�>���J�|����% � :��.�8M@�\��"������ja,���ڄ�����vT�*��&��o*�_�Mi����w���6�����^�q4`���"t?�b�<�ã u�m:��:�ѓT�T ��`�x����vv4;A_�}vSؿ�6�\\�%7��s��>Wr}1L�i�E�����&�ȍ�X�Е+��;�ƍa�ݧWԏ�*mh�UR��܍+~���%b�9�Ҥ�<���,�����T��,ZcuP���"ľގcO?����]�=�b��^pՆ�뿮���Wt4�Ns	�Q{T��?{e'U�H^��t`2��{��r�����fzT���D��hUm���3`i��jQ�v7����|��U��~_�� �y�������Xգ �;����s4 �k��⥄����������ӈ��ٴ��%z�4�Et��7l�O��p�n]bw�g��;_eMy�Ţ�9R��?l�Y|3i$ϝ1�.��r��q�4m�[�ʅ�����	��>xʁ�2��jo�X	��Ӻ�>)���P*���?53)���}FY�<�@��G��BF�s�p9����:d��1�[%�P[F��X��-��ך���C�uX���Ml�/�m�"BC�9�@��Yɒ aLO����E�R���}�HZ��?t�r��({2�y��\T�������� m_���q���}@����&=���Wk��2\Mަ���㓏'a�� [�=��[���;s��m��Ҵ���*p��s��a/S/<����B\��q:3��aMk���VVou���m½RB%���E�N��Å�>K,�Z%z�P���/���x(�����<k�};/�p���N�&�����*4,
���Ac$+f�5)�YG�Pn[�J2��t�F���A����6'�S��6���.���j�j܈IG�3���ʒ��Enc��Ot�gC~J���~.|���Np��C$�(��nG�0������u9ši
�.��my���u5yO��2������rul�,&���:�1uI�x���H�j�8J�붆6����Z`P��Af_Xr���98]U$�����o�`x:{�a���9C� �n��?T�iD�s�fʓ��!��yd��H7O�[e(������H>Հ�:�=mb��>s%ry��qݣna8$`��"MN~
'�tx��k"$Ǎ�x�n��8�E4�E?;<�s���&�p���E�0���='�η@��lH`��nn���E򪭗To6^����(������*��Kه{M9�Q%q�ȼ@���9��뀣[H��/]Í �{o�(�60F�w�0S������ㅦ�͑�W��i�gI�E�p�n��yA_K� �-��xW=�3��^�J^���R!#�\���R;����0�������"�H�g�B4�{�۳{��䢠q��E��8�E�cML���-s��6����~�2v��OWs<�ߨ������e�0����JH��5Ra���՚:�g��3��m���t)d�f���2'�����8W� {,� HH�`�̬��l��α�!W7n(7U�Z���L1<P�#�V��v�Y��e�e9<�j�^��A���y�B6��t6�E��
�R=#���1��;��o���3�"Iwh!V�}���_��x�C�q�m�Ex�p����#9`�.��"��F�`��?L����X�θ2MY<F/D�o�>���1��1���t1�����>�m����q��%\.����(�f��N�₆���~��ܦ�I" '�a��W�k��	iO4����3Q(@�	{ݼ4�el���c�ܦ� ��^w����[�ȕ�yZ���w�	���HԴ(���Iu�	NI*I�
PZo�R]kub�)W|f@с̉O�MTQ��%�s�ʇ�[ޫY�m3�Ŝ¤\��	����l��<����7�Yy:������j�N��~�ӓ�͵4	���C�8y����$�����;�����A��=�����ōx?���=����-����du�X�B�y����?֪&�=nӺm������f��_��M5�A��]P��~�A��G��%[]��Hi.yq���%�"��ȷТ� �;f��^��c�U+y13�_���5Ƽ��*���Z��V�,��a5�K
N�<��Vӎ5�7^�HWG&���>�%F���� �~J�f�wyP�!� B���R�H����]�taRF\�+w6`ఊh��໨yI��T��ZѬ�� ǘ��\j�.7xD\:srK��	X"x#�Bs?"*�x��.b�6Z�r�Oc�sD%#i�	������'^�t��xQC�B2	��x����%VD�Ab��X{p�L���Ԕ�R6ױa��.dvےChLj`��҅AR^QRi����p)\ό�9U����u	���G�����u�s&�lq�� qf*	(1w�pJ����!�M��T�$�~j�f8���T���Xc�hƢ���f�w{hڐs��1��OR)g
�Z��-�i.�u���$"�yS��Ɛ@�_�H�ŞnS�ƄB�&�c�f���2�r`qʍ��/�����?�v��Eh��C<u����a��Quv�݉KL����Z��a��P�M��!E����>��.K$ծ�F.o0�b59x�]�H�n�mb{H�1���<]�r�0�K��"�v�Mt�w߼���������2 �q^VO2ҍ�RƧ�������7K�|_t�{�#����!Ԃ��c�����.�4W�:� ��� 9��N�Ձr+]*N��yri��
N�:��Qq#
.$�ᝍ�Nή,Yd�E�g�!���=�Pq�K1=�ti�6��熀H���0֥��$��C��"������K�/�RO� S@��(f�  K��Dx�c�z}=\����4��5Y��T#�F3Y�mbb,ͨc������z:	d�jמw��,���Y	��6�P8��ѣ���r�AN��Bw9�H$�GH�z�m���tH����U�A�η���0&�r��o�%M؟��v�"�]sܲ�C�U&3��pcl��h�	W�(�7�K����&�200�p*�Z~e͘Ac�����ᜑ}�C~�%B��x���ԫyu��Y�S�Sa���ܪ���s'P��s!�mU��^�:���J�v�@�چ��i���z�D{~��P�pC ���Ȓ��P?�PZ����q�B���*�m�4���;U�Ǌ����i�V�5M�ѽ����T���,S��ړp�ٹȿ��f��=ը����DZ;or$}��w����w@�e��X �+�P�_�L�Y���+8������xm+���N���i�/�95��1rM�?:$˖�T��d�B�L��r-@k�t-[n���lZ3v�g5�����S�K�յ�N��险����ޡ	5#�fM�*�J�����( ��Yp����rlr&T~����<?2r�}ݏ^�xq�f}s���Ң����*�cv��N��� �.��,C�è@�~��p,d�_���]x#��h�~[T�u�^e�iq�h��߀@���u�B�k�� ����Ј��P9�)�	rV�λ�>���V��'}�W����?:2(���C��|.�x�7���&c�v�õYH����������5�t&�҇m�&7�ň'*�*�eD�,�ދ�.9�wp�^U�]I��K�����NˋjN9�������6�@ ��c��m��i���|+В�]�������8�z�f��(��6�1+�C��y������ߟ���C�����'�H��$�C��q!L��,ʹ�Y�FtU-���F�#�2y�sv��KAtiw�L��_�Y�b��^9����[oQ��D�r��Zt4wk�b h�u�ޭ
{b�e����#|^�du:7�r�P���DZ��n��GߠAH�ѪHa�����r��Ar�Tk�� i� �a5� �����|.�Y��Ω�=���n��~@����N��z\�]_\�ɛ(Z_��:p���۰(åX���sY�9ׇَwC��L��c��%���b����W���hֵ/�յO��~d������1�<׷�s��=�z1N�ғ��v�@�m�-�����},��{���O��º��}Wf��Xo�L ^h_Ϯ��4���s�yW�"�[�L:�	�9V	D�zq���P����1	�\/�����b�R�"'>15�z� ����T��jǟE��.9	�I["H����Vw��hw��pв*4�oϔٛP:�o�.K=��'�45H�r�mT�柛���ƉT�"\���S�Q,�e���9��M�U#�oʎ!���f�&#�0�Y{g찋��i���@�89�A���"	��?�7�0'r��5�������?zq!@m  �}�4�<����`@D��@�;��1kC���*T3�����&�mM�����n����i*6�ؽz�r��_���#��kf-ֱ�P��]L�l�0#S��j�:屶&�b��bB��:�p��F� 5�	�Ҭ��B��Ƚ[k�(`,�?�b�:	Vaaw<�X�pS�ʕ+�6B30ҳ��=��VK���P��>��';�>�E���5+cg�/b{��͘t�^�0@��2Qf��2��Y�u3[Uؒ���z�h��@�Z>�ܞV7��\���j��\���s��0\�Cc�5�����n!Lυ@+�m�\����U9��aO��(u���՛��{���=ۤ/�m�>{���_zq��K/�Mm�h�L�.���z�X��l��-L������j-�'u:V����ӭ��_��{WG��e��~��?�Ý��;��TU;A�/�tҋX��J,�츜�~TP�M��U/��)�[4�Wǡ�!Y>A�G�u(�ߨ���3��(�	2(ǍC�R婢���K�+,A	'�~$g�Q1w]z�^5b�)6�֌��6}�\_D��{����f]ןw�8	��.��o�-k���t���erh�����{�a�����]�=�`"���&��Qˇ�~59�m��^��^��q�+X�b���]u�˖BP����+$F�*���rzw�5�TO�j��M��O�]]CS�!�CLL���$}�n�Nni��E�D�[*��8�l��b0N�)f���U]v`���垚��r0�%���p�  ��D�f(��55�%X�}�ݪ�/���ZS
:�������ޥ�9ұ=��ݸ���q��Ņ5��ID���ؼB�#*2����#mN�7�X�� � \4��u�o���I[CM(l��q��CwܕF����}�u��m��H[lS�&��� �ꚇ<���Y��;������
�T0Gp��/τ�JЇk��r�M���.Sf��6�eKI�E�"2�2����yפq:��"���E�G
��U$���� O���"�2�X#��B��&�� �8/�H���4X�@-q�_�T�0�f9�V��>�������y�_�:?w�ڣ�;4�e2�:������0s��_I�ź�����3g���0�,.��'����/������ps[ Vs�[e ȵЦ�ǩ��&(LЍ��u��U_]�O'���ban���������g?����c7r�����]��Թw/�5ok*'��:&�H� 9�S�"_�|9֮��� ��4v��K�8��[��k�s��N����#���ɓ/{���$�fG/���Y2��$?�����̅��y��|��y���P	N�U
�J���CӢ���4 �;�c9x M��h��.u*X�����Ԃ�2iP��W�ޫU��|�L���0��昄���l��$�rS��v�B�����#�0���� ��Ҳ �A����-���u�;k�K�1��$tI���!�z)]ʘ�����nyt
�9�L1ދ��ՋWg5�,�œ��)�4�m�&�i���t���������o	��)8Y]�0[�*$o]�����{�ź !!%eb�-}]ʺ@цlD���	���3_�~�$ӏ!<q_�i���U6�@Gd�����
$ˁo�n���<���V�}m�?�oJ��U���䁽itp�
�z��#[e�86D(�ׇ���.g��8���� X:69�����!etNkP�bΰ��E�%���
@�FL��h�S�Q��� (��)+��	��gY���@� ֊���	�~���`.�a�x��t-�eNzl�NԵj���_�X��?�A��g����kg�"l�ư ��F�p��E둕�F�qr�S�\^��xy����:�Ǜ������������z}��ɩ+��4�.Y�@/�����@a�nd�叚͍���b�=u*mJq��c���w��#���{��������;�n(���O<��W��b�����C';�X�X�^�ƭ��nPQ�ОR��5����bi�r���e��t{��(r�+�)m5P��9[M�1��@&��z��!-^�@�i˰ �p��Y�s:.ՙf`��5��w�x/K�;��g��t%�hGw��A�C�R��,J0��z��l3��;\-��_W���.���~���߭��}��w��������+W�SC�oH�N�11H�qc\u?_S(�P	!:�X-9�����ѯ� � �J�d��^ W��e�^98��'�BtU�!�\��ظ������L�;���W%�S �*@�B��M9����@�K����I4����q��i~v�z)@��� ���Rd|�7WР�+ԴSW�M�]�{t��]�>7�l1�tbTsDc֣�u�&�X��\Xн"�G�Y�B�=
��Vaϡ)�ɗ�m��uX-1B0*�T�]ieiũ�| Ƹ��<�P�H�����s�q��=ڠ��F�2G�N�2����;J7F�u��X^ﳸ���H����c3Y�q�@�!Tيg�Ws�pd��fͤ�1�d�i�gf��?l�� ����s�'�rdm�g��ҳq�`��
��0e.x���v]a���J��Ԭ[S���M�c���~Td��̘7Ed�a����kЦR���
k���^�xׅ���Пnh�l��������կ���wv�ٿ�MBؗgW��mnJ<�F��[��Ȁ�[[���fkx���v�|:����8r������|�Y��çV~������K��S����������Y��U �充��_��^}3	��3��עm];�*��~fg�BN�M6�������,���Ԧ�yuo�������a�e���9��ےC��E��\#���+���8��a�[�����Ph(a
�[�.��|�t���t���ZT�;9Mv��zۡ�q�P�$lA�X��H%g�L�$r-�-�{U }E?a,]�>90 �-��:.ߛ	r�O�&��� ��J�._��hٙZ�匨��y��ŕ�:Ir�j�*� Xrw�B:h|�1��:9��uσ�L��{o�����43;�ώ��4oս��3���t�%靖�c�СC�J
�ș^�$�K�s�2�]^Msr�;	-Q���uC�c"����0R��u��J-=�ȣ֌�`�ˈtS[�FM4�!�]��bb�����!����T��.�mb`� պX%��M�T�����S{(�B���u�8ӼsQ ��f0]�z���u�
ѷ@���eؒG�!B�U�	ז�(��G�L�u�G/��@����C,��h�4�7U��9�s���4{��_'9Aǆ��x�N��F��:��C�/����#����t��c,xh\BA�D�i�����8�`#�fԵb�<ﳚ���]�_p��!9���-6O��ļnT,������H��F_X"�%�7`��`S%$��o�N�(h�����ϼtjߛ	�}��M��߰�1t`�>���Ƴ.�*Ҫ�R�gYi�P>�{k��nľf%j������zm�t[k[�\��z��z�:z��ܥ�?�����W_|���/����c/����=�5Ϝ��]�+��.IMH,�ey��A��0�p�+v�!y�n��&�푢�ȱ*��{��5��%@�KA7�;����.��pMN�`Y5 !�
A�5��QU�M1D�[q��) <��������9B\�1q�d�hX�1��O�:)Ჾ?}�Y4���1�(��% ��sx7�Ε,)�'v��!2��˸Z����juP�g?���H��+�p�E!��PKH`gPi��r7$�~��w�xG��G?am����L���A`}��ƦT�&�%9ܤ{��Y���k����>1}n^sO������
48�k�SH�G@qU�G�����2Kb�����ۗ����3��+�=�t�ݪ��e���#��cD�C>8��b'fu{U�0 �yhj�$2�z �-�E�ی <x�kl{)��sN��7���-�m�2�p��b}:� �T	�����vauU�"}��`"�ȨD�>"�&Р� ���+��d��F�a�*��ӛ 0a47�uȁ:�0��6�Tz�/ ǈ  ���Q5���`�(��ЗXBh�� N4i�/�{��y�#,u���͓Mh�gw�و��� U�
GP���:��<+;
�}�a�^�f\[X`�8�`������*$�s:�ԋ�.�����9�������S����m�{��w���/_��n]�ҕ���ͳ��_����^n�ru}���nÊ|m�(���
����\�E���( ��Ya�����`s��ٱ)�ܯm�v����ty���qG{��]_�¥��w^ݜy���w���G�?�y�܅����/�����R���I�������{�7�Kޗ�A��! i�Ԃ(�Eتg�H�4� I~/�6�P���}n��Խ�&�8]vt .^���6��FM٧��V 28#��������3�Q��R��Q0�U�Ē(\��eP�s\�����k!ޯ:;_���Sȭ�Μ9��^�p�@�;W��v�G����c���n�W[���c��iF�߄�6u~��%�!?|?�,5v��ջ�p�k�ȹYD�#T�lU ����4AZ���mͫ�Z� ��_[�2��Z ��x��쓘�k�:0b:>E
�)`�莾����*���9T0׻���m��B���o�٫�g��x�,Հسř�tE 
!�18�3�O�����I�ti �^a���؉q���Z��I}��3�
p
��oِ&��~t��I�L�&���� ���d�l�<=����Q�n��,�� u�4�\t�&�)`��qm6�O�1���4(0D�!�!�nB�͜D<LY�Ua�k���)�Ɵ��^Ը2["�d���˳�>���^��#�/ؾi��\HT���	����*i@S{��ƭfh�C��٭B�yJ�g�}�-/�EU�� |�wb�`�)�1��B?_ ��B�CH-�������[q�g�o���k䦘�Im>�?�*���}� qQ˥3xv	��xΜ�|�	��LP~���H0�`���b
�CO�r�;�xF�p� ����Ͼx��l���t�*KG�i]͎U#hKu�J8���[����i�Z]Z�������DOtO8�٥i튺����~�l�볏�|�q��~�ѳ������_fYZZZuy��ѡօK���]��/<{��^���/��k}w�M��C�.�q}�&C�#9;z9�G综��"�[ٕݫ���� zQe�@���ȠK��H��%���[HѸ��DÄ�/�n�]���^9]8%�';J�"Z�I9:�t�v�rh}��~#��! ��}"�$J���/�O�iT���H�Z��HM����U-�����^�i��q�)�%�)�(����n�����{t��n�)]���0�ːj�cg�V��|I iXί��7Ȁ�C�+#j�H��>�����Ki��ai�4
`Ɏ���}���<k [r��REZ��@sd�Bx.�h1�@Oy2�hbz���� ��YW������[�#%d��Vh��2� Y�
�"<�S���� �`�cj"t@-R��rB�~疛oI/>�\:������ �/;���Y6�FTǘQH��a�%�f,cM�l
1�j,�լh6$���x�)(�j��a���-
X�	�.�C�HE&]�lb�r������ƻ쬪�{�S�R�{����u85^ǣ��xW�I ���B��7tx�kI�^P\���� �M�W}ֆ$PG4Ӧ�C��l��#G��e������GR?�TU�1��EB�+��f���8�D�+�a����P���0�{��E���[@v�,�̋�Cb 8�72��[�!<��<4E����9B�6���nȎc#���S�>�G��~~�G���/�n��Ͻtf�?|�_s���w5}��m���'���P��(��߭�߂�+ ���Rc��T��K쌲�Y��ؐvt�[Z��n�觟�˟�L��mǧ�>�w�5�SF����։ڶ��陹��/^�������zsO�k|O��d���� ��j��UP�r��71��U��k!�p
y��f�m+䑛��Fm/�G�&�jȚ{
qy�J���q�uQ��.b)�ʢ��ށ@uJ hM�A�4���ё|���8~v�%4h��uEQ���Y��an�Vt�9�1�o��Κ�rD�����m��:<!G?R�3꠷������i��&�_�u�`�E8eP4�ژ��E��;8��r> �6a�q��M�kn��F�K�c7�<S;�P�����*��4.���^��ka�t�ԅꧾJ�o	��6:1�9��0�Ì:/����(dCas Nw'�;1!�e�\������c0 [b��*7�`�j��1,ئ܂�Ԑ�9wu�B��������P%����!L �J����K�|"s�7��8�2<O�c�l�y4�7sbì��h�^��,ӳAq�,%�ܚ��{�
����*�H^�bUz�74n��1�j�W��P���~O�<�8�p�N�����s�Ⱥ9�j�*���bߩ�f}U�D�N��c��}�{ҧ��P����κ���[N����t��e�ߓRާ9�����s�L(�[�d��q��% hvthɠrU��}#��w��Uq~}ܫ�C1ǝ$;�ݐV��. ��y�r����[Ͳ���	�[-(F+��C����ە�^���0SS�T�y���g���_���+������B��S_8���#z╙?��8ᢝ�h�	�������S)�Kw���z�X���j��;;]���E��F�9��ӶfqqV@H����������j/��Т��Š)jޑ����-��Ԋ��58���%� �j
���&��P��m��HD&)�A��a��Uy[���k�%��r���&rm���Br���h�A��� �ɉP���n�2T��Q��sreI�Bv�#�ͦBAJ�v�m�1�PMyU}���Qe�W`lP����)M�:��!���p=rN�>�.��e8s	8ӱ"<"����@�uK��#��R�ՄuPE�n�*F�������j�s�V�, �F
��a�
 ���X$ݶa�1���k�JӃ�"����;�Cwݞ�z� �<�=�E�V8X�`n�0;�����#P����f�r�NQ4��!c�0����Q[F�l��d¹Ѯ��R��[�@86:��t�����{��w���S< 7bu�"3��[�ǚ�քlҒ�V�E���b!��B��v0Sݺ~����=W�/���s�p��!�?SefFsJ��� ���M���t��8;K?��ֶ��*L8�1fR�Uf����0�!�ߖ>��f
O�H�����mVl�����
��N����4���.��l��i:ΨB�\�^�fk��!��C��u{�G���{�������<�������r9Z���|�'���`\� �>����P�wܮ�E+��f�B\<����d��b�=�^��YQ���@�l�Z�3N�s��f��0&`��lP�/��4F�W��'^�x�;��~}�G�#��?�'��f���o26�?�4��ǟ8�����詗�}{mp�N�bִP�����G���Z�y6ހw(}�X���)�5��r��[E���%�a��K�,!#i�H	��V=.4yZ���%���$,�&���f!�3�����"�ϩK�{ׄ͟7�;l��D%H�LU��͒��0 �M-��*T�ӭ����N�u��3`$X>��I��#�MιWkLNAj�H�k�f�,�d=ձw���a�v�vؤ6k���ظ���`���B`4 �F�@�M���h���qU��-��5���V5"�W$2ݡB0�b�&��BK�8i���8�
68�jEa4(�=����)��J��nK���+M˖2�`H�����G�gj<�똿��O؉q��xU��;�X�ʳ��a��L�
�-�w�
K�J�C!T��p���7t.����W%�������0g�*���T��R�]�>X��]>sN�D��N�c��)|6�N�>�fp����P7�y����׮^1���1H :a:�������b� �d�g:5?��F�
MY5�PtR$����p��;��M�kM�)�Z��6�j��{*+S�ѷ~٥q#��0#�6��'�ӽ^R��3ʜ���U"aX�V�X>3$ 5,�CB���Çһ��٧n�'MپG�}Rs����<M����o�`���H�H��]ߕ�x���_��N�Ȟ{4������\���10�^/`��/� �� �Z��n�� �C��Ue�e�b]���C'hh�z�^O�iM�D�
�D�z�y(|i�yLs]2�pK]$�<�~q�q��*H �������\���c7]��<���w?����}�C���=~�������Z��v}�5;7ףJ��Y�/mn���|���ϝ���k���&w��u��7��Hg�iS��R��Em^Ƈ`E��z��|���
����I�qy�v�n���3�I��V]��V��P���������ve��q �}����M����dQVl��4����ܪ	!�v{<�tp{R�go���oC]cqvb�@�5�aW�_�>f͌Ő,|�k�R���?�A��{�43��F�ێ�:;��SS|8�G��h;�$T��}����#��	-�	c�1��)��1��BȶbJH;v�\��y]�������_\�ty	R)�뱨[�G��'G�PkR�	��F���!�#骄��W�l�!՟+�r���v����ߚ&GG������@�,�ft\ q�@Ì����u1(4UȆ�
C�B!AtXb>.���Zz�q�'����!������ 4E�CU 0���uT������ �#��"m�����(Ao����F1r+��G��Se����6��/=�������'���~���/������c4�� ���#K0|&e�kT7�J̰_[�W��E9�TB��}6"TC��ǳ��>KU��Й75=#�<0O��L뺄�u�fkn�q�m��<d/ ܟּb<�~ �s
�ql@���SW�?��e���GD�K���ӫ
�1v�.�"S�Mڿ@1��*[����;��/��/x��]<{&=~<�sN��tt�y�7��Ok���ؕP+��
�m�؆ ���d�w�D3Ã5`-yV*@��5<���E?<�4�!�}kg������f��3�C������F=У��Aj]`N��P���t�ۆ6?C�#i�������S_x���/���-�/��412tq��{Y�9����_�z'ֶ���Ӂ���}�jh���z���#�$�k�	mh�ԡ���D�ʁpP���&( �Zi���ROR�OU���kI��שJwۢ|����C8��5i"�{G;"��m����+���C�Bq((*����wMo����r�G2
���
���o��D;��r-��a�X��q��íBYd-���m�[8M�O|��r�E;W��]� ��)8�7��ǽ��̈́$h�J�⊲�S����a@��~-R�?�,�*2']��3�tk��.**6��!W!�>��7xw��w��ܣ�e>|"���:k���+N�)$��g`�X|7$&}��5�4�b!	�j��.!�gD��ij��E�����+ 37�=w:���}����dﺄϑ^/!��:�ώ����ү�c8ɵ�p��38vv�%�Q�6$�: F�R���z\����)a=L#U�	˸E���w�}Pņ ���MM-a�:���/_��&�����ߚV�i��x<}�[ά;�����C�/�ȏ�����#?����F�3?�����E�#G���cH�N�-8�m�7Y�{�x��x���"�QsDv�w���;xPUR��v��_`��KEl�w� @U���_��@}v��"g����qL��[��[�G>��Qi�n��v���<ux[����fc,u�[�X��皀Q��306�Ω8�ɓ'U�aX!�=b�V�z@�$�x�4���j�K�ږt�9����b%���P��N�E]T���$JB,�� ����#�N�R��Q`���j����5�c����F�����
��i-���Xd͹w��+�Ω�Lm%�{t,6	�kZ'���|���0�59�n�=�|�Qe?^M���B����g��B�H `e_X#4}5٤wd�Ca�	i�&^��|�٫˭������JmyeY����>mV$$�JkN$jt�Q�:��^'ew�?��zV�=�hú(OZ^ot#͂е���"ւc$�H�|l��x�q�#W�_�B3�3���C�(Zv����{U�3���K����U-�v��?{{#��k�v�.MO�X	=��}��4,r�Ҥ� �]8Q� �%V�N�]ZP��H�eEK�jA�#�\���fP\0�q��:� �/����pֺ��%���Dz4U������^�h9��JA�-?f���%'ֽ�/�(|�0v@�uZ�F���������4������+�@v���e�N�;�I��.9����O_xQѓ�%���чK�+�k*[`��x��=���`�	�jQ��`�l] �
��(T�ۨ�6�����)���q�Ua��0�d[�Z�7&a��b�L������.�z���~]3�$�x�%���]L5Zq��E�� �%��:9�}�t�=b�v��4�THqD�[N=�E�tB�k���Ŵg`8���黾�}� ��!]�~?�J�����k�腆^��6#�J���6��e�>��O�6�L�qe���Z?�����eS�aCs�2�C�أp4Yd[ꃖ�����:�������O�TZ@޻oOz�;H�z���=\!m>�˦�����Q���i�� �L�Z�RqC2g��Tl�@tՇbp�;�p�E�n[s�3�(���X��e�>U����U��=`ʤ��D��}#iVlO��-�-�_�L�{�i.~���(ݕ~��~>�]��z�[��a�UϘ#�$5T���Yj��㽺�a*u˾+*�@B����J����P@����г��u��1Ӝ��<E碤�;v�q�7�<���s 3��\e7j?����M�r[4����ξ��eK!C4H	81���X��.k��jy��e38D�����w+���
���fCыSr'��@� +��C>G�H�"!��}����^��ya����L���E��>UhF�H� ��P�충�B��.�DMi���E�"�#�^;n QU�gE�2炄�iȜ�E�:�j�ǖ���X������g�B��ٖSǗ�P�`p&�ۡ�{�q�B �b���Ҏ[�ƃ�ɠ01���؀��%�h�9%V�N�^ՠ�Q��bǉ����t;r,��K��{����Mkr@�I��U��Bs�!<�0r4��I��~{�h��-?ܣ�
b�X!&uF֍4m��uL
�c<�w3U���3��y'��svZ7�
 �<R�`���&�T�|���E��c�P� W��a.IɆ��r//9�m�GCW�W��2FT$tb�;]Z��{�x�B�b�ݿ��i�����8�#��7Zp�۟hr�O����������N�jc
�mi<z�:�g�L���!�	l��k,��@8�K�<�P*Y}.PIͪN�	1v8{ݛ��%�:>�%��M y�,p<59��7�g>���#{'�J�2�X�M�f�3�M��9��@V U��}�7ڒݩ15,�熼0pKR�́/Bl��X�O�n��MR��w]����V��l�;�i��P�ĸ�i��yN/��y~/S� �K���w��xK��ŕF����*}�S�R�	���)h�A��c]``�& Ê�:F�\x]@�j
�\��i��g_Nt�Kk�N�"��=�&[�����7?���g�b�ٺ�P����s9��W26v��
c���ye�:�#z��n�_�k��$����d��i�ƌ���
�Q�b�����釼	����|��b��nl�x��2����??���y�����o�V�����{/ �;_-��Z��+����E�aBX�nm�`�i)��8�/g��"�$c��=j!�p���.�n�m�(bs�WHyMC8?t1>����]�'��ӭ�#������I��c����Uw�!jȁEJ>�M����)�]� �4�u}�
S���܄ T���rP��#
mP�fa���Y38�#���gt@0`��I�p:q�z5���w��G����\Y��i1�7���P��>ir�q�r�b�?�}������,ׄ�c  ����\ǖ��9u�:��}�^��Ħ]�9��Y�#��#�˂e��|~Ga&*�l�س3-\&4�ݵƆ������bm����;Q&d�x�b���>�������7�QZYh.�Kߠ��(g�/�G7�����t*�l2j!Q`@� Ӳ�#��S��^B[:6��v���(j���&�F�} f4w�/%��w�l:]���ۤ� R�歃�w���0c��������A�Ic@}*� �0�#mK�#ѿ ���u�z���N�G����QL���^�/��M�$<�-����Fu\���U���316,����;��)����lBD�����tTz��Ӣ����?�>�ɏ��S	
6�\�L��B�� �QK	^�ƽM�'�L ��Xy�����+:<�]
�څo��*9����VʆjfQ���t�ٞ�^?�̎����Y��τ�d�pi^*ɀ���b����#�5Bˇ�lS5t���P8���Z��	������[��`��nly�ՒC�a�[���A���f���倝׻��R<�;Y�p�|�ز[N�L"hkJ��f��7��� S��K���X�U�5�q��r�0Idn�c�y{���GU�%~X���-��8�馐��:ęjERA_ b��� d����s��zA>x���Y̨��ҏ�M��z;UdN�	���X����A��eǣ��K���R}���p�8�9���hx\���k�I�%ݚݤ[�Ȧ��I��9��֨�ZOVZ��Bf�<�v�q?ts�4��l�����y���i��ElN���zE�����ލ��Y�T���@`ѕ�->W�E4%�#(<�����;��u����l���q����9�9����	4�]��;��[bs@eS
����%6^iu��#!��N��^�@�}[ N)����]I��@ˉ	[��iga�,���$���c�-��"��P�pC�7�
0�!�o����fz�;ߙ^y�e^��, Y�g��S8x~i͟!�kR�9��4f�}��J�M'z&X3�l�
�~�7ؕ��W�Ƚ����k%T��.y��h��j������[k�n�1D�E���*�`K �B���*�wHn�>{D���[
�1v��`t�[b~�._��a�nI`�{c�cG��(��x��q;�*����|�Nic0�q �![�HO�K	�I�@�'p��Jr����*�S�T��:6��C]A�Va�j��F�.�X6a~����:���g�}�h[!8��"zD@�((�c�JB���ࣜ>�ETscΡ|��a��n`�x�[��(	-tR��H��ubb�U&^���o��Ui�o�_����@�Y9Z�W� ��	ƁE}YRT��U�R]�(�n#O��$h.efh׫�&�+2��1�|�j����S�0 IH���/�,�\C�
�[ab�u#J��AP��Y_	�H\�
��n \�cO�p_C�+�{�= �Hq�����PX�;�M*���ZG�Цt���Bg~��qũ��Td��g����0 �r�M5�DD�����Q�ٴ*��C�K�(Ш
F��@�)�+�}c]�D�;�ޏ`�����j��F��p�a��ơ.P�!;8=Z�min5��� ݒ��k��Xֽ����n�д���f���}�I��ݷBH�
ڮ/�����~^�O>��3lV6�R��tVs�c�=�
��J˲��y	ʛ��(F��9���ngGV�;�H�B����s-Oy�7rO��+��ԔTP�¬�����9�9�p!��t�^��9��QAS��W��{������v��X-TY\ ���KU�E���k4��(��(H�z�'m��XƁ}ҙgt-l(�R�#��F��~�S�%����Q��4x��y���[o�5�^�v�i�y}?41(���A�*�y�D�$-�E��F4�������WU-}%�}�-�c?�yN "|�%@��z�E�hj�Q������2u�^(e����j[�c��L�U�9��u��Ɲf����Dk8�B5�X'�>�M���r]2�����~2�i�b�Cm)�3F�\N�Gn��9����,�fэ��.��_��\����r( ��L���'�;';0����:���[9735~h_���9u4�Ĺ�|8��_�f�����I�����d1h�;|X��g��q	)������i����y2�^:yF�W#�w��2rX(�q�,��	���>-p�C� U@����&V$�)�J"v߱������\�h$�T]9���hT4Qѝ���v�P�M�����ٻ���	fڥK�)�,5sQ�O��qF̎mRlqbXH��C�0�ZC�~i4?��f�uV�BϙE�	��}JQ�`��� �����hPz�����%F!��=F�B;���Z+-�{!��G��HN���f)�,�j�G�Ύ�GST��T��˺:g������p��h{!' {��ձF^�C�3}e:X���zo�[Il.��P���+�J_C�x]�Ϩ�)#����}>��گ{XT��`o�B��:.���zY���E�D�X��QhJ�X~��b����'�dv�veM��h�� ��=-�\ �����:����Ջ��2тD��>�o�8�,V�l��V �[���X"|ZS�.	{Ra ���b��w̯FK����E�(����^fP!�G>�Y�T�)���c��^kҢ��_(��P����,ρF� ��B���/C
ա�!4��� m\a��jt[�q����׻G�	�5��f�N�p�rR=��P�˧^I�/��>���N�������a*�ܰ��Bx$i�%Hff�M"�Z@lN%!K���yC�َR���^��"A���z6�W�n6ȜU!O���zl&X�Fp$�nj�p0m��l${t�x +���C�\iz�����6�Uڿ�6���%]���X,cc`Pz'/�:.���jَd��z�X���i=\�8(:-z�`�����Qv���ľ�K_�3?�b��8��x��xe ���gr�_��o��~�NO�oC��[S���b�~��φ*�6�ׄ�dKd<�
�\X�0r�����#ZMW�5��F�E��3�`bKء�|��6;�j�=j���ʙ�RR;�4��������t��iD�r��I�J횮Y�4 eX�7��H�s-9�%u�v%[3�g�~���\������F9$�ա,�.e��G�P`�N��G��um����vP�4�������P	Z�B�F7�D���!���"0��Cg2+��sl�tc]�C�
֜V�v����BX{@��
���K0U�:~}C-h��r;��t��R���řn�@_-�X 4@�Js�{�17P=th_ԩ�(��}�۰�]-N_L���)>��;ӿ�W?����ȭ7��'�����g���c����n�Mb���W����~�sk���H�0�Jc�!��/�x�޷���.�)�R��^ENjQN|D�έ֪�?����	9������/�ZtK�Ʊ�nN�}�{�3�>#��B|�=��r	f]��Wl^=�x.��.��S���j0"�`�X��å�CU�yA�ې0VB��ѯ�ބ�O� ���8b<�oT�R�w��DH���5�,��Y!קIbM�dW~�:|D=�&�?�ph�����ds�p��t{b�t�>��e�����C�.��N���-1���ZP�[���ҽ�1@��3��W�L�%��q{���z�"�I�ް��E-"���6I��\e��	�	���K�>ܣ���wަ>{W�yղSA��=jƫg��6/��0I'��
6�)u>K�}��ҹ��������^���4�T�u�g6�޺Fo3��Z�!�\E���6( ��:�ڠN]i�".���F����x�}�� h��(�ֻw����Ϙ�@���(�3(����;1eCF@�d�@�*��ЎJ(4s��������:�g�P���pگ]�ჇҔ� ��A|K3O0#Y����kYRk*a�tb���*�J(��E��ǟ4a�FH]F�����RD�4��n��M]�95����S��L�K)�aѯJ4���]�6x����Wt�,J�k_���}��Tm*%�n�t)�4 �=	u�I��룏�P�8� |��\����B� x�~&pJr��V��ϝ9�{YO���S�6i�;륅(r������΁�\���=�r�83eI�αp�##��������P!�5e��f��8T��fB�a�=.� {l��:sE�PHK�������O�
ǜ>uQz��t)��Z�VbU��ȳg��s��O�����l��?���;�Eao��&eK�N�
=-̥�g.lq�Wԏ�:�11M�.N��Z]S8S��Bt��9b��q��iR��Qm?4�hR�o��؈�P��9��4�=�"�S����H0��i�M
\�m(��*��²6�Y!�%$yYU�����^	ꕄ �2/'���z/}9ds�շ��	9�t�U�L9���m��/�=Q�0V�b=[ڌ�h�VUoHa�>��}�d��ҸB�=�I��C#b�$���;���	ٗ.MO�g$=���\�/ϧ�E �4z�>����~���vl�\b ���1�e�:֣^�l��kda기pu�n-�8�<��A������!{Ϩ��d:02�f4ޫ�
e�l°��t�Z(�Zm"/`��N�l�;����E��d���� g 5�z�a���5��[E��6/�z�>?�\D��[��� ���7,��Ǘ���r���bވP:���p���rwx��h��Q��#.�0b�F-vBQz��lsUU�U_�S���u"��-�K_u�A/�dU�_�@C�gT���B�w�P��޻����f�M���-�d']�4m�r��-�v
΍�+�t����2��I�:��`2x��㢯SM;�&Y`�nX���K�d^�t���wɡ8Ӱ��nBB���{C�u��]w�)0�ߡ��.�/�2�A�Q:�~L�k����8 ���[^ZM���:m�nxV����r��K��F�J'r�a"�����	�
�d��3ϼ�z�Ś��MKk3>��@�m�S�e���h����h$�}�b����h��:�S���M_��Uꢎ��f9�G%Խ��;��
ƅs� =v,-�Yx�;НJ?�o~A�ߢA]��]~ŀuB�=��p����ӓ�=i������L���#�>m}՘��q�(�p�4#����cj9|p��Ƣp�2�>��OHܮ�Ld+"���#5{fTaN��������/��
s�.�|��~0���gĨ��kr9]�f�P�=#�R>e��!E��;Op� �7h�ک{�O]]ivA���ae]Q��܅�tN)���Ǐ
�H#4��ZLoem1oǾ��t��^����(=����E9�p�knf���H����`��O��X@� �p�0k�#*k1��Ź�E�a�-��+��vҾã
U��[WAL�^"ʔ,����cK�c���H�g��/h�#�G�<7��Ph�������@��A��OD�K������0��D�^ �na��:���֠��1�5r�*���ޢ���&�6���������#�{%tJC�H�<�Z	������D�ȶ�r�4C�E�#�lT�Hk���=K�k�ֹh�����r��p壿�,P@�F<@�gAU�d��Bp_Ʊ_��ˡ��;�, �d]�f��Iņ�q�j�FqCv�0A�/H�7
�,k�S��_�?�wT���	C*����D�������Ϲ�z���W���Tz�v�6~`���4�����3j��k��t�X��'o9�:6{���%-����s�������EU�~��e1H7Yw�͏�8�p�L��{:�"�,�02�����4���~����s���R�ȣ��tn�ً>�1tQ@��^vcО��t,]����M���߸�w�r�O<��Ğ#i�7|cz��g�g?�i�3�^y�q�#��t��K�������5��ܼx�T�]ɬ0�=#\��yF�����B@�鲪2�t�tD�L�������ω�9cVbJ�Y��G��/�w:�!�c��^��s/������t��=�2�����f���y��xN��}D��ų���}Ea�i�/�A����R�d��������О��r�Mi����w�!1�z���B�U�>���d�x洳�p����E��MX\�C=؃�n�%�& H��9�6����^v��;n�-=��/:����':�%�)���L�n���˳��|N��a�����/�1O�
����3k����f�&^��"�C�����l$H�Ǟ�<��Э�{�=i���mب�)wl�pZ�|:���K��t%M(kk|r��g�{�!��=궮�K�#���i�BGp����_5�Tn`c����^���A=?bFHP���͇��ҵ��ɢ.fߖ�[1/��"/�~A��A�N�鬧[�H�|����
��.�
�c_���
dV!@�"���PԪ� yV��1�.����iI�NՉ�;��Wl��7����~��P���0�a_O���^��o~2���s*Cp ��_��tEl�O��_�5ϊ�����5�E�{�	��b��l�h� �p]n�C=0�I#���%� ��>;�^1�N���3��V���md��n`���S�Tw�U;34���5/��
��G��i���5?�o��'S�|u= b��b�9K�
�� !�"���ҀH,�t
$�@���-���E��&h$�j
�I��"6��wh��u(Ty^��KD[v���oI�	� ��$<ݯŐ��+�O�a��{q^�刾�;����R<N��u�����=��x�&�b�Ω�����E�>,�1�rp���M��=�,��
q�X�3�+xS���<:��?�ԓi��@���ǟ��q�^ph뀴)�NZru1$'t��% a�}��z<--	<������$��F���*�'i��Y�.�M�4&�O�u�E"�[��_T��lE��K�EM��7J_��w� J}^���M��)ܢ�0N	��ē\�	� M��(d��4�N9��Ys������{���B}���뜯�������ޔ���ߓ����#E/=�����KgӃ�zH�t:=��z�	��,���|L�����Oֶh���?>6��҂f��#��^z�Lz�����{�I�&) Im@L�зʾ�� w]�gK"�=���8}����:A\oKs��ԁ�'����Fk���M�y�"�*6���oV�W�ןx�	����u�l��E���z�g��5V��ٯy�{ҷ��o���!fQ��=w�cG�X�{I`��[�������Yb��@�P�r�T�Am�W�bH�H�t��+�/
|_����y��&ѵ X������{U�u��%e�Ix|e;�����ྃ���~�����z Ι�jl+P��x(�T�|QdZ����X� 6(�9��Ԁ6{Լ������d�� ��l)L!�:J�k�k��Z�s+�,V@cq]�IkG��{S���7L�����A��][���7���tif%�z�X��_������MiN�8�7���̃>�G.'K���zk")��^]fCKZw����%�ޛ�'�笣s�X���G�/g�z�|����x��@���<����?sq���к}N��0�X� ��`gۭ�����X���k����
Դ��J���u��3 +�[2,���X,*� {)6C �-X �C�'�'W��J��)����	�
�����f�mA(uSD�;kI��H�GT�b� �!`�*�Ǌ�-�0 X��[p�O�$�J��q�|�^�/��iPo���d����Pz3�\!��܀վJs����B#B��S�-�T�L97�|��
���Թ��[n5�N�����51���̬��ȴ�q�Ȱ8�U7s�"�%SL��$ȥ��Rck�g [��sCL�\^Ĥ5�	i��&��p:�>��1�'�h���U��qF�����N�O��.�� RJ@��t~�{�������(���'u]׃͇�A���$1�£�O�M8�= M�!l
�a@
��pP��4X�;�R E�h��~��#bY:�A&G��hs��ü��d	*�$�̈́X,� ���y[TH���Ɗs2g��% 
�}2oI�� ��ӽ�48�h&.!3�}L�1�E���Ze6�c�Ӣ������ �5 ]ծ�ܫY(��W���*��XX�1'��r����W0S
�!���(�,�h�0����#-�΂ަ�cQO�63���h�*։g�J�$,�=��Ç�:;�)�Af�������~�5)��6�������F��-x.�A���(�U��֔	�-��.��>e�W=�K
�]R�փ�'�50�����pz��l;v{ZQ�vM=�ԯ�W �=�JenlS�T�K�7n	�4:��LN��|HSE&b��6S��T�-(�"B�h�A�.�G�\��l���~����w��W߼��/Y`�/�"-P��V=JJ��nzU
�I������5�X$���N�H�]'���!� j���G��q��Wquj��?ґ������ήyJU{7��j(KpP�Z8K�}�C�IB��]�WBM�	@�{Se��:r�z��'c����h9�ye��j�cG:�P���j�Cs���E�Ľ��㡗�8�4m�USC����*�=t=� 5 (�;]�G��ͅs��TwF �].Α1bf��d��%��>�R9$����*��3���X-�
sىj���^`by�,����.07����G�u]8+z]�k��߇4M����5��P�5��@���&��Vz2�g����d���q)�&mz @aCYt��~9:@��3���2���bAp|� hB�3/�
��>����Y�V4�Ԉ!(D�B�W4PfJ䬸���H�<*�ɹ&'��"��ӂ�H��r����x�{���\fI���!���U/�<'�,'�y��]��͙�*HO��
�ҏJ8Y�9�{�-�<[��.Q6s����+�1"��Rr�l�"��%���w!�F #6K�_�a5�j��u�;����=D]�R󆐧�kc�,�HB��ss邴L�c��X
⹠�<E�E�Q�s\�)�rN���Đr�%�N@+E4؉��g�j�T�����E��zT!_����/���3x�-7y�_��r2bn/=ۢ�a3�ߜH�x�8���$s�RS�uv��w�s�ΦǵY |`J"k={�A1����0X=�=H��"�Z��� 5�Q�Blܧ~i�-������³���uI��ģt��d36'nz���d�u�=��(�s"�$E��u��%���o��nh����5�Ru=��SHVC�u�q�Y��P;�b�z���\�z=��n����k��:vCi0G�u�U,��s5�pL,Ξ�b<7;�n��f�E��iр��'�o��(��B[
���84�����/j� ���^br"B#cM	;�U�[b �  3N[6�D������j���M�N��jĹ&N������u�5 �Zd��ڽnlj��v�8V���b���%�?(x�Seg�u�z<UW�~��j�p~*2�^����k��rVїL�t��`g��Dqj�Ú����s��C������%q��(x^�*o*M��
�/ؤ7��)�77��@�_!A��4d�K�ӗ�h2���;�
z��jΰ.�۬a��6�+T6n�gB>���:2�)2�65\��N�*I/8.��QR!�|d��~p�0^+�WUÈZ38������cӓO|1���,�	]�4�#zb�Rd�E��q8kw���n@�ٶ��r��|�A��amqO���唙� B 5�{�5�b��I@��۹��k��3�g������و\��nXlд�ܑ5$[�9�֘qm�AF&�}U�Y�ߙ0Y'�k��V���3�ƥ�5��c���y���^_08�����F�>��%���c� �\7��;��.�#��( )J7Q��f�.������H���<?��ۯЩ2��i�;�7휺���J������Q��6�k�Ц������w?���z�K�2�6kß�=H�H�Ɩ�	�S8K6��P+�_iB8�En��Nھ�>�mK��7�I�!�Q>����#�]�@(@��=HdAٵ���J
;���/����z- ��D�e͐�	�U'Q��SL��ڑi7��L2���[>$'ؗ�y�Q��A��X�q �ä́�`Q\��d���珤WG5ޖ�a���������$`ҙZ��DNH[�B��V�Q̉B���a^�Z2cƂ���s����%�:}�;yt( *v�,�d��&{x���C	9B(-�2�U�F��>id�h��u�}��1' �� �Ь*d�]1eq�>�#��ġ�f�a�wT���'�	$��qЄW`��,���Z�G���7���ȱ	�^��ΰ5��`\�b��Þ,�A c��sƑ!� B�(s������CA�fg� �)I�
�ܙBUצ��D��=��l�������� e|希@����A��6�bh�{EY�̗��G�&�K�R�>v�(2n�έc �"+}Γ0�YR���ӿC��z:�(vP���ؒl  S����y`��f`Ђ�3;S=�9k���w�A0��ha�x~�!<�k�S�٦�X��J��mA�����u�6��L4 �eF�7���y݇�m
T���f�yX!69�dZ�w����?�ĵҎ�1䙀�@�M������6�>��������#?��Nec>��S����騴Y���`�$��iG$`��y��jp��Vm���WS=��{%�oJ�7�.�xg׺Z�4������1؀RQ������d�$����҉ae�a���7H���x���?tCc���ʊic磇hQ'�r(��H�%&O��x�Bȷ#�u�+3>�l^\�7�&s�����7��W�>9���w3ͯ��X�̈́��[�ܜ�������`Q� -���E��y3+��,�T��  p�cڱ���n�q���08ZO.�c�G,vktt�U�-��s�\�8ֲ�3�np����b�~��m�3�d{];� c��"���'c
_紨�j�A�;X�i�1qr:|o�O_�<�n�N���	sPtܫ[R躩��#ॶ��q�f� v�d�P�'�;y*�g
j Y��a�4+�Ыv�W�/�X �F��?)��+*�R���+'��������x�2�F�궉5g0R�S�0���/�̎R�N�ת�UP}0y����̬����U�!��9�j �K	[��+V�-j4�C��9���#����w '�^�!�M��q�{�h�mL���"�\���bg~�+�]tXp߯q> �μ��y��īR}��a��* �"�����5�r|7�����j	�2 �*�� d�L]*2�(�9�{��WWdI-W�{L�o�0�:6v�=���]��N��p2��Q����n�c@u9���]~�=�=�닁�d�	�ӭ�R�{.3/XS��X�U�h�O�&N�?��:#P��c�Z#�*��ܓ���V��ꏤ�nR�Z�^����������ߦ����tǝ7�����?}����G?�x���KE8�K7�h"�������9�Q��VsK�dӅ	�!��V�pA76b
�G����	$@��+�iS�±cǵ��*��x��M����3�^㕙�b^/t�+�8�6V�4p�m ���jw^���+��c�#vY=���P��agG؁c�T>Ο1+�F�솾_�BgQ"�%��?��MJ8�4#*��3���tt�'�=l�Q7��iA�,B�葚�G�Z�?����Q�/�!���\�J\K]L��������/�+Ph�B�	¢>! ��o��@��GE��ﷃ4��=�^P�'H���6��K�$v�f��w�jnݑ��� �S��\4��e�_,0�}#�� T?!0$��rxF��,�N�x�8Yvv�hR(9 ͔� ���$���,�Q\]�;h�0!(������"�=�e��0ЉƵnJ* [��D��J��s�� Pv��JC���*�n�j{Q9F(jOMN��q��z�|�"d@+�\\�6���95{W]3����A �h�g#�	q�Ց-�h��]�K`�hx*�K���ߖ�Դ~�V*� ��|g��+��QX��#�+𰪐@��I���_�5,篪�E��xƢ��������S��%�ı���9L]��-�mk^Q7,6��B(���(�#(��ϛ�̦�d� ��,n��4�k�1��CL}�=w�.�*z���1Ӝ��ZWVY?���--�)�S5��Lz�R�隵�.�|6�\:�nW�����?��u�Bjz��~,uJ5e�R��Ǜ�6��P�V��c���ּ����zMO�����n`l���ŮhH���[S[�!	�P�����E���z��k]J���g���Z�͋�w�U/���$�Ź��+��� ��+fح�||��F��g?����A��x�t�
H�����������u���ɱ�@�� 
���P�&��#�w�-��:���v�,�#����ET�p0-���x���]��+��A���z�+'S�;N��@�G��7������ٹh�\u;u��@}��)�������8 �1˃�z��~�M��N��2��Զ3mZ�XlQ�~�����A�
Y�*V��XTڥҰ�V�ɚA�c��]�X� Ж�{t3V�	���o�Oq /�J4��热a�Xo�{��Cv��¯u(g����fe;��`Ć��p��ꡕ�>�$����ju��^ )Y[��ҍ��U�ul;4H+4Q���|�!�Lc��ap͜ �	���������!?�=�3b��J� ��Y�=, ҂�zc�D-��
���Ǣ7�5��f"օ`� ��(�K�M7f��q�~���C����Y��<0��c"��7@�P�x1�
�m�S����W��k��䚂��S�j�bv5� �lx�n�!|�W���	T�q�/M����Z����	������2��z-�l�����c�k����CN���������/�L��o�]��u	��u�G=(h�K���"@�7�?�&]����<�dW�9�~ۊY��J�@A78�0�0r�������i���.,X,t���Z�a�|���ko�៵H�]�N0Cw`�������^	v��r�,�>�#�G�
����y�s*�����*�\M�k�A�׊���y���-�=/�i���H��=! I]Ǧx\�?��ԎI�w�R}�H�IKa40�:��]@�ԘZH��n>3`>2�B 	c;B�#Q��O�\*�G �:Cs'kl������gsp�B �
�Q��{�SޡFgm�h�ն�v�| '����3���}�Ҷّ�N��q���A9<Q1����_.�� ��k����>��b�pr�8i�� ��{:��񘹪X9dj� b�]dvˬA ��u-���GpK�,�������� %w��V�����ED�ss������O����~��p�\E��z��� ���sP1u�^��E�Г��A��9��\Va�G��?[��쮬!�Uq(v�z$2�"�	&�KZ�(y�&�Nr+v�Z�R:�8��(�����T]�5���h�|�+���y��_0D=fNSd{�06}�{%2�h��<>K���U�L��<����>���я}ʡ?qQb�g��魴Gw�T������ J��-F�v�*!�������O�gU��&���M��GT?죿�;��q���߭�PF�J�+s1�ɘ �h�<|M������x���me��nd���(4���ŋ�2�!�ƙ~ܴ8�v��A�������노�P�{ ��ڭ�Ʊ����N>����Ԏ�ÅAT������@����A(���S�����<D<�f��Wny7�Y��%�G��G���S���ZVZaG�%�oD���6X�lĪ���R��cf�q�;p�P��� ��[��"؃{qxR��wQ���M��C��w7�Y�>e�Iu��"�ܣ���Z�T�!�?����^�Vs֢�Nٙ16��|���<&U���T̀5` ��sTg'����a��Y�| 33 X�n���  ��z�TL�� ������!�Xv��(^HM_�O�
���J�gF�V�Tw�ze��	��� i�zs�߮��_�q�X<��N��
'�ōT��ܩ<O�;��d��
�
�G�*�/�\��/!t�W�' ��F!�T�*_`{��{蘢�+�J�(��1~�z��y>�t�O�; +%�9u��J�3Ĝ @Y=��-���~4h����۠���J�8�z@/�&��z�G��WNk�@�OT�����+�!�z�;�zS��U�?�$��
MN�ێ�ǀj)��gYa�Q��P������>����[|�*M�j�0�ޠ��[���0k�ϸW����6�Z@��]�<R'�X$a%H&D�߰��@8���ӗ��uA�70�ޟuA�y�^0���9B]��Z�w8����_��_C�gRi�CC���=�]��� �%�Cw�����iŅ�$�`�Wy�_�8�� ��.����E2ĴСu��:�ߡ�!�-����L��n!D���J����Z��S�A�����Y��G�T��E�AF 	E�2�tH
A0�S�T�=^L+����b ��lv�E��札�?��Q�$�+�fj��)�r:_ճnU>�!�D80�f�{��v��X��g��X� �h;�*܆�B� �@��b��k-�BQ�i�b��D����C�D��vE�b��e�+0��ư 3%iM������"C��P�u`� ���eJ4�\�.T04�˜EU���r��.���2���s�9�s��=8�����B۳��V�b=e{�tm%��m��.��Z�e`�Ƈ����&�/�b{i��Fu�j�dMZ:zg��s���1�L ���5ޤnU�N��<�z0 k��;����NY];��@g�l�P�]���$�� ���Kz��Ҡ �Z�l	,�m8:qo��{D�ɶ��k����B�ϧ�S5x���ծi����U�W;�餸·����Q�����̛�py^�y��o��/]���/_�( �؋�!2���B�]$R42��EeYB��y�*������^��}���b$�~��, }���xy� �+����G�%a"�s�^�ݳ�=�N�<�+�ʎ�k�I�C`_�E�(.����G�+R��y�v��u��B֖�MD��OX�z��5g��������&v���8\�0C*��r/5] �!���6-�Գa�cLO,Bh�q���w�Z����=��� �/�Ѱ?/��_ΒB��3����1��rbLpN�3��	ge���˘`[�2��?-��d���F��x�tXW�<�Z)������� ���p�<
��$������b���b-64Nd�p��A8ƃu3kU7�Jg�)L�k���N�ah�jNȆ��\ȦZ�c����+c�0��	�� �^�����<���_Fx2XK^����'ol�� ���*8����d�t)Y�_� һ�`P=���`�u���pb��K<`���W��+�Ɵ뭴B�����D8�Ў�an� }M���e<�ޔ��1Q��W��-��ੲ��"��V�2
*R� �=��	���8���e�9w�!�qe��U���ǞH��P�cbxb|(��-����H/����S���S/��o>���C_������>�ZHL��6�VT�r�[����~G��U6!Ɨ�[��D��jm�`�aH��Q�!�X�</�_�m[��[����i�� VO��m�, �Sv���wd����j��m8vw���/;�|��s��p���X���Ñc�X��ي)�n�b�u�e�}^8��[c�(!���R�O���ϸ�Zv�A���Rz,��w��L�7��y�ov"�ʐ5�� �0�=@���~pB��PΪWY0�I���3�Y0�/�uX�96�C��q�슲m��W��h�����0��E��"/��ٮ��������[#�6��m��Y
E�"�j�E8�T�(�3�xy̮MR'���}.��Dx�q1;���yFc[�	Pv�!���c l�K�ܰ��b�]���w������}��	��}f����a/��P�X�����7�RM-;6�X8)D�����z��쒾���ܬj1e�n�f8�e������+>����󳗻��>��: �V�h�0�+Д7j�� &���&Ѻ�HK��?�"�0����{� ��� ,��9�ˡ�T֨ut*���me�u�!�ҭ���[���M �b۹:{<[�R���������Y�Ϛ��;�����U*����~�JSx�Jh�=c%��ܯ�aSz^�g{�e�5������Hz��ϥ�O~:}�7|M�����a���H{հ��3�%��]�.��R!͖�9,&p}��:��fgws"�Ҟ�Ǒ��H�`m8J޾�B��sX��ʱ@A70�b����Dvj�Z����a�-��wC$��\�rm����1�	�8FZq ��^t	����T?
����?���~B�wv�~���8ip�[�H���8q(htU$�2��}�Z�n��v#(��"Ev��v��P����C ��DQ�������0A�; �$=s��$�uW @�6,�؂�3EϢ��rc����^��1��L��rj�r/&>��w��ϬL���AH����$C�0����c�do� ��Z5Մ��Ɍ
JUx�c�6�� ���@P��F�}��0�ò�uS���!b  DYU�dν���`#B�l�g� %g��T��|UP�خWc�]hQ���d���ۊX�E�b�6���w8Xq��ae���E,����2��L!Ć�'Bd�x�0hy���Q<S{fs�У��`�w 
~2�J�Y`@ ��I�7X&lN8��"��r�ޡ8��f��ɫ����3�A�k2Us�S�����}���� ]�@��F���흡��`5�2��a���\���w9����L����o���BXqe���>�5+�k�I816����>�9��:Y{�y�"���|.�-�N�S�ĥt����g��;�D�f��?���o������f␒��*G/ϜK��b���F�[�'�֮\H�c{t�z��.�a��"k��(�bW���W%z�yh�vTF*_�b-P@��ŏ<�dh J�	*'��v�*Ȉ����ݰ׫v����Z Y8��)_c	�q\,v��+����q|���� T��w�����[hГi3(oiX�F�����p}�(�F�`��:)8�\Z�EH�+�O�Km�N�#3X(�ƚ[.�7�X2L �K�$9/@����r�1�i���p9��a�pX��ݱh�� ��w���"��n ���g���}1_BZ%
*������b_Z�-��:��C�N���T@�V�?�F�v6�Af��5�}p�v�w9ę���T�-�����z����P������s��c��k�=�dܶ�4���O�;�!y��kO�ϟ�kf^��:6a�<g�O֥�����G����,����JDϥ~O�c���}سhIr���PT1�c]��d���|��+��L���W���b�}����^��m���@�ȿ�� �s�H" D��</�^�r9P��cG��)�R�'��&�k�Јjw��r����<���ȁ��?�G�?���N3ϥ��qO�'�׿M�<���J��a��?�W�w}�itl ��?�'����ӿ��O�ob'�y�0 쫠S���bp�h	�fr�Z#:{<vz��T������`{�(�D�t�~��ơ琉����k��ݹ�ﳳΟ�#m[���*��j��gX��
��� ��r�.�c�]���w����e;ӌt�l�VxD����P�:BN���v3�!>^��d���Ǜ�V�� �;��8qt2���؟�+ʎfTUfI��E����p�.������l����B}|6���x;�g&%t!�_ΔȎ#�K�4ؖ\K��f%8��#��]����jg�vME��]xv��:wY�G��+g���h�dp��(�;��2 �Ƥ�g�\�C���w��/�J�l�>��=gJ�����אs{j?���y��8��j��5@�F���z�����"���=,WU@�kʡ8�*Ӕ���ڀT�������̸0N��lg��}�5__�e{g`���������E;j�����Ξ�s��l���pc�?2��!�&������_�m|:�o��� e@���N
$I�S�V&m� g�ZS�U�`e�R���iY�g�sګ�?��%�ӟ�����1Z�<t�	�W�Fu�T���w�'��o<�Z�
wB�-��-��Ԑ�󘯊�Lj7�v��IL`�T^o't��J{vA<M�2��Ȉ��o2{�z:���Ũ}Qs���][��]�S9*��8F6���'��Ŕ��"w�vh!X��c�A�+07$�Uj{%.�h������o��̠�㤚v���q,.��G����ݮ#*\��z���i!��P��δ�W�q�bprd��{r�C���uBUZyδ���`�||��Z�ɋ5�t��l�v��N���%������w����PSe;Gb��[W����k	&��fdG�=��U�ZT�_;��E,�|F0*`G�q�]�3���<U�I�f���������Y>O�_��8�R�#! DnF�_�u4g28�X�@(_K���}�2@����S��X��A���b�2C����Ӟ�9ڵ�ϣ��lH-^yN_Ϩ������Ή9a�G���r+�/�|�0��$V���σY����v��k�6kg��!���:!d�M%.P��[k˅��s�=�z�^_�������g{C�������:�����ӿ�qi���&������'T}],r�v������Ks��JX=�������C��2�$��5����C5h�:)��Z�X*��<n�ύ俜�\��ֶ@A72~A�����9[&��*QB8a��^h�䅟�U%��`�'c&S�m`(�C;�l�Cw�M��~[do4�k�9��z��%RdQ��d&�_�bݍ�F��c#lT�Z10?�?�^~���o��2�,/n�}�rF�C3�"���]�v�R9;Z�M�?���I�Z��G�\��3���(h1(B٠��vod�j�Ɓ���z�B�%��0L�E��#L��:��x��y��k9~�w�\��Z&���Aq���ö{p�w2kD�̙j�Ai�σо=\z�p��<�# �����^�Η�v������D/�-�>\{�厪0bv��[(_��<��9���<��͈9H��k)��X��t���ܱ����g(�_���/^��l��L�#D������u�^ZZh.�Bׄ��Y�L?>ü�=��B�و��q���<����t2E����'5����T���ֈ��u\}����\��x3��{��
���q��3�m ���y��I�;����F6�j�#Y�Z�\1Zz.jt����>Uվ�������m��Tk�.��첢=-%V4	�S�[H������2�������FLY�U�jC6��Bz�����+�o@��c��m5\��I|�u�[��~t��ŤK����k�p��GJB� (ov���W�
����Â
�o�U�Z�^��B�Pe�x�Ks���f��n*�S�+;$��m�bU$�XY�I�]�r��S�ISo�MB	I�0� �Z J�8e�ә��
0�:��}����N�N�v�`n�L-�Ut<"�q= �@tnc�����Z�Wɤ�D��T �k�K�CF|Ζ>5ObQgA��C�s0]�fL��*������<q�0-v8h��69��w���|�<��� ��?�Ϻ��w�9�9W��1��2���l��=J�'�M��EA� f�c�(�r�^�P�'Ӎ+�˅�48���C��*�s�,�\1��%���Y���=�Q���{?�a��!� �U�r����~�#��Ρ�0�ưC��{f&�~)��s�a����i��$����ɽ����0!p^��z��g���x��hZT�΃�79y��ƢP�։f�yn���������-gp�pf�8e�9�Ky����P�'�J,\o7�ٶ�p��z6���*�]�-7I�Xi)�>��j��GL<���QC\���^HT8q�ѩ�óʜ��3�uakD�qT}�Ⱥ՚5��GBt�Ue�=�S�(����t�5�e뮫���O��ށ�jk���w8�O�(=���ɖS�j&��Y�[%$���+���n`�]�ǆ�k�����(�H�|�6�v��� '�ȖKl�5�E'�>߂c�,����V������E�`/��m;�H9��7�ќi��E�ؙ��,k�1�	zE�Z���@h���Z�����,�)�NV��q�
}��#b^Rh�3�H	A�.�3�T
�vyv�0/f�9pO�~P�BdS�ɺ��j�}�
��8�e ̡4X��D���9;��1�L�흮�ag�C��}�踕���5�Y�p8��r�j.U�7U���^P�Y��"2Aa�.�@s�Kۡb��r�9���a�k�s���qf�<�"�ʫ}��Gȶ���|��jKgǜ�'��u�T���sw���9��������'�S\��!�LŜsH���Ffo�D�&나��ޓ0D��������2�k�z�.��'<����&F�!�x|���U�W�Wf�4��a1��W����g��EMK��rTѮ�:�Cy|�����ꁹ'�Γ���S�и��y�WZ�.�p�4D���IG��sZhc9����t�-��w���H���w&z�҈��h[@gG5�:`�7�錊*>��K�"�]N�lߧ�iSi�0b�Cc�1h�S�=S�il�xz������ϦgN�u�X�޳���T5��̺��(���.�{k[���7a��QTl����Z֑uBժ�~j����WC�k�}9���p�_z��Uq��S��^G�{�� bfF��A�!����bC|H;��z@�j�T�e�"x��H�%����Uub�wC��)�hc�ʵ ����)��������q/tg!5��������n��Z��* H؂]7bk������>�� Qt���\s�F�q����O����-[��i9sث,"��q�륪a�Չl1��}~�C���4v.�K�&�F�0'��Y�g��cG�8�qW��A��r&`u|�o.֗{da�-�6�"/�@�C��p�赢�|�+��'�z����}�2�j���Ɏ�g�7 �����p�k���R�Y�� 6!�e*�ﶁc��
��T�����v=� GNq���s��0&��k 6�箻����64�７1�S\=��)�8߻Ǩ2fhŘ/h�\�gו��"�.������g�eXf)��.�s�{Ό_imx������	��4��>3Fn��zAhv�ldd�R����{��w��Kcb~'�G�g>�4��8��ݷ�P��B��?���@��;n��J�h�߫jLs����ڊ�"��-b����)qف�o=��<pO�V���z��ОT�<��*F�n��Q�^I��Q��L���җ;���ߺ( �Ʈ*W�nC���\U�#�A��pp��_�I�]���>�ŧ�3�_z������9�+رR?d@�b�z'Nx,RU:&��Ml��X�@�]g��=��Mqo8�\���a(m�o��֕��w�(`Ȃ�N�0:W��"o�&G�K΢��PW(�E�ir�ܢ!gj�� ��\�k�εJy�ޓC/�/U�%۸��iw�v�m8�ރ�u�����3��]!�������{J��3��H[ �H��z|e0�GȩЕ�Y��,Jf0��FA��dQy��sD��1��= $1��C|��P���7�q�dV�}����Ο2
��$�2�k	�G"�n����:v~&rh�lY�2�[b�۪ @�_>��� �
=y|�^�N�2�`;x��O���z-���1���ܔ׹6�s���2��#h�V�l�2l�5�����٬ |���Ҟe�{ܪ��̲I{)�6k62��*�)*�,H�M��N��4�d�	eq�x�c#B��U���J��������������[��c�	ZO����l����c�~���4�sZ�۫�Ѭ}+�J�P��m����|z����<�zǦҠjK�=��(�ZE*�RFj�;���@�'��r�7:�����( �F�O���B�YO�cY@�v'V�W��|j��������}�K'r�{a9pZ�:i�.�� �P�MgW�R,��e��*�2�X0�㇓��[A��{v�xQ�)�B�+�Ąi���=����1S�uX�Va�c5w�X�V�u=���g̰T:��H�����0��]����sv�����dX<�:���F��s1��5r��U����_�{�ﱑa��6���3 �nt�4j�1!R�:,���u��s��Y'�Ӳ3����mƞ{��'9��E�@In3(əKo��ɶk�d�o2X��Dv�y12ۘá\C�c���� +�7�<�.g����A�k-��p��e������&&��Ŗe]U~�x��_<_�����E¼)�]/b\�}3v�;�v��J���%�N���y�SE�����}��h����)���WM�c�!���Ǽ���y: Kd�*³k�K�Ra�(w�7~�7�G�|z��j�XYW�c�;x츲��B�W��W���z	JX}uz.]�zE��H����耲�.��J��M������SuX5�:h����u�ֺ�O#{���7�ڕ����5�u��|m��"ݽ�8�v��7:����R( �F�+�UZ7"��A��c�nn���r !^�lMv濙bQ�V��d���vГ�z�nU��k�Ϡ�pJ(�Cג��P��Q�:@HN��*���k��YK���ѫbuz�e������ ZZU�C�C���Ř�1@:O���l�
��b�?��_�)��4��(�2m0m�����g�9��V%
#U��2�$P
��@�1��l�G�uL^��W�OֺXoD(���haQ1��i;3��З��~\��v-�ru�.1f�S��,ZdD(��{[,֎��l��Q���؄��qrϙ!�N,��tݙ�����t0�E�K�������dp�>gہ��\{fX��8Ute9�
�GO� ���=5�9R1{yNy>W��^��*t8١�����C�]f��v͂��3�����e�����+vK.�Y]���sߖ��+���D'�1DCG������wD��vf�k6���=�f*��5�#z~�Ħ�V��M)7�}������V2Ӫt`���0o�UC��)���3�H���=��`�V���Yg�޿_��GF�����)ė���H���P���� i�N?��G��.���f.+D��^c{�hyM�ohCﶦ�w��M}���3�����z^���K+�*�^O/]M��t�����J/]�����*2��Z��9!;2;k�}9�[���� �aN�5���o�X�5��� ���,��_,�uA
>X�W�|�ICT��w���0܂�n�z�1gMƓ9�}u;yb�ľ"L[N=R��.�܎@Y,��.ޘEW^P;����N��.40hk���ڷ$h��`�6��4�ۢ��@߀T�uD���Jݷ�:fcv[nha�q�d�H�����Pz'*튮��#z����7Ů�zk3hԩ���0�*���Ԕ+W/,/�!���+]�#���]�Ȣ�` �	
p��]{$�CE��*�X�~��B��{tMjsВ&�~R��DcXgV��z��"�2��l�a�3�3�<]3��z�U���U�� Ե`�B�0A=�n����XON)�#����[ti���!1.ن���Fֱ�@����=NլW>6,��� K��m�����X�e��я�{U#&o:ܚª�pfܲ3Bbͭ`W*��ff�����!\�V�0=λ����j:�k�ޖ�\�Z'�K�]���*��#�HQ���W�&l2�l&�,�Ě<3���	P8BH�gW6Y�Ƃ�����a��h}⢄�jγQ	p�}^��YD٢�����CG<�n��k!�ݛ�{�Ζ�86���ٳiAa*lb��6��N�s�Z�� ���OC��;�Ÿ���~!}�?(1�������[Jm_]ZI'�I��#��4���"-@�o�^�G�.S)�kLU�WӲR�;d�~��U�&�t�N��.i�&�>m+����t�i�؉4<�H=�;;�Щ%�m���j��64M_�������߿( ��F��j�"�ˡ����*ڛ�k�D�|i
����.9Ț/yw�����ô!~�.f�PJ�-�C�Y^"f �FD@�B���om���ڵ#���{Mяǎ6j�X�]�`bWkڞ���-C#ғ�G��r�ⅴ�^Qd���S;�ɀ(�y1%_�o�T��*�d�Z�oto�>�y׍#��[�NO_M�OO�Kt��f@,���
5�A��W��i7U9\�!�ٱ�rQ�и����-̾H�	p��.���dG����U�0��"k9�ʑr<7��f�SV�O��S�Ք�&FN�ά���Q��?YKE=ܜ=Vμ7?~\;�%i9f� az{w,v��7�������-s0��x�Y����"kX+^�|��)��}�Cfb�#�fM������;�
��53K��c��RT��[i��l���0�1cn�&��܎ۣ��}��F�sW ؙ��]0���A6+A��˕7��g�:\�bZ�d{J���o��oN��}�e* ��S�BsY�o����#���du;�������PGJ�%}sm�w����!B���g>�~��~L�X�;��-�++���]bnв� ��U]��ŋ�
�t�]w�!�η��ѣJ�2�h�+0pb̯^�I�
���t�7Ž���I �/�=[N��,�7{媎����oJLx�*fh+�6WӰ�*����Ӓ�ua^=��6Ԭ�G��Rw��N%�KȤ^���j��_�( �6H�G�	�uo�3��W��p$�<�ηS�E���T�8�����رq�0"��8j�IU�Tv����~��ZY�0�k4y�1�D�����p�Nd@�ܢ#}d�D��Z:�w��}�{M�gMC79��>���*�߶��u�Z7�f"B[����2 bAǙ�����Kit��n��Q�`Ɉ!,{�`��c��m�h��-����XiQ�r�]���p�r0R�11]��zk��?�i���Ύˎ�� Ӗ�qe9V�l+����`��М����9��q����}�;#�l��r�^�Wr�^9J�J���6�`�^�ۀ�'6�T`C�0&�	.���������w}�w�f.Qp3�$���x��y�����[;k?,Snw���7O��7�?���@����-k�r�0�١!�6�fi&�o`H����|�ؘ�ߎ�̡!9���]�zw�_��#�ߛ�������Ӯ+�&��0<W��|N�@a�{��y�	��ʛ��}��;p�������7]����d�Ǌ���/\�ܿ�[��Z�%^�银"@G6�#�<bM�7~�7��h���F��6Ŷ��ы�@E�]�1�7���@����<��X_z������ϷZu�s�lR�gGzƁt�������l35S���k�4���}�0S&Zss���#�z-���
����Ro,lD���� ������]`!p2���%��xs�+ǥE��ͺ(m�U^��3�P�:����'ӷc��p���Jt�'�� �����Q�P�����*������_U;��x�0A�D��13@q���bސCw:���[�
{ 3+� 9N��`�^N��|_z���ipX;X����	�  D���3�K�Twg�!��,�`uwm���[������p����O��?V��;����Ä�e��9),�x3*�ŎW;`6��a����lH�2��-�}��O���O|"=��fw4��w!ʪ��+S@�-�P���z5���$�sc�X�C7,&l���[^I�|�C��sߟ��m�e�t�^�K�.�^���Ei���xv�j�|�v�L�g*>*��� �(4CX	���ރӥ�p���59�V��|��Z����`�ٜ���PS�I��n���tp~�#j��mzF��[��*�6(M�$W� d�E��^���t |]\T���(�������.\Z�3����y �����?K��P�z����=�q���}�������[f��U�bC�u���[�w�T:~􀚪Ω% L:����sS�;b�-���v�jg�3@���
�i�6]��i��1b�R�C����s�!����O�m���"	z��"L�X��?)���Fmg���e�&( ���sx,ZZxs�=m�<���X�_ ���_Z���𲣮��)�8s.�~o�A�'4 $x�i1����t�}�Iԧ�⊳�ܺ0����u�2*}�'\�g�ӒRsYH��k�&}��|�ŨgN��uf�s��ώawW�P��a��w��E�ŕ��
[9�xo��ᵤ]h��[T}��j��#_��`P�KQ�:��[�ȶ𢻦ٮ��@C{K
��`����w����ZD�otIPuݙ��3ϺFM�N��0 ˵e�c���,h��xe�;��4r
�y���4�GB6�����O�9��^�v(���뤩˞.Pɼ�ޭ�i>l���}�]�/�~&��9�g
�����Р+L3';|�?���	q'+mJ�-� �}���+S���#�vɀ"_weF��Ie4gR����	��^I�o��t����ҬCG�����R9�����ML���8o���f�w�����;q�Ҵ�9c��c_L���Z��=����^ �J���m��	�X�j'Qu�LP�Q���V:
�nT�G ���s��F� A�U6��r������~��ނi�c<K04 �?�?��t�w�Y��B^u�J��K���+.����w>��i�Q������1�����Κ[[k�q!�F����W�]��ӽ�ݫPۢBi���Z¨�ز:�SChyI�[5^�R��rZi����v���ꍸ����i�ʹ��`G������6�@A70��o��;^���ڳ���k�������@�|c�^��^��W��y�� afK���%6[a��dĳ�8(T�D#�LiC�9���#��8d' "L��P�3�d}rT�m8kI.i���l��_x����w�ig�vf�lvh��?v���v��b{��bQw�����By�f��[o�9����w���?��:s�t��N=�}=�B���4��Q23���W�A.��5y�����,�n}���Jw�f�SO=���������-�����x�w�a7�Q�{"ٌ�Bt|m9D�ٛMi �4+�O'�˯�z����OX��cv���-G�� �f���B�U"V�-ɺ9A�+��)\�:�^�������ΨH�%�|~����������wλ�T�F���v�0f�=Ö��"ff�~ה�h�Wd]99A�0ٺ"�b�������x���?o��o����!�=}���������ܸ&���A�������Y���Z���a�?�����J����t��)����+�����HO�8��`�t� �&�@�wg<JϷ�Y/�\�~��Y�K�B!����N�^�2x�Գ�6�����Q����|������~o���|�����=�d��u�h�Lv�6<���(�}4�TK�Ad��]��Z�أM���\�j@!+͛˗.Z�`FC����-��r\ӈ ك>�гt��	����t{��J��Wl���}�/}ʎ�@�0�G������� Ͳ��?�cwUu�ӓs��f�����` Ex�
�$�$A	��������a209�ι�+����}v�3=��L��?�z�����>��{ιg����{7��L޲�o�6z�����p�?���ge����A����w�r�P�Ŗ]��r�{sq5��X�@po� ��c�GcPŤ��®ҡ� e�Z�>�b�2`������V���92@ۖ�\c���gE��ػ��U��H.�}j1���pQPv�ZV�n�x��y������c��򒗾�|�/?PN:�$-��eb�ds�w� �����iP���Ge��
������Զ�2�~q˽���QI���>o)�׭.�~��ʕ߻���������m`0��7>���?���n)��0�O�� �ņ��н��/�+amy�{��0����1~ի^��o�fRk�L���njdD�8����$�7�f_�%C��Epޣ�>�;�O|��C�Pٹ{Yѷ�<��*O�姗/}�?�"Qe�"jǟQ�Z�+�i�Z�iD���dL9b   �)�	l#��)a�Qrý�o����7��|�ӟ.�wn� �����Cҙ(�7ŵ<���܌$Өsdcj�`	�yWb�v2�;���c��s�5ה���_�˯�ܺ��=����xy9�Q甯~��:z���M���;٧|~���9_y����F��������]��� ���\nP����9��{��_'v�!EG�	L7`��)�x���"WW ����ϻ�ȕ�AkƆ�,R���}�|�ӟ�u��Fz�ﾠ<��Ow�����7�7e�r�0��D���Sc���zѧl�\�c����G<L����>�պ<~�[�^�֐pѹ�46���ͼ�����K����� �� }`|o���r�-7�1=�]j����A1��{U�LݲO����eU��H���vn)�z:Z��̝�7�y��̎�_�;�7�{�䁡Ѯ�ˇ%؞�Q�f�=oko�
��sV?3�9G�-]:%	�)X斞1�0���w���90H)L/k��ŶM�)E�Y�ҠiV��g�:N�d�8��uP�]_V	��	}�ލ��ض���.����ꁀk����	�%s^�{��u�гkqqH��N��Hj��EhQ�"����"�� -�]��yR���{`��q:Hn��kWy�w�o�;^�6n����@�>�z�a�)����_�0u@�1Io{��yQ��<X�_��xg�n�7�,߁�O��l���^w�,�\�벀��q���AC��7)eㆍ�������(�Ʋa���w���q�Y忾�������Y�%�'��,0g��yِ�����aCW't��܉��-�|�3��@ h��QY]^����a�;��������]u�gZ3sZ��l`�6퓼��5���6�ȵw���iW�x���'?Y>�5 Z�r���}�s�)g�,W�x����]�I�s�2����R�8#\�b�9���k�d�E5~fA�
�x?�)O)'�|�������s����r������=w�`՗�a#R��1�Q� ����O�>i��G�t�l�pls����B��G?Z����ҫ�9��򲗽��Y��ܦ�y��u��J��2A���P S&l���.��VKP�X�:>�3=�.��2��8���EP���-��|}���?���=��e��NLC�O�A��M�^}f�(�`�������:���7K/����/��^�yĜ����ny�����#�K.SD뀑��<9�)���a0u��H,{�'�sĦ-t���Z�tTEs�ca�����j^S,��DX%�L�����i��l����,��T��2�	X�j�-+�^zi�v���7/����S��KK˃�z�X�����o,]-�=m������ۚ������ͱ��M�M*tR"r��5���ԾwF�ш��P��wN F�;��թZcg�'iV��h�פ���r�c6����bKZ)4;�ci�d*��tV�lLl�>�ߴ����;{P}�P���5�����/}�.��9m�O=�ԫ�>�+�CM�O�� �0F|^c��P��{���;�{[$�������TM{��6<F_#�K�Az�F�(!��wP�n6��,�?�9q}.=��d}�Q�%�d�|��֮�B�{���Pn��E�*���b�0�0�$��A���ǜ��^_��W� |�_2��7������/g�u��$cs��+|<�m���*�n���
��ݥ@VÈ��}�{o�R%���N?�m8]�������=H�y�\ ��B�Y�@Ȼw� b�Ƅ�h��~���XM�U�N�K��q���x/��r�]���w�׼��e���2�������=�l:rS��5�h�骰��1}���_C����#�������� ����rĚM�w����W�W�9��[�̦��B���d���_A(�EEe���qM\n��	�(��E��42Z�bæ��S$�P�z��c�)���3�]��������UX�𕯲�Ρ����sA�O2��u��'P������%[c'훘+�͜���`�MoWoy����x�+���!O���;�0� etW^�=�9��w��R䍉�B����R��Ѳ}�v��?��﷼�-n��뿖e�׫4Ĕ��p	�O�*�n�p�gA�y�Щ�c�o4\qfv�ϸ����>H��s�����?��.�eT��]��qDs�R%���r���[��5��h�y% �V���4����l����vq$t$�����:�`��� �y��Kӽ��%���=9W�"͇k������H9B�չ�>�\s�5嚫�����	
��9X�%�����꯾�%e�e�ms��g'$�l���kmk�`M�RL�S�}�\��w��v��ܬƱ�t ���Ҝ�̜�g3��3���xN�����]�6s:fN� �&m���� ~��zf6�75����Nj=��'=��#6m�������}����_���0��O�WA�����4�zḿ������{�EŬp�n�mz���U�'��~�py�cD�G!�3J�7I�0��X8-R�y��6Q6��߹u[��p�)'I��;|��K��c��I�T ̤�\nZ�"��6U�W~ �R�u�7:��Moz�싾s�������򗿼l�$���3wև��7�\�<9ћ�w�t/,��;L�������_e@.��2kN8����w���r�)�[n1xs^��%8d�%�^�}#�<������#�wja�'랓j�;��)*m� F��IO~�ټ?}�[zv���ۿ+W_}MY�c��$C��z��  z/rN�d�</ݤЁ`����X�p��6Q^�◖���۠n��b`y����o�9���.J
�6�~�H�9	�i/��ߓl�e�&��dKg�FRu  !*�2�j0D�/zы��A�>=��o~.�k�xq>�~>�^.�&��ZTXs Dx6�,=n(��M7��{�� u��@�s�����?ݶZ�x�]�����Q_�:"��$ &z$\���G���Qn��A.B���.�`�φ�we��|�Ϲ01�_jX��g{k�2�9�b������?�s��t3[��J�2(`@j~�8�21;�l�]J�1w���r����+���kָ3��v�~�DKp3N��]e�`�p�"�_��֖Ve��͑
�Dݢ����u��?��;-&�r�U�/�vl-S�=*��?���x�1eǖ������\d��Hͷ��+��ڿoN�[D�4�uv��u�x_��5I{47�bE3A�<��rF��Ts*�ɵk����Ӥ��\��m�C}l��S�6# #��J7��A���o��U���9�E!��a}4�N=����O>�G�����M��}[�]uǌ�ϯEt���b��$R�i���@X�{|)��=�?tq�/&�����y��ު���3㢡��"��t�@����9+��E�J���&"�N��f��M�s�N�u4����B��%���+F�W�1;��2��A��-R�<8(��}v�K����b`q��U�Vڨ:^�җ�=����n���VLǰ��a�%uR��
��I��2(S�!l&[�������Z�I�v�j����K��h7.B،FÖ�+�q��V�)�b�������q)��(�1�hX��*_ Ӥ�\y��~����������f�?.P������UF�j(3p����M�V8���r�/�vW ~"j�E��v�1�KUy�촓N���V~�)?�]+n8�"���v��A��L���E�6��(q��\��]��=�E��Ι�X� �8յ�y����c0 ��8|p��)T�&���|�����=��]�Q�t��oZ��
�ݤ�C�D� �I��a���]�l��K�� �
���ҿ}�u� �,�Ò��}Fs�%�����W��k�q^��g>�:\��I~�(l).j�W!�i@��"e$N����=�صx�:�X��|�7��ՏU~ƅg�1Kw�-��O�y>��~����3�>\+F��c�ZX��o��\|��z�������[>���T����v���� �Ѯ'] �_����_�)%q"����g��eҰ��,k�u�c�*M��u��zB�����ȁ��n.����̌�<�]��jͪ=�㝽KF���)Bv���D����.���葇wfF �S@��j.��y����O��aN�O����j�Ӧ�jQ?�h l���6������S��K��i�jW�~�7B���u-�7u�c{����ƢYk���'�x�>�G�C>_A����Ԣb'��HZ���V�k�w��K;쵨�'l�yy�3�d�}�B_Y,��1��,..@FwZ6e!�H�ء�|� ���916�ZX���.�k���Yvn�M#����2
{��uJ�=H��=��`�5F�6�rqӈ_��|���[�������W;] z�$�|�+^)V���;���ZL34=��Gu�%=J�z�;^���Y��$��P2�#T=�"�9]E{���4>��L��駞Vv��N�pT�۬E���Q��ɇD?�ֱ��q�ӎ(��;Z�,�d���C��:��(Na�P�N )��s����/~�\w�JMp��ĥm�;�6� ���5+�8�>B�N�U�)�Q�"/�� y��Uv/<��s˳�9��7+�x�4'\����-ޠ��2D���u�"MIv��ġԎ
�t���pM�t���U9dd�	E9�.�j"�RL��0�-�H2��n�Zz�'sSOh�`	8/._�`�hDJ2/ �f�@̙�#�U>W�'�Ͽ͞�?\�������D�x�1��nW����=
�)U�9�Gf̘/5h 3fG�e \���ah�������@߀;���/������1�^_�� �+�J�ad��H��G�gua����U
@���ث�ӹ}t�۴� W��MG��Qcܛ&j�m�_yy�=�q���//;u7����/~�<���v����F$�)�x��6�M_̨� �{Cr[�M*��k_��ǋ��㞻�a[���w�܄�Q���t��^m�Vo(�.�:x�ƳM9�V�9;E9��^��ѳN:�?����(|�U?���" ����M݊xY�U�����?Z4O��m�{V{}$j\��q�G�9�$�����uz_O�^b�[�<�]�ڪ睷c�B��	��t����3N?}��������v���zFv���s&�� �0�}fl�yv�%U�>G�y!0v�'�C2<
cB�{�X�Bg�lR��o��g���qP"1��5! D(�X�v��e}�on�
	���U�hQY"��Gn�v�
�2d����d�D?��*C{����yO��3	�z�����S�l]���b�^E	�
�/���N퐹=���TbqB�D�!S�j+�vьLkGv���)c�F`��J�j	i�c�B���U��->�]e^�CTvC���
mN R�����R���qF�x5F�y���	'�\�ؼ���k"��KYF({��([�f٣�b�����Nډ
Q���ݸ�?�o�S?Kd;.W���$�,�BH)0�62:]� �}h��N\��1�2!��\;� �qjfL�$ˮR���Q_H��p�EA��aZLaP���M��'�~X7��Ssc��fRV�=�ɣ��!�9� ���9�&�H�<e@?�L�o:e������H��µ���� w��g&L}�.��ф-"c8O��;�z,���h��sB�"�:�(1f�`1e�f��Ä[sR��V !Q6�9v�Sa�sN��P����=�r�F�۸360"f��'�`:��J���� �=K��$������4�:":;4�y�?�9�[ fV����/�^��%�sP��nX�	���+��,�˗��;f���@��Hխ�b�zB��2���˩��#�]�����Ĥ�}l�tܚ�G���{��}s��f���G>�a�B��G�{���|ƕ�׷�I0���$�mry��R�h�	x�J��lE�~Vλ 1@ο"�?�&��n��N����bug=r��X[��i�*]☞�Y1���G��L��ڴ�����O>�������=��7��b��������)?^-YA�1^^2XP�����Q�ÀN��W�1L��s��/��4�\�ݻA=�*��퇗`J[��(p�\Om66M��o,���&Y�� !�J��z��`D�$�!�2�C^����.�X����)�9���_��UO��ya� ��;��^v�S C-� @�!@�����F[ �@��	T�TT�����DG��3U -�a#�r�ɲ���� T��-�U9zB��1�b� ��w �����e7
cD?��r]-X�H*�:�_Z��ႁ^p�jk���伄�ʘ�=hH��ف�� ��9�)�׮8�(J+A�����
v����+�������zFet8*�WfmWh�  D�*��E�� �)��U��#�{D(2��
�{ڗ����uyk0b�Y�䅋C��G;�1Ր��k� ��<�Y/�$�!�7��Wj�RK�|������Wf��]�ʢ�p/�V�x�`�`���5�HVI?��D*��j��!��z1�R�!��}	ۅp F4}����   IDAT��ȵ�fdTc�ry��^�Fw75��;�^|��fLp]Პ���؈�pw	�;j�6=[`3@��*��ȥuwII0{�x� �������oܚ�����C�neEV�!s2Q�R��{��r�uוg��3�G�9c]���[F�}���z��o�V�'��6�<��1�	�A_f c��g���z�-��OQ��Xtm*�ڶL�H��jF�R��n��!�<5*���1a���i�Etx#�U��^��=T�G]懂 ���R[��yJ������E�l��ܦj�]~�wV�)���#6�n-ڰB M)9�0�x*fԙ��EӋ��<��lU4ǔ.�#�٥Wy7n� � ?���v���Z���(E�C��%,~x3Aj'T>fT�����1�H��X�7���N�|LA�����Ź2C�d� �%͈@�%b���n��ϫ>�4��
X��31��}UgЇ;���9S�l`-�/t1$�P�bIg�Mqo� '/ra��]a\&e�ڕ�������(s�.��.�5��V��)��T���R�R�i4[�5�Co�9nڴ��OZ�� ]�I`ڄqI��1��:��=�r�`g�y7*��W5����$�Б��"q��N@���L����H6��*�M�V���H<����R�c�oW�����3��W��6e"C� �k 3�U~��7��|j��<Q(4�5;v&x��^��C&f�I\p��H�5�H�hw����(N+�c ٤��+M���:�MJ��1��pa�6�9?�q����%֣9��(5��`���q� (�sb�`�j�i�	��}=����c�z%�~X�� t@-�l��w��]J�U�n��W�������t��+N@�7�c0��'c\����>mtT�L�$���TG��A����kS�T=�btG���J�g����e��yj�Ij���OM,���j-bɵ�xY�
�K��E�*@��,�;w3���šY�F�A�;QS��y~AeaܿOy~n+�u�(�E��P�w�X�(P�!dmv��2;�V�,U�V���O>E.�=1E���hTK
Cc�g �A���Ls�?�7���QUH!$!�Љs��
c���*C�>��]O(|��a� ��!w��\*A��E�AuX��̈́l+���#�#��� h��4t&n[�l/ ��$zYl�(t<�Fz������b��B�;�\�Ղ�̑7	%V����>�63ЙUԞ .
>�0��;-s�p-'�������꓈`���j�"��7s�[�#�����p��]�� 5��	7i?�����\�Quj+F��r�F��5�| /�4��0KT�Q������)�Me0��Y.����l���{����@��!��Z[p;�!#^�e�
j�>cd�Q ��WtM�7�3_�$��"b�dY�|f�L9��g��.�M8�s3�d�Ft� HZG�;ˀ8����O!h��2ĳ��sTm�L]�w��q)~��D��h����?�Dg¨�Zֿ������� �c��.f�6>KNe,Cbg�����Tʊ6��ڷ3j���S�	��d�O!�׵a�xx8��vɅ78>��\*�*h�
$�+^�_�u�-R�6&�Z��:���e\l�"tv������q�����kA��f�\��esa?�74.��vM,SdC��creQ��u�Xt`г���c��8+�* 
�NMg["��O��R�^��[�k�+�߫Eh���Ұ��=h�u�9稀��f�>��ăJ�ȇ��A~�[:'׶�cgk�1-h�0��@�C$D\��B�6j]�����6���X ���@]�C@�I�&��aq��Q�X8�}b����:�� ���rn��	�<�\) *
�E�)�^�kdHh;fG���j�7Y��?�`?3�*�dd��R`P7b ��\]]h��>��U�dUG�2uR<��G�*v�$���4�e `#��耘r�2�H�QD�ъ�Bn>�3�A�̆���`4��0�#� ����s�|_�W @����>G5�97z1oH�0����{�KLFS-����V&��x�f�)���B�X��G�D<�9�ZN�5���=��,�|F�6�XW,ܶw������y�{N��?�Y�{P��������w ��abn;5�cF�����dA�J��/D��f���{����u�y��p]���B�+��&r��e��AT�;����R��]�g�7�j�w:ˠt�����:�+q���zmJ_"
�+w�A�?T����D�Vvw�9�GA�)#���K����+�vPE�>|%gT��4qm��p�)��@��Y���1���>��䨀��T!¬a�5�t��C�էr����&�Ώ�Ո>��\�~����%�5��X��֯3� �T��������o{AA����'ѲY9Q���^(fT�͊�K%]eր�c�*�B��pW~1�e����W
���CJDYͫ�r,�a�c���M�UBs#���Y��f��h	��]Vƙ"�0S,�Q:� ��6�8\�"�òTwE�؏�&7�Nh 2���F��;�9��DD�XlЂ5�}(�/�~`b��Uf��>c��3|u��ZO,�5���n��*��
`��]:O�Y�	��F�[&C�.2��0H����E5��w�h"b'Jm��2iWe� ��qz9��3ˊ��cB�	��,�;�GbS׃�Ǻ�`�t~�R0K�S��߰-�:�T�h���b^h� ��Ɣ�w����s�έ��;�,Y�����TjT��L��k�z1@����{�,�k��u�P���4T�/A�YT���Wd��te?�3yz�h9j�6� F�8���|�M��S��A �% �ov��� I��c����Iͅ~�����0��d�&!��ilzڴ9SZU�P��߿ҥY~��^~�!g�~����ʐ���t������3XfO<�w�QX XZ+'�p�O�jo&ꆫ]s�����<�S%�n-��8P�$����UR�A�16V^+�v�6�U$E-Tg�⯟�Xd�k��(�4�^D2�p����#ռ&�����s����RP9�p��h2�щlB����p��Y��Q�'D����17& �b�M����hvh��ѰvSc��Y��.����0#����d��n�ܒÆ���;�&+D�c�Xܜ,��A�~���H_�F��04�F��"�J���X��ŁB4	�#r	��H!]�*@Ӏ>B��Z7��ɴXڸUMNFq��#D@�T�
#�9Bۓ!��Vm�����̔tOji mD�0�� Ȇڠ��6�\+�0����`E¥6_c*��0q��<��"�3�^1��O�������Tc0�G��864-�� �/ے�@#�A�����s��xL9�3����>�le�~Fy�C����U?i������T̃|��$t?��C���@�ܟ�j�`��B�7 �v��X���>��H�s��{v� ��EϺc����-:3��x�8�ɂ�
��8s-���v�����Z� �lW^��R���&fs�Ϗ�Ž��e�ÏY<~��&�<�w��9�!�ϱ������:�(��1��h��hk���+�?#GV@�k�G�o"��3?�ĉk��g��qY'�ED�w�����Qf�E����ٷ�������;���u�l��)�o�6_o|���:q���8yS��tp�6 ��LoZ�|�e�����L�a��x=�aXb������8w~���Q�>3���nl�1%�z>�By0��ڧ���V%�ӂG">rgP_jRB�Equi7�����o��"0�]��(�� Ǯ�X6(�F�v\�Z�o��z�v{gժ����B��?FA�\_�x+��	�ɢ�D͠q��i��+� �=.*�S�W�V��G"�(��ϵ1 DFQ*��M�@;<B��u>tA��tYv�Zxq1�y?.���ʈ�CV[:I #J�ȱ����R�&������ �Q��������Y���dd�]�lPB|�g�Sʝ_ù)�}3�>�������B�թ���i�7Qpɮ.�M0.�����W��>�AAה��]�����zֳ~����,b\��w��u���!ȍ��z��8��O��&��n�lG��1C7S7<��TG��P`w�\qI�-0I��}�߸�E8`ڭӍ�g����� �pfu.�gw\F<��������آ�0���>������3�{0u@�����y���n��'� �����%��Ч�b�f����V�*.aAz94��/��Y�k��~�Ck�9�O�������2�3W����H-3_�a�Q�eY���UB�%��-�il��6��P��1m@
֗���kZ��r��c{H!m�Q��� s[�lw�@g�"�(����\�a�"Y�@�M;��9]D�G���6"5FԮc�0W��4��^b���|���{`��k`Nq����@���b�F(F.�C_���[s�t��V"�&_�Bx�|�$��M��ain��cnZ��2	͠ȅ�G���ŤO��֞�t�r�vlDfj��L���)�� �����=u�[P�t�M.�� �*��;��f�%��,S�� 
��_��`���C��CaF-zYu>Y��1��`\P�D��ygN�&Ј����Ε���{\gXf�}14�:�$?���'hS�IjuyY3#k��P-R�a>�)�A�[<Z��v*�Q�� �\��ţ��0�f}%&�ς��"�P���ݔx��i#��(n�d�<O�6܀�­���|r�Ufʺ��J�=/>�9��tuw���v)�����#�OI1o���S`d�4B{��ا�s�
��
Q
�΃ԃ
�-yoЏ1ga��p.ړ�&YϜ����VkV���=�7P{0R2�
6�l���n* �Ne!87mc|<_*���������]&���\6 0}�{0Fzܰ�A�����}Ŀ*�K�i������K<O�����[���Rq����sM�z~��YtA�o4a�Hh��F�繃:G�;< �ni�@�P$U�zFѤ������y�7��DGح�oʬ0����QE�H�P��ܪ5���*��D�_�jj"�Q��ŵVe5V(G���Q��K\>*P�u�H:ʆ�/��/����7�+[��i��%߽����o�{Ri֯�:�M�XO��i��W�C����*�a�ܤ�aQ}v�����1- A�e�� -��� �v~7��hr�]j��3z�[Z���%!����Eƿ�#L2)� �uƴS�P��
hav��ܖk1�x�á��	�C+��P�
�w�$�h+��VX�a+X�X �QHS��I��|x�f �Sp D�2�J�n ���)��^�2�.����<�!F��;zYӣv��.ڋ� ��v�2�b}l�|�X��F�9ޠe�����6���S���8C��vH/T�C�R���'��5�@�u2:!���]dc�v��v#�R����W��V@�q�0�w=2�����K�M5p�u,�Uw	}�c<N:�de�]Qv��D����]|��v?Ў�ڑu�	�� c0y�P3�O�bi�Z����4� ��(���/�G��e��p�Et!�������-���i�) �{>T&	pD3}ܾvӆ��� ���{jk��h,�1�m�S���(8�+��s��]������'�#}���XF�`P�%�\�VnB�c\��0��i��&ɜ���(L�$S(�n����9ah}F)�C9�K�tTnz��s�A\�����q�K���,]��c��1\��F�"��S��q�>p����׿Z�UY��N;�l���T��%�sܹ���i��^�U���O���L�a�q�5��� E9��ٛr�vd��§�"3k,����-������x7It�Q*�w��%&C;+�o&�9a0��D5ô`Hud��9�X�z%T�i/w���we��~ة�q����)@C��Ek�Q�0 �s$���8"Q5��Е�!A!��@N��j�$����ذ�"^�%�r�Ο���~5�DSm�"���5��zA��1pVae�G'��)�$?�#�H��@*�^�:� ���Hq��pof�zlӳ�Ny�r�]��iGc���d�0Zb�� ��
�ŘQ��A�<'l�j�=���l�LP9'����f9S��	��5D�q"b�\;M�י�f����nL�<"�&�t�:A���fX�2�Y�9�h�6B�q�!$W��.H���V�l�����0ٖԝ��rm.�O�ie��N@)Z�Y�ҍ�&���!A��鈢�3�A�L-�j�+H�K ��� s�9�9�kOc��G��(?�ju'1ޞ�l"
�MTٚ�g��-D��Cn
��� �|��7� ��,��q����.���l^���*�F��1�ٲl�
�A�td���SD��t0��g�Dmt�I��XJ1�&���k#�W�r�맽m�#M��`&���k��}��R^��=_p�M�h}p��&r�0�~���%�������YH��]�J����ig�����+����v�ª�h^ZK��pZ�V�H���a؊ů���E&�0�F��)[f�O�燩i�y�#�8~��3��E�B-����4�;X��y�aт]�8Y��!�E�L�^%�;���S�-��z=y����%�G�U%|J(�(�)e�V��q��9-�,�$-���c�,7�~��ګ쪚�a��Mq���ʡ3*�t��˪�8����C����ۨ[c�����;..m�\���~�G$� ��(2@��( j`��(į�J�\2M�H�@6�ӂG��nh4?`Q��2��ԧt #�UvY�!M�DٷG�?���M(d<ht��"�,�unZ蝹�z�wg�� �@�v�wы �e7�O���@?�B;y�t�l�1�'��L�5\�������%�:ҏQ�+`-�#�*s�DԺ�i�S�ש����<4c���n[�'��v�C6t��k\3�i�	�+D��oGQ�ڙ�M=*�:)f���9�+�U� cءy1�Q�n��Ʋ�e�-�b]��"�0���,�Mt8bdGj&��Y��"�
(Q���p�.�9���'�v
�G���sűT6Oc�k ��ѩ�J[�9�v��<L@�����^�Q���%U*kn)��`��fʣ*Κ��'z�ρ3��(g���]?N����O���eY�̺����$e|u�V��c���p2ʇ�Ϙ���B�iPX��SJUt)��ʜ�ɉ,%$G�?���hS[ft!^̥p�(#���J��C��5Qɞ�1�?�3{����h���m�:u`�6�"����J��m��l��2��5��'@:�cg4���!��Y [[7ͭ����|�\u�b�����_�6cZ;�` (km��_��Y����"tCV��E@���?�U0UmKLK��;6N��#_�C�r�U?P�5���~�g	mfW�,�+���G�0���"����
p�����Z '�e�t��n�#�Ԃr��7�uJ*�y�rb˦ҹTQC��3��j���阘����K:X��]��!ؙ��c
�5Ô���Z$���J���~"�0Y�#�lZ����!J�~��+�r���iX߹��ۜ�xRmb�O
5�+���:"a0�>oU��
��a�yj-MK/��|���$Qi�y8F��mD-���o��5�G4�!�˱*.�<�.�ta��m"W���2ڴ���:�0����M��sN"�y�R��GT�D��n���@�N���� V`킄�r�^���p�`�Cfw������b`���΃��o��C��}2�d�$ÈA�~����w�v���2�����$%�c�G:_��sϹA �	p�n�f樒.��� 0Y\���e����؍�)"qxչf�,�� T��b
R��V��0����"�>�aD]�T��}f� �75�-܄o������=�F`z(ܘ��� 70��bԩs�c��)� E����1"!b���#�$��fb�?'��6�a�**l�u~�tJ�]֯f�Y�X�)G�+�B��Y	��~��)(�"�̳�<��q����5�;�s�u�63\K��`�d��%�p�;E�zLl�n@{�Y?�_��j^Sό�%A��V#p`�D��s&n͉�Q����R?K�D����W6)O�*�ؤ��ގ �M��B�wsm���(h~%���c�	:�1�3#;y����W��`��Q�O���7z�ͺ ��]
A%[-�r���~�������}2R}�\Љs�9����ZDHH�S��]8:%Hm/va��٨v�-Zغ�1jo��Of'�5���c�pQ�R��	W
����h6�� �R!D4$�cwR��ZA��'�oF}
r]2��q�m�U�Ͳ蜔1��i�\d�-΄u��w�[��1�\����PV�n�͆���2l�!���C��mAj��e���F�s��`��ϺG�H�?`� u^q5���9��K�>Ǖ�¡�J̙�Kb��7��Z^vu9^Cc�t
_��YֿRI�-~��r���hǽB�O1FU�ù87�����Uv#���Q�*���^���hG�D�	�F����ŋc�$���7�ol��/�����4�8'ғq�ֲ�o��׫,�$�L�0hjeUw>�oS��: ��L�yO�$Μ?���炙+��6��q��w�¬ߕ�t�'��o��a���8�tK�� Y���f�D�	�����2�ų�3�s1�VZ�铑�9��r��Mб�]����7��-�ɑ�~�j����y�`N@��qk	lV��2�Z7XwAX��[��U�ݴ��a%�lW(�D�P�sb���P�VT�'��7a�gt�ܖ���ƤGnᙩQ�h�V��Ea�K?I�/2A�9��_����B{����c4�@?\��b�w��6��8��&����v�h2��[�c0<c#���|����q�������.D�*1�*��ev(�<�m2�=�ϙ*kǏDQ����NeO��!�Ɯ� ��ؑ�1�Ckbwn��(�Y:���	$�c�ć��!��.��n)D�S���`���Ϙ�b���kW{!&Q����H���е �Z�b`�I����ar���6�3vd��+i��7̂� $�7bC���V���^h�Bf#�P�0İY�*�>���@PlND�D��S<�� �=Mh������P�fڕ ���Q?��q=-�3FCͱ�/m4�P8� 6�2�YS��ͰX�O|�S2t�˙g��q�`]�F�Nن>���_���__��A�KD^��y�J`\���Y$.`ˏ50���lT�K�1O(����)F�c�`~������ �1�.�u�p�dɌ��m�=�����`3�#�ŋc�K	x������fD���/!��l�*��|��
�׮B=���	�b�G!Z�3�!��������f���g��V��
��=d~,�h�c��	�0����M�RIV�ڼY�;����;����kw,2'{%wW;ωj}�/W��и���ݽ{�ֺA1A�c	 զhQ���>fX���k��}7��Gsp\�3&'��5�m�f(`�����LA*!_��fz���ô�?N__A�1Zf��Ө��;��!��Y����.���d���`E0������� ||
q/>{��T�&tW �?�y��=Щ�1�z�c��\+K���zbRt��9LRE!����{q�`gE$E
���aXj9f^K%�D�aw@	V�
NG��&��Ν;j�
n�������85�k\<�d��AY*&��0`���P\���4BZ�%6(�@�f��U��f����axj���z�[�b\޳b�M�{�mF���B�@�����d����f�N��$YG8�C2���O�+������t.�U�Q���w7m:� j����O��Qd�>��m��r�^hI���Hc���b@с�������v�3��_?��5;ˉ'��H��va�����_P.���EJ��d�0� (���(ے��1��6�$�\x(sܦf`����F0����� ~�H���W���g]��B>�f;��2��(E�W�l�D�)�yN6���^�J���Pdr���X��8�0���SG��:^v[R)����xڗ��X��AU|��x��x���/�LF0�d��O�!^v���s3��֘O5����� ��iLp�nX��������v߶us$U���L�p�w�֛#�?AA�r�o���mykY&`�k�N�X>;wl0"g�)�	F����C!�Z/n���#�;�t��*�PE���M�UǬך��K;��ZF�g�^Z�ha�-����� �0F��@̻��U���pe��ra�nd�~D�LQ��ع�aU8�w�,��4f%6���tT�a��$N9�$�49d�����1-ڰA��Ds�o(�t�	acH�?�4�-�u�^M�E���������H{���E��5F7��Q���lD*����k���(^ ����Ȫ���8��r�"=n���؝�;�fi��C�Kc �DY�m:`W�V�?��0$�hX�A|�E`���l�F1� X�FM��-��LP����3:#��t�ѩn��=�
���a�aÅ[�蜚Lcc������ ��A�v$� ���[т�v����c���0IR��40�N���H;}w�2�M �����@����2 @s�1G� ���6�%������ng� �x�%�:�&��Am�~1������S�=.�v�İ�蚍N�h��g(�*�G�j��6�5����'��s5A(׶��n�p�;����`'��c��t���PS���<uT�"�)�Xe�d���A��s�l��Ǽ�儕�5�8��)� *���R�d��zew�څ�'A9}i$���c'X{�C�ļa$r^�Z�������T�cWy�~�ERٶL�5B�Ӷ��,��~q��ݿ�ŠI2J1f�W딈� ڷ�?����b��G�ZE1�Kz`\;˩*�A$�)�?�P�m��i��P�}p/Y#���5�G.i-Ǯ��9�w��������1�R2Z�p�I-��2�����I��6v��H�\�x�d����3���f�hڑ:�X˔4+��yZk=h���mo�)�16�JTeG�-�Z|=�XA���=1*]����c�z/��K�g irw�;��|jw;�C��T��z$VHB(��+�biƴ�_����vl���A��أůM�m]F�A�G���"�:�g��:�����xr�6(X�K
v��� *��`!"�pDu��TE�1^,���p��0�G�t-\$��A���f��CFXt���p������]e��E6��G�#����/Ԧ"��s�P�^�:$'~� ���b`�:)��7	���"�j"�`b)��u�L��1�zd�%��#<�e#Su?K����n0|��.�6}�����~w�fԚ�k$�^m��F&�>1��lOʴ��O����=.�V��ރU=�#�M��NY�!�0"��D�B��;!󸬔jA�s���P;T+����|���g?cƈ]��@nT�(���f��<��d����H��A��F�FȆ��S�Ǧc�4ޅ���'�H���0�0S0-��z�=����?�S��_��Ѱ]Q��=���>�	>b�N��%v�Sj���\2/`�h��`#�F��Zs��0w]?�nu��V�9�?��V�<Rޘ��lD"�/N�~$� �2����j���J�ϊ�JPB��W}v��7x.;i�j�Q��<@S���scT�a�'�Q{f��8֪	=�۴6�yםe�j">���]�Їx�B�i��ε���厛n�i�\\Z.W���e1���%�	�����*�k>v����t��������w������+���O6�v�i�seF�	���l�(�/�mr�wv�	,�"�mY�'T�ar��XAr���4>��&̓f~���Y>���Gσ�x�]c�c�g���{��}��o�����֭�d^����� �~u��Ul?	����#b�Ch}Z�%�����
��)�a���������
W/ǠePv�Q�c��=ZHY��g�zQT�o���`��!!�a�٘�*\S�pSC��#ZN�-��i�/f@~y"� V�(Wr3Sn�sk�Ff���~��s�30 ���9կ[��«bf2��{�1�1!�U��Y�M��m��b���A[%��~�p�e�9�pBٲ9�P��!D�AQe�]��KE�R8?��2��"3!p3.� �B�Y�S�M���4Q�ÌX�1 aͬ��B����r!V]?��Q��R��z�Ȯ�B��Ex����,.y�ZPyU���]96�D��0$��o� `�r�`��A#����NY�% ���� ���q��N���`�y�8 5]3~����`e!�yIC���V�]��KU����>Q޲Q$�E�����E��C�Ir��W�Y�]M sZڝe8\�������k��I-�󽸿��u�M��Zus�A�6Kj�(Λz�dar�Hp���\K���������;�eo�<j~iMp��3��6����q�Yֹ������i��u��Rx�`a�5��gրSN9�<��/�w��U\�c=��m[��%dr�W?j��������v�˹��;�,�.mH!��zV>RRPv���=�ts9r��r��e׶���պ{�{�FĊ��,K�Ԭ���=hfp����c�h����ޣ'��7�L�U��Y=�3��Csʍ�����*Ay3�Lx���G�,D�KӐ{5�cѤy֤1֣��$���ޜ����={����Ϫ_��w )~�f�,I�65~��'m�z>�l�_8��f&����>��"��]u��\/z�S,�7ҷߎ�	��B�O#͟W�$o�z���C�ª�	B93�;�,%�Wj+%ج��>�� ��-��"*p�,�"3SA����uN�6Rj{*+�ع��_�����2���Xpt�R-�i���f��1��f�,��z�����[,�D�X�����YaW��1I���Bx����$��}��� �FQ�@�o�����^�牭@ŉu����|�
�=����BM�v��lw�r!�}��P�`" ��11�6�Du�1BN��� T����'�e��$�~YЭ��^s�ϕ�GqU��2�`!Gƿ�E�P��M���.�9�׀ň���;Ŀّ�&'�����R�D���ۣb�0�g���/���̂�-R$��c��]��H1q>\;ˢ����e?A	2+�r������FC (uX�^����0@�1���C���&56��ʟD���\k�v�k�7B1�	�l����&�~��Sl�\�lB�>}�k�Pju!�Ʃ����P����5`�{���}�K�Sܢl|�'�և$������։�p�`���7�0�r��R��ti�_��ؠy���� j����G�
0��}���O)+=v@i��ե���NI����σ "���=��rm*_�2cM_H��d����K�W���Q�|����="�}w�"#�X`����y�⒋ڛ�g&2�r��֞��&1�M]��M�+�^��ѓ�4{��=8�wL ͏3��pe�9��p�)������G�L��#[��FS5��_/�����f桞�qM�s���J����qۭ�/���(���g��u�f���/����a��/�C��t3���|�&��\��F��ޚc���F��{�`�Y�u�A�6еt�YQ�����:�墎@TWg!.\52f$�`���.}����(a��u�)\��+n\/,�s�Y	�'��s*H#) P���.��[jw0���B?אav�XO��'g�K�8��4B/���}�'���X`�ѽ �F�3�E�.�<D�D�9�cT�m�FF��-bp!C�^(\�c�Y?��Tʂ�:.h�n֒�~�J=����J
��!�r����.���X3WN��3��1�;�bX1Xb��Y6�G��5����D�״��%1n* n.j�9�Jk���LW5��/��a|q��( Ee}��c�x�`7"�Hԧ��*��ME����p���ۈ�ͱC7������y�Դ�{��(ߒ�X5�O�p#s�n�6y��K�K�r�{�m�λȜ5����j;��b��n#���4�bt�����I-Tc!�!';�s�g�kTc�yl����U�]�I������ Hce��ƀ��������r��m�hǈX��{:'�"Ƙ��X#��n $�6z�	��� ���?��'	�<�"v�g��-w�&��z
��C[����+&Y� ֨\����9�bgר�R�!ˀ�9��(�P�d�t�4u�@U���_�H���%�*��'��Si���9�3���:��έ���ۮ�٥�V�k��Sv�I���MN���ܵ�u��AaE]��)L� ���.lV}������B����:�c:^�j����푘�q=�Sz�E�D^�0�@�yi���;F����~}w1��=-�|g��.�o� �maG�'=}d��}�5�Q���6�7��ޮ�e6���L��
U�d��UB�̭Z�z��wꁇ�=��	n1�Z��5Ǳ�ڙ�j1bW�}Xa���԰U��={mb��r�E~xv���홁"���퓗�<gb72���� ��z*���"�3N\';�q�lk9�\1��`��$������N>k+�ǎH��������a�N�a'�Ӡe��Ha4���o�v�<��Q�� q�
����oټ��`B�/.���93\O�E�#���)�5�S��`��C�		L���i��2X܇� i	*���Ǚ�TB����@;>cl�MCBԣh�+C�D~�Pr�(�6�1!��=C�����K�6��+C�>8�5�T��f3� ��lP���lq4nf����_�T���p�nC��
���6�Oj��d�0ܩ�q��\�w��$��ݩ��ڎ����01 ��`�]�{x.�������nV�}Οs#�,E�K� �1�q�<E0�� 7�	2��W/����-2�G���B�|_��7'j/�6H�� ��{N�����au3 H����sJ�Jn(x� H����n\w�u�r9N5�X3wn��4}(�n���\)�Ї��J�z����2>]e�r�9�h�z�X-���;��N�/����v�TT\�+�������=�����ԧ����
�Ö���3E����+����7I�<973���;��ؽkjnJ��-sJ͡�unJ����a\hf���gi���&����I����Lͨ/g J9_�r�j����������֏�j�����o�����9a�ZE�k�$�W���6���X|ݯXA����~06[p>�L/$$C�������].@(��=�P�} y@��s�ߴ3�eJ-��ј@�`"@!��,�$�Nh�&wZ���+�ɕ�_c����q��[sd٥R#2J���r��
dAC{���l烵Ц�2���0�m�ŝ]L�o6Վ�F>B����#�}�_�����dOfv�9%E�А
�R40�	Q~ ؎�Y	��b������ט�H9�Ō�W��Ϊ�W�-P�����-��e�M�?I�a� ��0Ҥ�m���x��٭51"Q6%
Fm�ۅ{1��Q�o�k�K_S�=��,��� I�/,�+�{�[_�83'�YƽKF��3�x���#r�!�U�^�~��JȺݮ�*�~�x�T���D���1�0��)!:�������Y@�P��p#��9�Lח�ߐ�j�H��Y����g�* ����w�սH f\��_�9�>s�~E�߭�c%v��;D��{�Q�CT�^������ʫ��G� �'�`���� ���d���@HX���7솎c~����T`�L4��cC����1��殻'�c�����q���zp��6か
�>����q�2��]��M��ǅ���.Q%�J�m
9g�F�C���w�Q��r��ǔ����9��E����g�"
/����ȇ?̌���|���\����5�����u޲m�J���1�u�Mײ���s��A�o�jW\7Qg}+�	ýLAc�U��nrwu�M<἟Y��'������,<4��$��":��S>����fB1:а9� �)�
4��Ր���~Q]]#���q�b�a�Ij����:�~,H����
�1� ���u1��B�;jn}L��2-�r�Ѧ&��E��vO_iV��Z�Ě��TVˈ�|�lA��sfL_Yx]hSL��3�mj�A��Ȁ�9�+�	�O�vU����u���I-XD�E]'j*!vh��D]+��V�}ø�q���(�5,����]�!#�Ga�,�d�&�G�#A���V������t�,��RV�l������ʡ�Ӹ�^ppզz��p[-ފ�!���&Ѓ�i��A-��qR�^�@LYgF��`ȴ�ӏ\5���|� *��%6Z�kN�^�H�[Q��lR��4�}��ic��(T�%*QQN��Ui�=�ZT\��0�  �*���;lZ8�I��
t8t(�]�� �»���C�NX׬Y��
�Rd$%DՏ@�����A�&�W�~&f�E-�UUH�&%����xRbě��41�S$z��ʳ1*���KpB��!'�=�n�~|��������Ăp�ԝ�I)`�S���6�H��:a�HE�KʸØ)���A��u݇Kd�H�; p�x�Rp���\�t\�,���g�t-�U�m��~��z���l�K�賌R$�r��o�И!�Í�����E�1m::�ĭ�`C=;�	�]�vX)7��ğu���+�+�W~��5ɥ@5�t�i�]�$���zr�S��q����&���oH��Q�Q�'�Y+0:��6���|Q��6+}��q�'��=JܸO)%��?�׊��|߫2+������Xq����>sfa�?f=��c�`�����0vQ怄�5ח_w�D"�Ljb�������kMGDJ�Gi�)����M\�n�a�N��:�DD��'�/v�Ӕ�Htu�_���9�\0EW,��n�^�@����Yg��Zv�~k^B���O9�!�VL	�����������3,�2 z��MU�.1�� `<�����ȒL��
�߸�|@�̌��9�c ���E8j������]�ڟ��G>�����C�=h?F��	�� 1_V��>�Q�Z�ЖK{aם�qGya����Z��@�{H����t�߰CZ��2�P�#���Wax��& �5A$�Xq�Ї��1"�����g4Rf���
E�	Ɩݻ�zڭY�GQ(Ww�"���N�dR�#3sɂE(��EF4�I|02�P_����_]`��o�Y��RG8�b���`��U_9c��F�!�$���EuUq���{��%���E��WIW?X�ԉٍˆ�^;�,��byX�5��(:*�7�6D'���(��� �\�Mmh�6q���l\[|ϕ\p��&
���7�G�/���2�\��]��s���I�s��y��#�<�d��*��sr̅��۔;�_�zy�c'O]2%�F	���=��~M9Qn3���A�(��:\����l��������ԍs���wͳ^�Kl�Z׺tyYջ��a]����~�Fk��Vj�[������ڴ�(�G؝���A�a��>o.������:_��`-���O���K�Ԩݸ����{6�6(bL�v(�ho�arp� �D״Kǔ_�{��`d+F��/F%� ��xY �s`$Fw�28:b�F�\2�-b�L���.WH*�3��	�ЧqC�Q82�W�E��^~|'��oY���� �ES��i���}A�햱�z�V*�M��.-�,��p
�-[��]L��1��R���H`��؀\��j�wؘ %��������~ZY�Vn �-b��  /e��D��ukו�����F��U
9'pH��h�uN��܊�:���Y�	�	�3��X�aX�$A�C�RM�5�W+��6��$EH�q�ܮ����'@^�fK���lW�p���� v�G����-P�AtD�\���t	q�4M�lٲ�Y�!��=Dy�`�l�a��7fNqU����(�q��,��������"�4 $bޜ�hY�)�1	�8��B�s��:i���2z>ȭcM.��}�縌��hb���G)�|�]�'�t�57��O����7�G{�8W�����z)VOV�k��Eغu@zq�s�y�Hj^g�!�v�]E���'=ɹ�`u�%�&�'?����}�s3B�^��NP�O#��vn�J�0��y�c�Z��CNi���	�X�Ʋ\�7�>�hi�FU��*/�p����5��s�v�_��aΝ�Z�@th��>�&6isb�F�r6��CG�蔫�˕(�p����C{*�Y������������":���0��� �&�ҹC�Q�0a4�`�{a��`PhVh$���h���g#;������jË� ����b�NI�(�H�^,"Z�v���z��N9�e(�,�L
,��+{��R�
_��\��ػgo���z��"���oVE��N���)2;���4v���i�^�pQ]�u̴��v%��8l	��Z��KeX�1N�j߰n�����fu����`Y��;`����wA땺�F��]:G�y@L�.19�(Wʄ���=���˥�^"�q�r�l��a���%C�>%��6k/8 n����]��'�- 7�d�#�7eIb�)� |���"@��"^E�Q��?�A���?g]F���^1Ǔ}��T��cN�D��<ĺv[yΔ�n��|�_,����A�~�ܮ�����+��a������fƷ�A���̂�+�3^�:EZ \Dοd�� Ap�@��O|�Jhy����^6K���c��?��r��T��ps3��ݬ8�[�·���ߩuJ��<�/�^F�e�E�
ox����k�i����v��/��G�N�� I&��s&�I�'�w�K���s��O��f�*�F;H~�3˜��۽|��_��_����s~ٺm����g�ē�v�aa�z��`� (h�8n��-c�$�6�.�d��{+Uje�uڨ(7�zs٣5g��b,��y-�94�[�}�=I�Dz�a) OWeOO�<H�����vP+n;�oFa�d\_�D	�3�6���G��Y����=����M%�I!,��tdT��C���x%�t(����cTS�T�ֺ�蛵p�x� B�(M~xP����~Ƞ
���W�\CcZ�����@a D%r�m!+@P�&�KK�dN�׾����x��y��>�h�O~��(�'pСE�Ą�s\��;W��6�$�]Q\F�@���>�	��E?�x�"�F�W@�ý�����]P6m�Tr�C�7ܨv�6��я~�|�ӟu���64(�@��e�=���Q0SQ#A�B�x&��q%��J��+����YgA�$���הo�;����.�[�6+Ae��D��Bb�l,��a�vb�I�X��:ܰ�Ox�C�p���y��(/��x�.pّ����q��j��s��\y�{�+Q�v�t�%��\(cya�+jӹ"��K��(��Yើb.� q>�э���i��_��r�"������|�;˷��-�܇�)ǞR�:묪�R&��t!��Q��p�|��B=1sF�N�ӣ�>��$#�n���}��o�+����=���ɟ�s�{t��W�^>��U���o��\n��k��`^Υ�a>�� �d�8ֆ��¨�������o*�{��̚|�0� ��Y�����5O���@��	�
�D�_\Չ��P�y��׈�c��|�����|��Y.���b}>�����_(^|I�� !�s�4>�@�mĦDz)�>K5��EF�P����ފħk��c��i�ֺp��7I4���Yܵ���E	��*�=�vz>�~F�'�>�OaZ#�W�A)�G ����r=��dL������&�{��w}rC��̪/�ǡ�~�z���OF,���G-d�dy�YXT�25��(�A������Ac?�Y�0��z`��<W��֪��L� ���x�a��%cW��(����;��ۋ��c��M��}�-�Eь��f����ɚf�3�(\ﱳ���>�Ϟ�+�RViW7������{G�¬�N�?t3vi�v��L��Mh��*���q�л`lm���Q��;E��� ���/��\tمe�c�O�'=�g�㽫����)�������J"<9Jg�� h��s���>����?�:�s���} ���W�,檩���b����~����o.��r�2�����>�<�ϔ� �����W�0�E��Sb�N���8�7�Xd�V���y��p�J�N$�E]T���>*���c��6������� P����>��t�D��p�Ŝ
=�ua�IP���h`�4�� N�[�9��L����*���»��.�3�:���MZ.���2:3R��x�����=��h&�mDv!��#`�yp�3�׬��_���9R�q3Sl�c���-oy�ٯo����o,�|�9���//_��r±�;�h�X
'� �]�Y��dGV�ŸD2�2_`��|>V�X�/���z	�/��²{��r�
�����q��%%�
�;�|���%��N�Y���$"8+@��H�2�M�ܴ=���sIʉ�E������|�_q:4i�T��y��}��5��	6#]����o`����:n��W�Ĉ���S�y��̒��:a�fs�D�%~�siwf�(��2��U�N8�2�,�o�Ԧ�U� ��@�d1���Zs�Y�>ǂ���)�Et��E}F���S\.D+�?-���$�3X2���Wh)j��y��|��j`4'Iag���G$Z_)��|�B�ךw��|�h�FW�ő:�^ #�� 0�����X���v!�۵��%$=u>��0Z�����1T�޶m�w��׭+�>�Q��o}���W#ˮ�Ӟ���{/�]-����P�~ja������5Qf����sF-jb!��q챻5���\�4��З���r嵗����m�*�-�)$�?�6�+V��� �4Bڳ�C�V#�n�
T�'��t��>��{��q��»\yQ���/;���3�(_��ʍ��X��������/��8U���W*��܏����-Q�Q��@�evC?�n�4������������Շ���T��'>�	�ÊR�lذa^��C�n���`���p��7ㅻmF9��ah~��'�\F�b�)�p��������90t�Vm*/|������Z�K*��� �3�����A��5L�X�t�)¨2�¯v���tDy�K^b��[�EW|�lZst������聲G./X=
�f�-Ν0�"�_ͣ�  ���o�Cߥ��.�Z��t��@�s��g�ּ9�s������%D����p�&�.GRD��s �֯��Nm��3���'������ek��#��-�� 
n�g�E��O�W&���t����]2㙿�Lύ�r�1q#�U�h��-��pR��w)�{@c�};���)��<�X�?e=m���|=�w^P���O+���i\�����y�Ѧ)8�[�<=l$t�ZFHr� w��+��?N=��s���(1V�>�y�"2��Bñ ��
���F��7"ن\�,�$���h8j���H4~�0�hm��ūߏ>�L)�\}��XY�fU9�Me�Ļ���j�Y?�0s�=�Q����+_i0�[��L��򗿬<뙿&�i\�k3jwIƛ�<`,-���87�KU�k�:dkn&����ҭ�Q�-n�׾���6�ַ��r�uז��#W���!��{v��zY��%�J���+V�Qw��zP���u�+��h�P�
�K�V��w�m9�r���_*/}�KZ~�U׸H)������@,3̈́0<j�����D�!M`�;}��n���a��o������ovx9���J�.���lF�x$ӕzG	��Ꚑ�(�T��yE���fH�� ��s�u@J�G��g�g��g?�.J)�v�Z�9	q:�=?�*�k��e������a�O��3��m��~���屏;_���o��mxO;����W��\�2���n�A0@�`���"{�y#���?la�Sxm�����YC�t�a����'�׽�u������g YƈW���:Q�=Ϡ#�"��8�"�^��툣�>�y�s�� `���������|�|����&[��N���Qr,����!�223b���*#�m����f�����кW'c���x¬c#}���B��2e�?��1��~��Տ�����-��vq��"��](��FVYm�4S�70B-�h����,S&i6�c1X6.Zx�������XA�7X�0;)M
ތ�v�z@CC�����1�����)wL�4��ra�A���P���C��gA�-`aA�!�<�O���'��c�._����������� �T#ڭ�u��]U���ᢘ��Jų�+�����׾�<�)O)��r�v���EB�5`�ڤ���Vi�F�f�$p�!�J�D������O�)�B�۶�Gi7��?z��Q_}�U���?J;�9plV��i�ltL�L�4���թ���e' 2#��L?�+ƵO;ߓN<Q��A����<�)�U�z�uS��}B{Ө���ŬScU]f��b8�_�=�[�7ƕW����;��y�'&���7�����L���N)�5\�>�e���Q����f���
� �t4#�~㪠>bQ#��`��@�r�<��/O����k��N�㖲jժ`��W��2�!�1��Kw%�]�js��H����I�.F�?�ؾ�i���)�́���e���H����<|�1�k�U��������g��J�� �{�_������8��V���W�O��dܸЮ�$5Kk��_�j�]��F���
Q�\���$mUd܀�9�5֮�E��k��*t<v�Ƌ�y���eG� ���Wq��|�@Q�"�D�j��$�ޠT�5����r�r6FN��} �b-��Ԉk���v���K�{Q٪����m$�Zy�z�t���Kz��c��]�'����j���XA���bLv�ս��,-RH�Z "��������@��?�i7��S�4o�ݔ
0`sXib��ѥEN�,�{�;˙g�!�+�\��;�nw.
�N)�N���FgU��]��c���n�ŋP�G?���m��#�X|qP�#�8�l�r�Ԛ�Hݡ�~"�������
����V��b5%��
N�>L��E�P�nz���v�a��u���E1 �}ܞ��%�a<#<�b�V@Ye��wF��C�uP�����c�H�~�`a=�łq�|-aX�X\cA�i��`�^X�4���䈢���>�*���o|î�
��B�:�0��`gޝꢛ��<4ڜ���� ��U�v��ۑ���`<��J(H߂ȗ~�I�1����ZD�NnT��k�(s3�3�,�w}�P�y��n��R�Esf���	�a>r�5�\:r��r�^f!2lz����|����9*��>+ǜ���߇������8�h�F�q��\�Թ�ݵ��b�����}���Y����D�)W���с���h�����W�!� (j&R�-`j�6�ʚԓ��H?��<�7)��ǟ����6ou�V���+��Y��kV�&�U,�˒�J��{D��{�z��?�.ߓ�Ɍ���08��j? K���� %���N~�Q�]����_���1ю>��ث���k7�#֮.�ܹ����nk�.N�hmU$�zp<Z[D7.��=J^� ��ڔ�+��C�Wc��;����+#�E��s���hG�����������;v��Uu��ԏ�J�to��7�w+�GG9��ːč�e�B�^'�d��9Y�O���sb���[&������8�@p��p�R4h������O�t5mc�Hُu#s2e( .��`�G���\SEZD�#��T훝��yPٽcgy���Q���z'r��&����Z�T\J�p�e���˖�{��	��;��py5�2d2B3��
�t����?B������nAeܽ�?.P��U�7�7�M9��f�ʈՙ�������O�!�/��@`|0�����.-��a����~��}U�!��V�5�& C�SW�n9������#<\��8�0@�>a�M�)�F��0C�b7���b��&a����5T��7��+��m���r�n�D��Y@;�̾�� ��9�����x�)������-�@�|���U>�W����;�<�ɟf��>�r�񱰙�lxl ��s���^��Gc��Lf�IkwԞ=J%���E/�}��� ��HGs��7������Lb���6Z+��D�r>e�p�M��Q	�a]���0�$���d�fܡR-Ѕ~��%n엾���Q�>�����.���g�>lg4@�j!���R"g�ϥ����9X{���r�D�9�\��&@�`��q__�L���R6o�Vz$�n����C��X�^v
��:"ti�W["/$���L�����WJ����7�������τȫ/	 [|���":��FX"��=D�h�70�.�0
���߬v~$�?Oc��c��,���F��<�.�C:{Xv���O+�=�Vt/^����N���q�-�v-�hH��ޮ������qS��KY]��/eFm�Q�UsRHD��7e΀[���*��J�`)ιC��n)�ַ�?��?�����w}@: ���N@��?R�"��DEA��\@L�hY�]��N���������WJ�i��3%L��׾�E�.���f�5Y�^%�C\:�H(J�ȅC����WA�{�\1���
 �O �����ay@��G�������Z.a���o�^���~��ڟ��g���R�����t�2*������
1O`G ���W�A]�DY_�#0�j����|�ϕ݃��	G�P~�E/*��0�[F�+_���P�@����b��`���	E�����NJ�k�r��:@����P�åyC�D�Q��8�fI�������S��d���_�z�K^�1�-��w�y������6l�j�v�b���B�|,A�1.O@9�R��Pz�Y�?�hū���T����|�3�g���7����;nuH�Źz�)�k���'��a�=�@��	 ��`��S��C�����o���t���e/~i�9�������hJ\�_�җ�7�PN�p�F���u�^c��Z!��Ө ~�� Ak7�9�ŝ�Åf��n�Hv�M�^0^��V�C�X�}�k�y�=߮�W����VQʀo�������E?�ݙ���P3�5�������])�s[������������������4S�G�K׈��\��q}�8�7�ֲ�@t�۾��p���ʋW���r�� �6��ԓJ<׳0�*
�s��y�a%����A�a���Gs��)�Pw~<�a�Q�;��7]S��
�x��ӭ�,w���N�:dG� �f�%t�(e�%�=u�x�_��'�jG�����;.��k	���NHfbbT�e�s�q��c6���S�i�>�B���(_a���
��� )UҴ>1@�U�pǎ��L�_�������?Ӯ�k��/UD�[�t�)'�e����˺Z�.�S+�+����r��LJ5�U�b`���Nѡ�h$F���?p�~�#~�C�+^���'<�|Y����u�/w��p��?$*����EB��q��&��RV/�h`�X�c(\`�p� ����ժ�m۹�,ʳ��[��������c ���߉���w����o�v���m�������˺�X����<?��0v1�j�ժ�Q��믻���#�ź��g�f�%E��^�Gv;|�;߱��Z%�2a	���Q|�+��`�\��/ ڬ��ss2�v�B�d �Ec1VKpt�ڧ� D����g���e��!	䟾�O�^\rɥ��\v��N���I�� �� �w R�ƜhBv�/Q.& �7$�������a�TDխ���?�1��/{�4Q�ʕW\��I��?x��������m ֗a�()ӯ�~�-��<rn1vu������jT# 
��l������C�:[����D>��϶�mo{��Z�	�spۭ���֊�"8FS�gk7$�`	��L ��{�3�j[�k��S㣠��0D�����E���V��;R��8��.�`<��qJ�Ԃ�0K��$�&7}r睛='tփ4Ǘ��%���`m984(09��P�s�r�qh�hC�9�rg�ah���Iz�� {�uM j��m�����+��Gʵ��Y2�kc7�����9�&)3�>/���� �0�O_�p�F�����̀
�A�N�{�[�M3��3���f排��ˢ�?�E�[o�N=�+��`, �U�:�zV���as$�X�~eq�$z�ݼ�B�)�`#4W0\vQ�����s�G<��7~�Y�x�p�1��/����o}K��eҥ��3ɦ�s�b8�X��.�;Ys�y�h3�E�$��]G�E��uQ2���4�v"��:�(�-g?��J�xC9��W)r��22�wlw$���v�T�G�Kn�X�3��� �G�?F� #���1�ʓ�~�~�������v��;���_��[7��~���ƀ��8��D�s	c���ꀬ�vs�(�:�g�V1WC|+ )��N�K_��W����S� �
:���+^�
�w.tDz!����[�x�� �s����LMQP���2YM\9�gK�B惎�Cٲq�!C����w(_�-�%e�"˙�5� �ח+T��5��mZI:�bOm(�C�
�+�D\7�'�%�C5x�~����׼�5~���9���?��#���W�D�p��)/C� �n��<sV?�D�֕�B�˔�q�>�Q����|�����v�;�=�O*����f��Fy�sQdX��E�ab�5��8pa�0.N�Ȅ�� :�s��ҋMS��ՙ�?��d��="�8�5\�h�.��b��>�_zu�s���p����'�p�7i��q�#��{��u� I-1D�T�]R��|v]�7ma�P��2~��H�:�(9�B�am:�]��֬��CC�p_��MS�O	������X���#-�~�z`�`�'b�	C��@�n,|�Z�겘��=QP��Yh��E}���>���6 zX�� PiZ�C���[�a�tZ��:�,�-�d�v4���%�~��*�b���r+����;/v���p[�m���ؐ#���-�'#�J߽��?A��s��\aoV�X�Mb���V6�2Z�ΪR���QIQ�"l Z�%���%���H$`(���P���<S9_��^֠�UJ������S�?($�O������T�q���J�8\`�aa�"�md�cTH�3�9��c40��-���1�?F"�#�R�s�dzYg�]�E�`�ey�pyE"N���yFL�<�P$^Υ"�ӝ��,O��':̾����w��{���<䡎�!�w�����F��|]���{�O�hv�2 ͻ�������$v��{/p"D��q޼es�V׀�qM��RGMP���q	0+��n�T�	�3
���#a��*Ր�:m �v�΢'s�f��݊��y_�D� .G5
ppm4-� ����i��2z��@��#�=n9W�B�G? P̧��x�y�JuL�����Qp����  05����M5�=fVt��N�1gYWߒ��.^��h�����p�gh�R�}���v�#̝���Ĺ�`�@0��s�B9B�؀*����A>�� �?&�C��\����&�Eg��LXƚ�:��!3��z���J⇵��g�C��(�k��:`z��el�D�r��U�����L�?6>�4>�'i����� �Fz'*�|��cQbMB)���	�7�!��Kc���H$b�db�p�r��+�6��qhfp%i�_ w�>�}����U�<�%�t���}��^q�ŕ��N
V�.,��;L�+Wh'�t�,����a�.M̙!��~z�����B�'����
<Xl�F��� ��)\7z9"E����T��ڽ��?b�M��~� B�ǔ��,��2��L���𰢣��.Eōi�I��ԗ0��O�u�K�=�x�8�
���x-W�V�c�b��	Y�=y�&�5c���w���v8X�{L�Hm�o�!���fW��M
�����HװOb���G�h��"�vi�	��V-'L$�#��#��0��*�4S˄��[���[2��燎�x������cj����fn����Q͉ A0 v"�2/�(�y�Ffm�45� X�է37�J}�X�)����> ߵ�|�	��@0N�MhL��qf��� ���2�	�v%$�2���A�ܙ���I[̇ ̐�B�j�ؿß5&��YȖ1��M���戂��q�����Jt@A�ٝ[��e�Ll�S'�7�&����1?�w��)�������и�g��>f�����ɕ~�p�r0Q�囪�G��cUw d��2eCs��Z�t��&���W��*�1X.��rNٛ6i� �������p٫��e�V�Į�r� �6"�#��g��R��ĸtO[�����5=�C��
pc2-�_6.������":�!����l�{r-���n�����t��9���8ޝ	����6�4&^�����xSx)���:�@�����&J���N�hOSC/2��|�k�co�%�Gdg�5��%�h��h10~�e�r�h�X�K
|�N&PC�@!�����H�����Ȅ�P�\�rx�������Y���)��\@m`��,��GwM��tT�ay�U�v�;֕W�F��y�m "x��6ch�RcJڶrx���.�.��"Z��1rfO��[ ��jL0�y&���+�`9��<�h7�@k�d��p{f��.��%䱯�1!}C�p\;�� pFj�0���,�4m�	W��M �;t
�"��j�	�]վ�G;"l;��z"Tֹ9�c;��*B�)����B_G�� �����\�9�9���!�%�W��F>ª�O<f�N{0���5a��&�y\tU��閲[G���?]{�\w	\q����dv��y\�y�e#�'�lK�=m���pvm@n�mh�iQH�YO�8��8+���K��pң��=�� ���l �k2��� ϊ��EYK�ch��M/0��s:r!��˼�T�*���>�A�%7�W��߇�����	�צyE-<�w�ޝ.��W�<�o:�E�Ş�_ ��ۍ�0w��˖�S��ψ�Գ�v)#�sv��4+y�]G._�~獷s��7�g'gf�Q�l�h�li�5#?Z�F��]��g[5�5�x&[�u��\-ad3u<���g���yr_��p��?T,���C���rO��"
�(jZY�t���{���\<Q�)�Bw{A�h1�7���Xd��#y���"H�� )�$l��`k�Ң�-���(�97)����eK˥��3�h���)�V(.F;��~h��P'���w�͂�b����:x�E�0"T�Fl�:t �6�&�ȶ���܄�g��a�C�̮��t��໬IDw�ؙC�[/T�C�&�7��nt��i�W�/ Z��Um��0�I'��y�[�Cl.��q�c�${=ae�_T-�� ��(q��e %��� ����=�F80,�h�ˋ��)-�h� 9�֌/@��XK��h|�0n62�r)�?�I)���+C�q[9^R��Y}�k�e#����g��^�gou��Y��*(��\JÜ:�t�eC��1��f@�4�W� 
���a���eܒ�3˨�H��kFPp�8��P�;�S!���P�,�+�}�o�4g`)���r���*1^ ����n���> @,х��}B[�,�cP��S�M"X�x�B�,}��>�˽ N�4`��u��^�vݼ����pO�7��iS�u�:�tS�
�x�mr��Nڻw�>��8����.�Z�����((A��I� {�;���_sF�kk׭)�y�RJ����'�)4�w�ջ�v�l���)��H�/^���/�Wm,���������W/Q4ٙ�iG�����jmj3��F3�E!�M�OM+��&Mk�4��0ݦ����M�?�z��kVϵbP\WrN}1-Q��9/�ֽ�+JoLc�8BJ���1)VSt�dOg���s�nk����6���������֎�aٝ���W�����-�ց�0e?�_]Ap�o�7����jL?�a�̏b��.�{��p�4^��:��O��4L��G�I����r�5g�bâ�]����
�;k/�=AB3��D.� 5Me��:ch��G*{�J/��c3���/ᦩ�A(j-fֳ�EHu��s��JhBT�=�:��a�n!i�v@ l�ݺ6:tF<��4�S	��u섄ڴ�s�7���w�n�
�! �k��tR���C�1t�c�}`Z���0 /���ON"�V�MW����`�~Kf$��=Ɉ��2� �4P�G�n�EZ|���?���I�.������� \��С0�Y�
&�����&�g �� �2;�a� ?�f�1���8�9���{�o��H�c����0y�q]��\?���id��9y�K'(���_���wf�n�y�d<�ېJb���$���;��,�#X�(&J�16 �F捿�N�Y�-昣/+S���c?��`J=H����b����s��/#�`WiO�DĄ���ql�~��LJ�"c�gn��"A"�G>�>-���V���WX�GAT������5�K`����u(���O^��*S��=��d(}�CU�1P�ʭ�3�� ��b���P���`� lK+�:��&�,���6yy$���w�q{�����ܵ+�ꤞ���|\�Be7f[�ȸtQZ����M���ilxpE�����VLu4��j�X�1���* �ǈ�l��J�6�Ƥ�sOb4db� ?n��-�ss�L���M�qff5�4��f���J�ߥr8����Q<��QC�y��sV��Y�z�����:����,���_Ѧ5��.��W,����]G�{0 ����=�@�������{ � A�OCC{x/���Z�F:=AP��Hbw�k>Z���i��`Ե��������\��oc3k�0��ᅒ��f��j>FCoe���������j(r���	uȽ�{�u"̹2,�wkDD��M��-j�S�t�^$�� *M��w�y�܇������V�<Dh-����O�c.�c$d�_]������^��9U0�)�M�D�Ic`�*����>��4���ۇ{G(�
ظ>�k��� F-`���HX�­�a�9ҝ���J_3��،��γ~z����Nc�ȅ�����`�5�t�L�}���_D����e��ڬ =@¿����2]p��o�D��*�q�@��xc	��c�}g��=i�pAu/ѹdx�+�����!A!mu~J>�0-h��C�S(�:�<��X��p_�F(�\R�N�`6-wF�q݅CF��<�;O�p���>u-�偙��������ј���`�_R!�Q��J�:L�~�`+��Ql�ꜭZ��T֫�TO4�p�_�V���\�A:K	�8�?ֹG�uH7$׹/�\h����n��Zbb� cb���K��2Q*�GJ||�[�)w*�ę���.��g�Z��:N��	����_9�Z �=��|��,�l�]��}@��srtBd_GG�ܧr����=g&pz�)�<� �ʺ��\ϼ�� ���<f��͐]����:�O,Qn)\O@�ǽ�,�kF���}���Z'��Z��o�c�_|�>��"�O�t�aW�vl��4�@w�%,��2D���7�	�hI.:<�Q��� f���صZ�"�Ц(���ף�Ŝ�p�B|����v���w�e��N������f�� ���&��!��̑��7�*�S�T���]ka�VD�z��n�i}֦v���umNXp�Gϱ�nA2O����Q&]���O��1��NLnTF����9G�ՑY�޸���������̦���ۋ�o[f�&$�����ٴ��R��t(:שF�sY�+0�F�Q@Zۤ��H����(�a�W;Ӎ�@1~2:.k"a8.�0�a�X�C�5���}���Na�r���ѷ}r��W\FP%+n�x�[�c�v�v�[)��[��W�^�q��>%�Fk\�z�]D��wiI�Ř#h���� ��M}�J����eZ�K6,����$Kb�
@��u�<ȿ���>���쇜Şy�F��ĭ��x8"K��ui�#�`	`�`3l�
է}z���y�h� �0�c�Hj(�����|�䠿0��7' ��좋�y��Q2�ߑ. "��6�{!���߸Ϙ��p�X���oJ��=�}�Q��R�8~D�d �1F�J�h���N����$�}�ވX�r��(��M���/[�s)G������۷��ؽ�ܶy�A�I����>�6$���թ ����x����H��%K��?��mV�f�VN����Jsrv�E:������z~,�ieIP�X+d����1��ߛ3MaJ4k]l�&bnvttnrj�����Uϑ���Y=6�*������Kc�{��&�=�[�>:x��\�c˶m+{z���t�MԿ����U�����[?��( ��4��!�9����[�Z�o�O�n�6PD��D[���=� ���%?�<���`��o"%=zv�l���ʲ �PH0�諕;�a>�lP������Z�0���h�csy1�
����P�ι��*��Y��ܷ�'�|�$j�a`6�^uY(�b��ϭ� 䗐n]�s��`�O�.�R��>�5����hR��<����f̽A�� ��,�����i�k���s��n�-s�F�)B�c�4�����ǘ3�{��¬��^F��,������r�l��s}@�@���c�(����}�ͬ<�ݕz�������+0)���x�h>Uu�3!�q?�d:���s�8X<�\�+�M() %��v�c���܋��ȿ -�Bg�*��U���*�_}nh�ѕɪ&0H`k�	]�@��Ww��F�4�ݷ#|46_k���d��?�\g<����#p�����ɰP����F\�&*�|U�7@R �n\���c���"���X�ڗ��.�-���2N0�Y0��ʹ�d���pUF�
��u�h?נ,�Sq�ޘ��^vi9�ӜHQ\ߛ��|X �(������;����w�( ��v��Qe�7��nO�t|G�ɛ4�lǝx�˭t)�]�=|�yڨj~(4��Mt<��r�)RlF�.�ы����][6�ݷ�i��hZϵĵL陚��gRB�I����x�֚&�f�:�U�\i3ۦ��o1Q��L��w�A'W	��ix���M�3y�	��
]��3׻l��1%����t� ���Z�w�0�\Gw����n~럽u����*o߱����bݿ�"��u���9�hT7Չ��4U�?/y����7'JF�З����G�"��qg�A>��ߔUD��9�R�")p��
QY��â�wn���+�b�@�*i����L1n����ؑ�B"�v��O���R��0FDaq�v-�?�3,��6x���&��:��BR�Ӂn� 7�lZ�5�t��2PD'�7ax�c�0l, ,89g`����ݧv���0�ܻ��x����ݬ�.=��#!C��r�z̓=c� �H�<����x��y�.��Y�p|� r���r����l�f�[��O���ܗtvi/wV�����iCAfv��ĥ�{��F���p���	8����ȅ+��0����%'CJ�)ݶG���> �ǐ���{]d͚��א'���s��8�Ϯ���ܰ[T�(�P�J��2v�T ��V+���Q��Ԇb|�tP�`z4�Z�#�"
,���5N .�?� �!�$�B�n��Z�Zc��U]P�q�]����'+U�o�����5����Y���Pb��zZ:/����02�>��0"�sa��͑q�0�r��s^!�1�g8�&�m�Z[z� Q��"SN�A3b�FT��4�t� ���޲��b^��
��OP߂kRm��r�-�O��r�
2���)O|�T��(�ץ�1�N���a�t\�Sd�g3�9��}�� v��Ng��3�Ƌ~#�&%zp��k��HC4���)J�g`�&��ظ�5V�]UZԗ�
�z�����Ǟ���֦z��I^ׂ�k����n4��̤��M�O���7�� 6�Zg`�b�0i�]����"jKԢ9�K�jh�ĵ
�=��U��.�@�9m<��z�dwWOc��=���7~t,���G�z�v)L��b�5�'����_�ii���f5Ɖ���t9���ֽ /��7�n4��j��XDxNà����"AZ��u´�A��Ov�z�j-�wo/k���#N9��ɸw("l�έ�̳�p��	r������/�4��W�B߮��42Ƹ�X�i���%J$*�EtF	;�ZK���bZH��ު�\�����l���)|'��}���]��Z�`�� �'��!1Ȅ���h@�o1��++GB�9��^Չ�G0���`mt���ݸ
���E���M�� ��I�"�}�]$����lۈ�act̰�H���U#ѯ����U�(�}?��psoD-!���*A����0Έa�*
�93�zU���.%~rX��^E��ݍ�S�9r��xh����hK����׸bq��D�@����ɸ��$���#I�(pe������d�k%¬��Т�x��,٘� O�h-��.N{��\/0Uu�^&�A ��{l�yf�"�ML�*�@�R
��d���2�#�>� � N�����'��eH�,1v����>E��H@=��`L6�jd���'���$8`*���f2{6ü����L�r1�)���;�|GlƜ��?���7d����?R#�a#Z�y��P��=�y�#��ی~e��T��'����(��L�Ђv�$�=z6'��0?�>���
�ɺթ�3l�p��z�i�"�]wp�U�+��X���ʯ��T�F'٧m71*�t�y�
�t��;�)�b�5��ɤL%�-�z4���MO̖�#x͊��҆���2.W5��1��R韶�ܫ9��)�}�lKSk�p|��X��yP�C�y��e�k��E� ;�#�]�"3c�f����\@�H��c�RT�q��%
`¡l�}mN.��Np�hK���p	̃�
�,�s3�Y�q'��w�_���r�QG����o�cV��=;({�]��ǚof����R��L�����-	��A0�]�$( �T�I����j�s��|�u�T�/"giFt�=TmJ�S0g��c�(']�#��)��ΞϪ�%Ȍ��ܩZBv� N%��� ��YÂ�'�JF����p!dY���@�����[�0#�����$���ƫ0��~l�z��7>F�U�9c-`kw��.�pO��=�q}*J;��q�n0�	��[��t�����C�Wא��4qs�#�O,g�q��!��Pv�T�W��e�ve��Q��8o���U��\h�>� �����qF"B������,p=3��t���6�Y��2����e�gTs!E��'��GG���-�0_�Լf�ý~d���b� �r.x6�{0��#ڐ��|F��vPi ـT�84@0��>�jm�Keu�l2Y�!b>��m�r�hS`���r��~�;���~�Źs�nϣtq�e�Rϻ�
Q�B�X\�f�6;�R.�f3Y�}��$Z�V>���(����Y*��y�:�@����pX��W���wP:�f��1��?0<�~��9]�X��d	`;�Y��Ir-�'h�"���f�������R	0�c�3$X�C��X�����53>�?�|kGkK�X|�T�����?�r�n2�]�Ъ��{��;�Wa����>]�G4{�y�W��3��id�Y�M���e��/W��������׾�\�;��}ʲ�\��]*�x��%���K���͡�����,����DF�pz�����0���+�/�S���a+� `r�ȖcYd#��Zb~�|.$A��7�g�`h��qI�u������LFHi�
,�%Z�~ff!�<5=nj^R?AGd'k�*��v�~j.��i�ÛkVh���/ʲ�<Q+������V�j�|W�J�3p�ErJ��{`���|�`�8b�m�d�Ȯ����"���T��s�qB���P������ɪ
������gq[�}Vn ����ӧ�#l
cn���v���2GM
j�KΛ��J�LH��'vT�^�i�t	�� ,��� #���滙x0�gy��MWZ���vr��L��85A@��q���\Y�H�8>��l}�w"�s0Hb��.8�8��Rk�nK�� (��yfGs�,�\�䍸�����g�O���<��#�$�1�(C�������)�>=Od��(�&J�gZ�y�;�s��5�D�� 7�A��h*�"w� ��_d\S�P��=�
 &oD%2Z��C�q�Pр$`�sS'�tR`~�V�̵�?�,/��y,��� #�2[�W#P !���i�����6#C��<Gw3O6�h��(8e��kWHV���A"����MG������m�*���W��R�WE�[��lF��\��F6��:44aT�
�
(33Ca���`f�pD9�����`���� ���,�hKԧ�D�F߷ؽ%��D��M�^#�j�4<'j�u"jTjH��rB�q;M@�A@��:v�+C�3�s7������ �C�
֊vf����
p�4�}C����eU��@w^���Z;R�5����C�Z��6�Uw��V(�HF�:gT��UU~_�~�ڲ_E_��nh�����?���I�@ ,єF۠
�%��V��S���:��#���V@�h�} �`��1��J�@p�}�Ѵ�#�^��>� b[�6�r��E��7��r����ՠ�K�=/�`��0[�@�v��H��2B�ӦM���n�%=�Pw>�Η:$Y�W2I�+���;.Y����Mmwm6mn�h�8S�����LS�?�7�s83�f����p�n�\K�9qe�s��o�UN�fm�V{~nSh;l��7�,�nf�߰�Q����{��O昂~"=>����b@�(�(o��$�JY'���"�6��Svj�6�s�g|Vc<���-��9�_?M=���h�4kQRГivW�F	w��ŧ�:U/�Uא;�\��O3�n��O� ^1ų,E�� ��������W} �%b�.T����
�d\ݠ��ZyE1I�R�d{�6��{e�:��>@�i�\�`D��ˊc��-'��r�ͅ��X�����~r�r����7�u0�|�����"M�2��8��HC��(���1�ac�lE�~����cXls��龎��n5Y'W�;\��PF�OV'ٝ*V�Ҷ-��Ic�ƕ��}\/K$0p�Tƭ�pfi�"�q�Xԉ#ÐEdQoB�e���p��}��j1ͽ��ۧ�7���q��������A\j?��-�N��?�2��[����z߂i�	lٺ�!��Q�@_�`�����(����ka@r?B�����L� �t��|�J1oӵs5�4�J����c0��c��W���-�E�'�g���"1��<���H7����T��̈́�-T�qnBpK�EC�<�.��K$�H�|��L��������:{f�A�uE};�,׊�& eu��>�t�9��>�ktЛ���!!3����;��c���UXh/st떭���.��Uש���Dc�U���ci��޸�C��Q��U�Ba�N0��P�ճ=FrC2�K�?>AnJ�Dy!�4�"TW���_� 聏��@s-z�%'q"L��w2A��n�L���댙���J(�P���w�-��(2���@X�b�r��%"[/MQ��\t35���ErP�-�݊���]gr���AJD��XT���Ż�LU�٢��źJ����k��b��pa��
� �%��п�{���O9CH�O��}h9��$�^�H�D���<�h�������y�Qdqo����ܹ�~ K���-����>0(�b�Ƌs`4�DaT�!X	X/"~0�yO�fg�7��)�e&��nk���xF��
;�yU�S�g����01��+U�;�9�C$`l|����w7i'����_���d|�\W�Z�{�XJR>�;'�$y���¥O
I)�:t�sNs&Y�dW�7�u�J�M��Ƞ��'�K�{K�"�`�s'��\++�3W���$�LSf*N<�$�1Os�-�U7�`�1J]X �V�[�6	��!�h����\��$�*�/n(߯�a %�(5<Q��N�66G���\��g n�("LٍА�π�d2�����ϙ�����=߽V�7c�w9c;��]�x��;KE��>�Liؖ�y� ZbiF�<�g��'6!�&�#�w�{G�Q�p8Һ�N�u�8���Ǖ����T�C��Q�Q�G�K��_���m���Y��7~����6/���� ��W�`U���Ñi8e��F$Z[/L!��>��Ǹ��H���k���n9�-���.JbE��*�t�_ީň�M�Mc eo�n��7lX�Z=k��v�̳� k2q����ga^4Q$3v�ro�#EN2�F?o7���#�3Z �ó1��� �����v�E�Gj�>L�;`���!ȕ��r׎1d׊�)w�!�U!L��5cH�<�����qs��w3o
;e\9�M:��4�
F�,�@�T��x�u��GD]���	��{�J�����v����Y� 4C�3 �v�H/U���Ũ��Q���煱A�f#�Y:JO��e0�#�0RT
\�("MȰ��w,��U5>�1�6�
�� �>�7�U��?�c�'@Me��F&4APjz	�wj�K�2�']�K(j[�g�z}V�t���yM�$��|���&��ۄ��|&�0�Q��qA8��H�G��O] ��AK���=��މ��꺌	��D�K3��]�^��p��k���2',�w [��;6(�+J���L7X�9E������/��9������˳����v��իW��N=���S�R����9�xDy�k_S��ǖ�|��J�y�}µ��)�7�v�o�ʘ����v�^m��sOt`Xd'����k�1UDf�@���4���ch���s_<�M,F�=С0�A�Vr��� bծ��6���ڨf�^�|/ڤ�����!�uxxB��Ouun�7�̪��f�0���#��L��8(wҖ���	ǝ�]3�iІ���0a��2�-��)��i��\w�,�)`�d�C�)h-Ad��Y>��z���Øu��Zh�m�x�MS�$����0;>/�����!�����i�K?蜸N u��a>����
�:)�9��)����U��]��R���dE��;l@�ݡ�Q,0r�J���T�B��( ���g��޽��h�Z�	���Β|0�(?X�HD{a0ƕP�	$ɩ#P�ѡ?x٠j�$`%�L�Csn3B�`#�k�N�b�uRj�m�Ů��r�۩�NiX�e�n#�u'�7� �Kԝ���b�rӯ���Ξ�&���|N�0��F��Y!�͈�=�BN��Y�q�y@#�E�����@����D�U���	]k��mkF�Yg�4�h���r-�1�FD��� <�����NX�`r���W�缀j�)-���A���xv���W�˦�2 �am���^�(���oh�"zrґ��@5��ɒ��Z��<���F4\��lh�x�6n�hWn�n��|�K_�Ɖ$�0��+��ԓ�)�>����_Y�<?�ڐ�ls^�,o�\`M�2.�aD��\���U�(���i櫊�����En{��]�4cc-���D�1<?��Yd�����R�����1�.<��|8��<P���6�+��d4X�����N�x��Ϊ�׈�����P���"-�9�2X, �S�}��E~��g����bM��1�����ڐ\��a��®��r�	� ��횯
���'��Yޫ��H��L�:/�G�5*+D!Lt�v�]t�Q�h�p��06`alc[�\ 
'مԠ�&q!���E8�1��['�S�H�ƥ�<��g+Zg�<k���2XQJ���|?vOx��0f҂�	��ڔ��/D���Y�7��q 9�+�_wݵ��~�.[ج�PqJXv� kv�w�q�˯�_���j�	���X@p��W�Ez� ��H�Sۓ�FF6�]?v%����6pOb��7���<s���ΕA�mH`�����xS�Eh<7A�|ޞ�R����4�rY����zX:�(�B42�1ܼ0B�9�XZ����F��7��/ܓ���<�!ժ�E��z̨ P���l��L�Y�s+]�#W����bc��s�C_g:�����W��o�Vey�9ڬK�|���eZs������n.?���GM��/+�����*�Wܴ�͜�樲��k�E��sĜ[�k�5���J��ҥ~�����H
ݦMذ�	�&kڬ�Yڊ��{�������c=��=ЮtR�l�vyAw���6�G��J�BR|���QߋE6���"���>�ì<�9�*'�t\y럽OƎL��%&��uʀ���g�񛔊��r@I�f���F
V�Z�Ij9�P��[O�sL����?�]�8�~Ȣ9.��@̋�h�q\�
�05���6-�U��1eOypt	�>@��!3�̤�-�U� v&5�����S������@��<� WU�L{�ݴ~�:�ÕLF�D1�3�(��_�$	/���Ds0T�ci�[!H3`�.3�- ���Ťy`�̶	a����D��F��BS�4P���{�SN-�|�#�\@�h)k֮.6�P��\|���i0R"Cv��1H���bu�o�=�	a�JR�t(;�<��<=	�2�<�I0$	R��ioj[�ա���Sp���Q{ӥh�۹�3E[�MLA2T��t�W��"�/�QE���Q�|U�ZD|����4Z7Ui����i��3S]�m�o@1m��7ne\n��ʄ�[�d�\�J���9���r٥�5Ks�ǘ��H �oc��Зըˬ�\�ṁ��5*���Q�zT������E1�w�G>���g��8��1�)�M��ct�ח�|�[�K..��Y#fH�Y����ISVe��)��O!܌}$���T����6:�18��P��
)�/���p������w/������{`=�!d����f��0v�0*r	9��u%��]���}���K������H��4;uv�,N���w�W^U�Ĺ2��2� '"@i�¸~�r�-���-g�ur9pp�CT3�cK.�I'~l�=����^�Hw������cw��L9�`N�/��<#խ�;�f�G�p�TF$�H�q踒�Bࠍ�٥����� 9��ΓU�'��å��"�Ti�w^�I�1X.�!��kV�I `>iu�� ��0 �n"�"����1��.�RF*"�B�E�asn��V�2c4^��K�>������$ߦ�D�;�\�h����s~c̸w�'�a���`���qS ���_��cv��c���'��Rf������~��V~)D����r�" 9�1��ZU�`]�%�p��U���`ب�΋�ѷ��i�Y?��Z�ψ���չ�wy/s��2`	���[8c��H2�G� ��Z]ɶf	�d���cT����,����A���"����wfm+��g����)�Y����3Y�!ږ�,*����r�E���<�bA������o��Z:�`�g��.R��b4+�:��>F�=:sA}Ja҃҉�~���ѩz]/|��*2�h��'�ɹ�����a��5EO(/~��#���򊗿����Yt\��0���q�	'8���n��e��4� �c�=o�?Z����VE�]q���_���e��3i��̡	Z@��i�]<�ǹA�=꿨΋VEi�� �h0P�����GQ�f�%O�B=�z��i��Qĉ�,ɸB֯ۨ��l��=2P�BZ�ĨM��g!����.���N-g��`Q�se�����M.��AIڪ{c�n�/��{�Nh�)�@z~���Re�Ɖ�����:K��J�����#�� g��5"Q/�?����i���Pu?���u��jakR1�cd*����ݫG\Xfd�kE�+�2�	�5ە�vF@�M�t���0I`c<�q��4���[Ɓ� �I��[9����]�i��/\���!P�M�Mԗ68Z�'&IN�NI��8AD���#�kF��r*�@9J�2�|Q��4������;��A��%�|2��.��o֣�"�*��W+)�Iy�����?�� �e��O/k�V�[o�Q��l߱]�n��a|\�Yms�
x�U��O_r_f�H� �&�T�)=�6i��>���vQ�!��v�7�C�D������h����~ m/���$�R��Ƀ�3Vh���x�(wrG�,:#�H�j~��[G||n�#t�y� m�ڥ����� �́%r�ڭ�����oص=�}B�ʂ���p�X��%��Pb���Sm"o�����,`�Pץ�v��{W^q���A������S9=���^ JPKK5v6*���ٯ�,p�c�=�J���\~�����C4�L�{�ψm:��%��I��lV��K4�>��O����-�~��+_��K��?��ҖY����z �{�E�:�@O��LMj�#uv�> �r������J��).~�]��-�+M��Ӫ;���J���맨A�l�Su�f�iղ#YT��`��Q ��t~������0^	x�w��7N��<�ܡ̬��EZ5��e�\&ZԦH��«�ӊVg��,�nW���ejh����r��.[���TX����fCX�����
����~�9;�Q��� ��ݞ^�?�Od�KA�0u2�T���&��	m�� �&�0yp��>MV`g��Q�WB/�vЂ��S�	���D�������I*3袴��w*�$��Mclw'�E�!-�T>GЬw$�kՂ�ZJ]�)�c*Q1�h���D� ����IQS�\�]��Q�t��b:'F�Q�P��eBQ ���մ�$l L�j�\c��/4#�+3C2��G�&�d�. |���
�?&����9Y��0W\�}e��ڎ�����(�E�D�U��#�в�#����^:U�Nî(E��!ͷ�졿i>G��I��0 �Ax�ߙA�5�Y�$=KRO�{��i�8�L}U�̙�a�@�%���!�+�v^�
�8��Ts��f�/��artg\3�c�N�9DS@�1\���� �#'�$\��+!0/g�gKĬp�{�l�W�4m�UD3���1.��
�d��X~(�
��o�"!�� -�N��ϪU�a��y�� C�U/�~]g�F	@Bl&\��`������V�u��w��{\��[�o�<`t睛ݎ��:��x^�6�c�:ʐua�@��?��_�%�ξ�q�3��H��D��K�lN� ����բx�;4��XݹT�\�����ƕ��6�̦��z�c�l�^���fT�Q3.H���OI,
��@������w�>�GP0?�.5� �w��,L�>����Av�i������;�;et,��ı�-c}��WK�x��]i4��0�.|*�3���2g_���D�j-غVc�EDQ�a�=#�['�0Q�
��@��9g�&��ĝZHDYc��
��e�\*�Č�/:���hV�'��r	s׵<������;P�;v�>�G��4_����@���!�M11��1���8z�� ����H.\�m�jf{��]@��Z%����3���,����T$6���r�KƂ�8?Y��sλʜk%�2��c9GQ}�Q�>�kP�_�t��#�BP�BE1�ލk)KJ�^��-yf1j�u����B/��0��#�ÑV���uּ����c���֧H���)��ӟ���ֈ�Uø9Ÿҧ��f���cT�'�&=��;����I�����m����,]�����q _N����:o��,���d�2.A����3�Z�y��:�s�2Wx���#w"k�W����}���p3F��F��mN̯��r91/�C�ںu���o���.fͱe�Mv����۲e��'�VX��FV�S`o�����������g?�ܥc�D��6	���ֈq�Iަ�����P�%��Lu�Z���cr*�h�ԥ�e����srE�j����63+�t�Ĵv�����Xd��Pk���qF2g/TwO�SC�z��a>47P,���`���$٠F@�2��⸅���f��"F�G��Vj'�e�4�ٶm���ڡ�#.~H�v�֓ஒ�b��S]�����K .���.���0z�J���]��������3�3�?����"�pUw��@������am��`42�p�p�D�.#���A*ꅾ!:y�|�fP�=`90��YD���MF`���,_ ���x��j�0��Y��d|:Čp��)��l^��"�a��\fc�Lک1�R?��Ȱ�����j �=�po'���!HrC��EL�v�s �0~0Im*J��o"�\@-M�$h��y�\ߠ�j���*�9��"��<I�b9�H���e�{�(,��'C��鋨���&���1�莸��?���K.�:7ʙ���k�Pi�s�ŭ�*�
`g6*�;�!����X����ߝ���'�4�eɌy<�S�@Jn\|ߺg\�fq4�̗t�s,�9˼�vtY��6�,Eep$��eɜ�Ṡ=K�*���&�&����q�b���B�\���.���D��>�;���������*aϾ�
|X�qnes�g�6�5-)�;UFc >l������[����|�(�77�8.����Y�i��:�1�S��	m�ȵu��t� ��sIY�98t`�R��-�sJ}�[qh�hW��T_�r�,�~jz`=����W�uGIT�o�ㅕ�H��@t"Qk#�� h!,=@ͽi�o0B7s�8ɞ��~�4���Xt��#]8�Ek%�UT�2�(P�΅h��e���d�V�X%�a�,��]���������0%m������o��~�ca��,��Ļ��棖��.=v�D��sgq�dօ�8F"C � aq���F�v���E!�
� �����L���V8"H0��6���C|����rX���xA_3���v�Ez��q{Tm]�� 3�]w��Ԕ4F�9t]F��s��.��,ӌ���-]nvg���b�*�J[S���8���D��D~ M�j�j��0��Li��VsF}�+��_��U��	)q�ے%��A���=�f�-��7�W� �d�B,��X$�\����P�����\c��%7-&�̃G�P�y�7,���ǚ��ZX�
�/� �|�_Ѿ�}@ ��|�&�L&7C~�v��jɒ}���.�#}��hf��v�7��{�$��h�O��	�U��ʹi+`&#iS�"><��}�KPdrF洳,70���r"D6#0�r+:y�ژu����f���y-�gnV��}���v��G>�b%ʖ�p1�g��
1@��=�v��~�ʿ���?�g����I'���c�W*�ǈ
�H��G���H��m��)�i#�Z��%��̜D�곎)"k��U˺��[�p{"/�~*z`=�a�a�;w�O
��:W�.����?�dq���o']f�+�Ʈ�gk�L�^ AZ�"���uk��O��ʄ��@Yrک��*`P�V�ͬ5�@� ��5b�"2�ňE���v�PqF#*��*�E��L���!���K��'��8\��QM���P`���U������M����){vc\U�[tt9��m�C����'�BAi�9Q5( >G���bQo��2#��WWS�aq��ާU��i&fO��ŵ���^p3�c�!hi�+2��t�"C��������$�CB�>�Qu5���6u����\ �&Z�r��n� Av� ���X�W�(0K�c�8���x0hcƵ���K]-���<��
�e��g�;~�x�"1�p=5�E9�p���-C�~��1g%�ձ�K{`ҍD{x�0��6#z���t�.i}"�LI��p\5�\��}�^�>�3�<�,P0\胂ť�N��3����&��\��E]�X t� �rʬ6�" ��Ͽ���|R����Y���Zh�̮DT!��T�	
��ؽ�`�\D�؆ul��?��C��zV5�hF���.�3Z��Ҩ	���[�~��y���Ψ;�*A��q&(� '��Ji��cܿK�{��n�x�*`c�\_�֬пr (��-�3~QI��կ*�\v��SS�L>T�<����(�LrD�'`ը�kX�B�ވ�c��ٵp�z^Ft?K%֢�ڰ"@�5-]�jtfr�@����w/���]r�T��-�� ���Y���Uy�֟Y�Y�o��̂7�)�д��S��	M>�xI�Zf4W�[�~ǏW{r*���g�A�m�ņ����{`=���|f�MYT��
� �=
o�O^�3�MJsɻ����:�)�F*5!k0��l���qtJ]�x�Hd��"�B�e�G�ƈM�NǢщ���
k�c1����e���!�"�R�#�d��Ι�cM�0<ZP� [N���L0F�2���K<����c9p��`���h�!�(�����5������W�#�\�M�a��y�Aمq����E�+Y�S�@ꬹ��;\����r� ��:�uY�#��53b��D1J ���7 �SQ-�p�&��<�Ŭ����G7l�·Qw�o'�����,tAD�	`�с��l�}�ƍ��E��WJ֗�aE���5R�X8	_��/hς��� A�7�[�Ȃ�5u+Nv��K�]'=�#��~�̒e��E�ʍ*� ��#,�s9�:�b�0'-b�U���rS7M |D����]�k8a�A��2�[l[�P  @ɐ�	WN�����(�f0��i�8�L��ܣ�վ���Z΂6p_��h.td�^|�"���Uq�D�#}�����4��k .r�1��Y��E�zn"�G�Gb�I'�l�\g^u�����a����)�5\W:�BԪ���%�;�Ĉ��RM� ��͹e��}������.')/��&��(���W�^���
�ԫ����R���Ǘ�T/��w��aH��λ�,�����#������	�SoUj�j�q;v�(�(���_#�NmV�}[�P/`ܳ������:[O��;{������˛;�:��`�Eji�v�1��kij�$�eNsxNk���V 3�-s��Tb�	����M�ݏ�� G@�� D���lJSlR�������>����뿲�[��њ8��Eӟ����4)@E������9=�S�ө�����kVi�劌Ea�u�z`ݯ�Z8ؘ�A��b��
�*|��+�`��{,A�}��	p�zj
x/ĮQ�'�����&q�K3���hؕ��c��"����6�v��τ ω'�\��DVZ��֒c2=��H|hL{ئ��&�+�a��Y����p�NWN��|�u̊@�u�rp�(���*�����W�8er!��*��P軴j��pu@��dKs�����t�R�� �Ѹ�����������.2g�óuo� }m��E�w��K�F9���7��_��dwϹ�_x����z��ﳋ���<~�?jv�}��U٠C�j$�f�K���` �B0r��qfgC��#�q��+5jo�r�,�����?�?� P�+5W�b�v ����C��>ùNu� I���+��R~F�p��0&�vSٲm���׳��dy� �N�{��;�� �s��="�l�u��Q㣎9��*�s�]���`�)^:�9�8�}�&
4lA������quz|��LYX����I��F`7mdY6�ӼD��C�����a�m�n�-��M
�1��,��A�=Ǽl�$E�C�2���F*ܖ��(M]�$�ݻ� �����s��\�\Z�a�>p�D\�z~��h�M�s�"�G�[ν]��˵�{$���䖅ɚ׎i3	c����i�֮Y[�R4٫^��r���f�X �$U%���6Z�s��ru�ީ������4���=��G*�gl�4�.��Gu�+�c�Ԏ��]G6�]���ܺjzjNI�ۚU"
tV��g(;J]6�����'F�gD�"S��bd���5+g��h����>�Q������8���ig�qїf�"+��m��r('�{����n�K6��o���s|���`��%7����g���B<�����=���kO��q��)��h�M����G�S���Xf�m��I�f���E&�;�h��Yw�)H]����@Mf�#J
@4ƸG�ݨ/4"��~-<�c����8��^u�D�BtV�_֭]gC�%ѻ]7����8���*�}(�����8�M�\\��X�p�5r�`�dW)�ߗ���J�xFy����ъ0s���.��)��!���M7�����-Ĺ��Eb�H�!�Ɋ��.F{kxԖ��dD��|����+�(�y���6���0,�c�A����Q��N���kVd���\�R&�����w0�>�>I��(w�~���]cD����� �r�-
-W�]p�bV�6co�	��xp~���Gm�a��Z~t�U��`.���$� ��AEf1�  ����_>��f�֯� ���2.v��[�Ns3^��}���s��E^��;�ӌ���:r��&���:ѫ������7�I��G��n��@hㆍ�B���g�
��B"����]C9��ǎ�:d���L|�3��&���3�E�c�s�?�Q�C�P��[��Y~㙿^���'��3�U���ed/�L\���)C��.C�î`��toW\~Iy���]����w���������̜ݠD���3i"Ӏ�O ���)J}�7�"��[�m+���t�m�(��ǟ�T�0�Y�9�!��k���7�5C�l�sK'm����:���.���O�Je>�����.){� ���s(Z`��z�H�m!c�s��bZEkOw�55-iokY��35;95�f���1���l��� �\񘅚_Զ@
?�f�=�����Y.�E ;	�}Nt�z�p�U0������fm�i��V�Gk��ά$	�W�v�ԉg�~��yȐ��_�<p�j���� �0�&��Nv��%2�f��?�u5Z�����P%J����y�����묑�p�X젆{���W䀉�:<�&O�X�4ȏ��,p#2��+���'���$��|��f��ŭ��hHFmH�׺#�Z���P,���hwyAy�;����LYٹ�>~7��S�d�H�oq��� ���4�R��o~�k��^-���T�[���jg]~�[�Z^��ז�?�g�nw<�mP�A�V�C�!D������ �F<JZ��8��  E2EΕ@sx�L���o�zWWw�������,��?+W_s�2%/�B�Ї>ԟ��Iב!�0��1A�=A�Z�'��re<��,�N�`���'�]r%�������s��\�<q��g�"xe}
���c�D�fs�@���x0������p���Y%�H����}�/^��姝rFy�+^Y�h��S@l ��LCM�`.�����z� ��/|W9�|Ԁܒ�����O˿~���ŗ]\���^^�җ���)e��@\��2"��������1F[��`&����Fr7�����gRWn�����<��ǔ��;O�㧛����/?����)�_o��g?����d D�.���[�顇�NųPۑ�B7�3G�VdK�VN8�1�|nڷ��m����"`����/7(�0�[���T���2 G�FBH�k�)�9Aw����t$$�6�80���	7#�0md����;��FH�<���,�|��5kVK�����z��t�4k�7.�q1T-]*'�k�T}P��1ԦO�1����隉���o޶�����O,l���.=�$�?K��sP]jQ+�ӡ�쇤�U�_�!���Z$�-H@���uJhJ)f%�G�꿦q�,�\[�d�@��s�%-�[յ��Uʋ��&1�Mڔ*�������EΌ7ͭP���N�ؠ6�A!�\|ݧXA����� ���Q�U�����L[�����l��W��n6j^EG��W�0�6�����ʿai�\�"�(��:���)�(Hbh�5��x�1�S�u��Ț�Bn����b���t�A�b�]b|?��ϗ�k��S!�'{\yƯ�jy�c��0Y��S2ر	ևQ&)�}�-�_s
��b�Fj�Ҁ(BI�w��]峟�����[F�Mox���*��c�w��Ю��~��_�N1
J���-\��w1,�M���﨤�9�h��\JΆ��~G׃��U��O}�S��`����7O~��o��o����P�0�s��7;Tw�����6n��1�l�w�(ѝ�9I:v��7,��_�:�A�Q����z�<G�v��U�o2`��><��$k����9�*���R3�p}�D���[���1jGy�J9\Z�+��s_��tZ��R~vy�+^%��,3�DQѧ��l�A{QǨW!���! HˬD�	Q7	%J�& �(��/{�����|�|�k_4�x�@ �����	m�/�5�3�� L(�}�.a"@�ƅK<\���nUN�}j�E߇�OpG��QɈ��/��Mo����/}ы�o<��]�d�^%��;�f�V;�ě���E��\	�����v_��.�j<b�._�W�����{�k�����g=�\p�N�@0ޛ����c7��tEE�f���EFޭ���&��Q�ct��ro�_��<C��==�����(�'��D5u�n5kss��ʎ�[�B��|:��qf�z���v�Ye��#$|.eUg9z`E�_�Z˞ܾSh#*�y���F�ygg�Ԟ��wL)#8���ۥY�Җ��`�R����t��^m��8�J����R��n���C��
�*`Ӯu���Z6ϵw�L�(�F��S,LO/���X��4ף��hS_��ζ7u��gm�T���x�C2'�v��_�� ���Et��,����0�Χ9R0FD���}���>�A	|r���?F�J��Q1P��F��2t@�����@`!���U'O�������ߺ��{�x�i�'�F�ta���X���u���r��w8iަ#�*��v[y�{�S�p��	�7�?����'?�I�]Kz�Bʑf앺�8�Ǹ�u~Ƀb,뽭�?ijD���0�P�W��6�����˵W_S���w�?|��G�5������け�#v��=�U��]>v�q��f���1��Q}a��44��	eF�WYk��|����r�i'�����=�}��l�S�����W��`�|5)(޹c���:w�I�9�`�i`�'��:U46D�-����s�9�%/y����֝[�>���O�����	,�r�-e@,X6�����Q�,U@��o${c��@���@қQXV�����ٟ�o~�>�)ǟR^���_{��wV�����}2�u��l�"MX���H��T@@^��WEA�
�Q`���.�{6�d�'�$�������s��$d���/����i�߷�{��<�9�9G �Գn��qt4REc�����5ϛ�= x�!�B�㔜VҏyHB �6lfֵT�<��ԭ��qLz�m۷��o�)��o6v�+_��i�V*,v��a{�8���"�����X?=;Vh�6 nm��B�T|�WB������U�
��mo+�v��!@���b:^���/|���"U��ߝg�Y�d�&m#3�� ����(�}�`.ќ8�e�|�	������2=���?��Ŀ�1_��/��������o��y�p��sŚ5/�{�C��uk���M�'!ǂ����=�ۤB���'��L��ic���T� ��ฺ��:�4=���h�l`S߯\��2SYkv���j�$�j��~��B�BQE���6�Y�\��='��:Ӷڊ3��^�׽���?���Kw'~r|pH&'L:M�s�������$C�$��=�mzJ��(-oa��2}t)�&'���bB����_����$N�Z�ʻL��C�@A�\o6�a�>��Ԉ1���DS�E����m,4��B�U_�ܩ.��-|�9��8�E'�-��N@A����F�~�����[K�����p��X���b"x2+)0(G_��2����1�P�#6}a�:�WT��ب Ԅ�}�R�C�"��{X�������Z�<�L�?>��Ϛ�MZ�y�?����#4]��j��эZ��6�.��b���$����6{-jHN	'ѯ��ze������W_}U���ß�����Oz�Q]��o�-�},�
4�Yt�^�M�@���߭��uFX0��# ��m�7-�����Y����uo|����p��x
Z���������X}�.U��RJ��ߔ�����`l��s{�̨�2mN�<s�����Έl>k١Ř6�~C�z�W�c���\?��O�O�&�(,��~8'�ɣ16�i�TNF*����pČEt��"pxpƷVh�jE������r��,:BcmSذnCx�ަ0���~�Q0 ':��ލ,�����bȰ;�
=o���x�C��ט�P1F�b�,��L�5"p�q�i����~�{����߳=�u�]� ������Q^ &Ԁ����%v5��6��AIF��}P�=����q]O�2�w	;w�1AK���������
�u�c*Z��
�eL]�[1P����9������jD"^�;c0D�X	̭����S2��K=�% �Y���!!���X�
���[��Ă�
'Z�p��&�@<'<���lN?�q	���zV�Q�k����;�����I��WBimhkX�5�84V
�L�h�e(�7X]+18���W麫�D���2�: [a3�p4��ֶ�0Cp�}Eo,��T�i����*`t����z��Aj���P�Dˋ���]����o�@AK4+,�V���� �8�s��|�e!&#��������Ђ�c��]�)�����`�0��!nR�k��#̻��7iW�6;'�`��h1��M'o��b"&���J1�q�&�x�#��C�S��v��	Q�0!����m��N �}Y{x���������`�d�j��{�S��r-�	�
  �	���W�N:�|$�J*�Grue(���7�Q��!�mwtt�w��]���H^��b
eX�'����}�� �<����`���!ާ8C�e���_'�Gv��Z/�y�o�NǴg�>�5����6���֮�HBeez��F��Lw1��i؊�H~:�cO�0^*'K]��}�c�G��V�-��@�bZX  �.�kC�l��Wҧ��O�V�g�LN���Aea-׸<S8�%V$o����#�/0����N�@<��0�ˏ<<F�^�%Y&@-��v?�v�.�[�����/��𪗿2�џ��i�(`��tl?;�����>>I�d@�h�b5c��,-YL���Mp�ҵP�c�ٻ'<�9�o~�,͛�%�M	5��d���_y��^RB����VX`����w6O��x�R��:> ᳔�H��^U4_)��@Mzc�v�1`�9�i	5��!Ȥ�[�f15=����+|�_�_wC��j�|���Zc�E��E��*YA���*��Yi	 �F�QY�:�)���7[� PT-cW���lLo�Cb�j[B��u�is9W�s+<W"�H�om���h��?Z�nU�)����_bd����ҕE��C"��e"h7��l���`���i�����pH5���*6z], !2d���lڸ��/��:�֨h:�CG����[mݟiat��RQT��|Ϳ�vX��nl¹N?�t9�W�g=�Y>�/T+ �c���D�q�
�%=���lI�G��l_��2��Z�'�2G�S�3\pAx�v����`�V%���h�x�'!p��*ɀ*kc���F��[ ��X������&�>7H�0%�8x(���_����H�3 ��.1Գ����m>TҎ���Ђ�:͉����t���b���s��}�mZg�r�SGȣV m�Hzk�i���4��ԥ,5?�	`(^kb��Lꁅ։9F6�O��իW��un����G�-�D��/!�;�}8m2�$
H�n�Rs�J0�,O���/W��6�����p��m��yn\S%�!��5 K�cU�� >���%���3F���@�zC���3��Ʊ9MB�+��2�1�>�g4W�p��`AGSa���(�a�j��Jsg1��J)뎎�d~����ג� g�<�+������{FG%*���8�T:֦M%����IB(�QB�Hy��X�]{wk*S=�6+����lEE�;�}
��ޥU �M#��oL�h(#!���]k
U
5��.�0��o^����[T	�^��AkN\*S2V�����s/8o���XɯG�2������l8ĹI����L�n".R1j��|����<5���.+��E����)ۮQuA,�]E��Vm���[�p�ֱ.�)�4V*d�*ۻC�:��H,����СA�Y�D�<o����G�'����
��;��賐�t�*�-x����S�ozH��zr�i1�hbV���Si��՚0ӣ�
�+�_s�:�U�}Ƶ'�v���R�9Ҙq5��u�pL�� Q����Ub��:OȋN��"6���E$4AX���l��y]PtTI�=,�!��7^] $�&���D�_���ݫ������>��O�hLH3M�li
�[�K����5�Ѧ��	0�S�U��R�;Y�vӦMV����
���1����z�i~��x3�4!�:\�,%���Yx�LӞE���d�5Klj�J�0Ga�`o�3��{D�b��r%�+���c6&M��`0�� +U��_������"2,��*]먞�q=�&��0��ZƖp��C}`�y���Y�(�_�m��Y�К�q��B�eec� J���^d�?�>�yr}��(9n=̖K���O�ح�>�ɮ�Қ12��}��c
�֯2 ��G�,��Y��Vh�8��5���5fn�b霚�V����*%ot:���^r���M��>=۴������T���>[u��������(�7�RY ��%��p�A;I��G��5+$�өoO]O/g��<�I�O��-�,D�O�s�Y����y�G	-U\aHn��v�ko���]�SB�i�
mU�����޿׼
u��x��(��RG^�J�T��bMEi25�����-#�^�ۤ����ᡧ���-��h�?B�I^Y�&��k���0YnҸ$�n�Y����h[�畧aU���<E��}��Ʈ�ƄU+�'m4�����Ru�.��Y��?Q����W��z���z�,;\��hH���w���jO�H�� ��A`�,!s�bw 0ǩ6�!�EV�L�T9٘�9����cQ��"dyHZ���~Y���9}cì։��ԛv_��	��|((�a>�a%�u>���"t34aiuq�m��?�����m�5.������f�ׅ���*L���\�bO����,%g�q0Ry���
YS-QT�ؾ�LiLW�\m�0��{��c-��I�o��ڻ��U��a�{�=& �X��&NN1ǙF����}�{���\e6oTfԘ�s꿥���X�V?S
��m�f�[���٪�D���4�3b\�0.󝂅J+����ˎ�⾱�G�i��c8 �ՎP����5���q��Th���?xP�̈́tB\��[���re��g��e
�K�#��a��笥F������w*kmO�Q�|,%��A�Bb�=*e��Nw^���+Wo
���_+E^i�ej�ºl�R�bq�QezOR�3�a� h����>�|a1ǁC�۲l�Iw�i��;��8����,&���N�N�qn��%p�U�b{NvJ==]��ݠ0ح��jq�*ղs�W=!�Â�%+6OftA ��γ�H�/vH[����VNSG9�u��*v0�B�h�_PL�ea��D����R7�(��O�L�ڸ�T��0F�¸��`_�#$��� �B��b�ttJk�"���:�<�.��!N�D�E���p�������_ �N�<a�s C�jF1V�W�Z��hhRE�n	7�|�;2i|2y8�48��B�{���.H��&��T�>a?>��[����!,�2T���q�F�K�V��< �t
g���`Ȓ�e1�g��f[ݨ�7%˘��\�>i�p�8�z�Z��6U�����LQr@Λ�P�B-���B�dʄ��6������i���_ ,�6,iNY֘��f*�c�b/�f�o��H�ta�3�}b S� ����jx��0��@����;��c�L`��ޝ�k���ya�`�x��t,k>��x[:�g��{��)��8��y�'1��LZsd1�y��z���5UO��m��:�e����Z���	t*�ӔW�3��?��OOz��4��"��)ՠKH� ��2G�,E{8j ��p׸a�ꉍJ'h����.U����p��+�?}�?Þ�]�6�Q��C�5W�j��5�r;��S�m���w�Non���������8�Z`%�DT�ܯ�8}7eU8�yr%W�9�'�\O�N��y�����b�"�E(��'����R{�RT�����k�AZx�G������ک�8(dF��
��g�Lm)�5^PB�8���Ǳ��>&-���>,ɀ�&�8Y,��$87����� 3�]6�Z�j��Tpl`l��Ο�EJ7UU�J[�y���} =
�����k(.��|}�̈� �����&���E�y��X�턔��g		�������cP�� ���غ � �� ����.վq Xb�e�B��\EP�j礔~�����g,�*�Q��|�X��㥦�	�azd% �~��= �ZckU��1�vP�$
��O���`bj~�����yy���,���Ǆy6),g� �̠��6�H�B؀9zqYX���5�盐S�o<'�HxU�����Z��b�3)��@QbL�`"=�b�\�a�#�7@�_�M��[z��S���̰1�P����kO�a/�Y���`����ÊN+�y�� 9p^��J��3mU|��=�浘�5@,F��Zix�u��>��G��j�ڶt�B����	m߼6��٠$�Xd}��
����A7TR�Uޫ����{D)���f�K��![?j`x�KW_n��P��2�!f��ZC���x/�o�u���[�w�7u�[�_�E�XAK5-�4ĳ�,�{*vI��.,f�.��c���X���.�3�"� �`q"L�:�yȪ��:�حӡDb�d-�4,$d�R�Q��Ѥ��)�sBd�>ȓHQ�Gk>�zP �h��筁'���X�V�A3#m4|�
�����u\�.Bl�Z� Mr���!4�^����hw��Km_D��0s���pOW�
-�T�P�L
���xS��	-�� r��p��R��Pd�w��F&��6'�k�Щ�c���9y�S� �rz"qO�z��K��"�lb����.^5�����{������h;�r*�w�
X�H��I��6�\a�O  ��3e��t[�@�݋�e���-��9ՔM��;�s>~oLU �p�Ř*H]� w�"-��6��0cccAz�q�Tp��޳h_�<$�	���XQ�BČ�%�b�*L�����q��92 !��5^��⁉����U�6�y���N��r��A���4R���Щ
	�A�q���=S�A���ФƊ2�nL�kгCr�=�4��o�xX=��q|���Y�M#Ú�B�C�'�R� ^����Eǂ6vT`fh���Oh�j��w�yW8�ÛCI��i+����1S����5>!F����eZ�bX96��*�h��-��@!Xt�m�+Ú�N��W
��BlϘ����R��B���H�@AKm�^-&���a%��1?�1&<�u�t�'��5���O�cL��CN�Ķ��7�&|�+��~;GC� ғU�+�	PЩ��P��@+U1�Qqz�"�+,��\��m��?v�83����. �-b29�D���5�S�K�Q�;:v�d���4=���w�Q�Q���^�	Ǐ;Z�g7�d�=����8Zf�y,���a+@f��^,R�χ&qq�mщ���I7�[�B���>vߑ���5�oK��}��y��7��&6g1h�'c✝��yR[cȘ��Q"(�eH�2�vW[��A��:6 �r��2 �u�0WN���|���SQ���Ƌqdl�����s<����W�M�#� ޏ#U+Uc3��L������yoe)�����9Q�P����
4�ƨ�FU.�_׏��@��n��t\� �\���ay`���J`&�͚��g�y��-3&y8��f�������y�`i�Vx��@��B���)�����;��+�d��٘iz1���e���#���{������.��xm���N�ْhχ����C��F1�e
��Z�\��NZG�drX�yM(4x5g2*}\׌�[O�1s��t��LϠ�V4"�Yh�s���
�I������MX�XNGs�M4�Uv���T��Kf�û8���Z ��%�;}��E�w�I�����T�O� ?���T3��K,P>����ź�k$\v���U,5RFBa�X'�e\)��zD5.Cǭ�-x��j8K�rQ������g�x�p
�p}Ik��O�<R��6��V�>��	���4Lp)�&�[��Sh���5\�!zv�쒓	���u���H�[�5���!��!�P�a�����rᑵ欂e8 N�b61�M@E�0���Y�L�da �*���ļD��Z1,:�o�����&\j�Fکs8���;�.@�l�(�5]�捥�+�Ac�T�29O�lM`�+�;;e9�̱Gc3��D��PQiF%������-��!�gc���³�����C��9�I�	�kd�6Sk�ڹ�Lԗ�����ۋ��Ľ|��Xڈ�f�)~>/>�l��d<\b��f����>~H���y����k�L����C�'�6y�D��J�O!s�.�-I��8v�Ҕچ�4N������͕3�e`�4wKsڠP�Q�w� �|���r�����tK���y����Ѫv=1E��XN�h�fB�F�+��!<%���
ڦ!S��ie���PѬH�R����@AKn ���&d�]��F����+�K���N
(�;��'��6��zBP���m�:wo۶#�t�-V�xÆM�[h�@�e�x��T�bU�%��ߧ�"���]~�(Mr�����ڽzuaB�r��{�Nӄ�Z�y!�MKB��>_c<��zM�`��T�����Cv��A�bIx29m���les���@�ĺz�����!���[@�Wh��"����DƒQL/�e�3^<͏U'ܥ����؝];��p�~���(H�i6��k"�@Hc�ӵh�l=� �Ξ�w�{c����8�t��u��a�)����l�����K9b;��Trމ�I��H�J!90�E �Sf��ya��c�%��J�i� �F���.$9 �Gۦp�}VV@����c���?kH )|EƝe2j�꘣�-��u�35����v���{[���J,��.n{�%��n��ɧ�b�=���O�Y�� ��o� �Tr ۧ��Tj<C���N�iKڌT��P��^��.��k�ǅg��9�߳D�>}��bk27�U}zLZ�	�?Kݻ�p�Ԇ�V�U��:���
1.WH��i*t�f�<cZVu���aeRm��䩭�Ą���gp:�-��V�BU�y�A�9�T�m.��&_���"����D�o'ydX ��%�3�0sr�(i�"SJ��h`�K��/�?�����yO�yh�Ʉ�d1ѫ�����b���J�S�y��y^�M7x4�q���?���Xh�Cc�����@O#a"Տ��ۢAB8pZm�
Uid����mtM�Ky;�6D��Fw�i��8��Y�q ���R��Ս���SB���i4�3�1�U�C=��֠����r�E��:䎒�^��
����Y��2G
��9ǥ��t<��7����|�SB��?���l��{aƔ���U-��ǜ`���ԯʝ���[o.9۽���:Yh3�^�c��6��J)�t&'T�!9H}�F��k���R��f��7�l"�DN���k�9s�~��R`�z5s0��;�j)��MX+���+��9%�ם��� E�DH��D�`i#]��f�lS��������XR0�j���f��ZS[a-W(�ȵ{�x��b �����b�A����� ��Y�����0^�@�?faY�LbMB�]>�;Qǅ�l�s�9�?؁2z��8}�TLP6�c[\I] 
ࢗB�Y��b�[aOke��Q�;�6!��w�czʘ��>)��
��ԉ��6v %B�����)g#d�727gTyZE �1ZZ~c���C�e��<T��t=e}c�̳6+��(p���S������tZ)O_��~o�K2�C���?�[�,2�}\��*5kEG
}����fa{hk�O,���p� h�C&'Y��s��&IG�2���py�X��?�c=�����C| ����Z*���&Y_��[�O-p,v��Y�Z�Ȩ����^��%'�T	���
�J�3V�����Z-6jv*@DL~B�V�̜�ZX�ݠj�̠܍��:1�!����B�.1Z�}��#��4EֿK��t��� �(�6��}^u�uUB���]�s���(�������vE<d�[��<����,��)p,�c��6�)��a�Ү��;��4�d����-�1%�
���s��5@(�Ȇs��S�I(��� ����y��X�ބ�f�,6�e�X�j}�\���Ӛ::L�'C�@��V)]��v�R���!�n\-�-��A0�{���=��3�9�8I��R�?m)|.��plv�8G�[��F�Bx0܋l�9ψL�S lm��,�rR&�EG4A�"�� ~NO8��@6���w�c�%h���Ɣ��զ�N�Wm(�Z��~̇�d�
���3}����SĀ�X��LKgE%��q�Ԑ��z~�<�0�����&"1�)��Н5�as��F!!��R#x1{q�z�3�2�1y0h�>��\��q��L'��8
�y�?B`*�<�k	k׫@�>�bE{�l���kDUC��3��k�)���.��y�Jk��h>w?����z.F���Z:���I���(����
vڦ�;s��Y�m�Ȑ��S����d���'���-��VN��"KZ1��(�Wf��,�S����O��H���Y	SYgi���VT�����"b���G�EbpD��Ic�(k-�c�:蹤�#��7�	�y8�_Rc'a��XM�+^|3��_���'�����ݩe9�˴� �\���:�&��v��<%6�
�y� �D���P;O�P"$��x,����{[ T�gO�Ŵ$�w�'���!N�6�9�h�>�ut|�\x�Ha�8�E;�a7��v��e�%ǏӤT�iY(��R���qL@P�;+G&Z�nL��Ff<���bEa��ϑÇÀD�h˘#n�/��X����Y�]#u^��\��T���#����
S�{r��1��)���4.q,>���_�yĴ`�ʅP�]����=ލ������ d�bj2�(���"*O�!z�U� B ���R��'�Y<�@���S�,L��}��!x���yd��+|m�Zx`�`I9�d�{��Ajݢ�M���p���;��9�9atH�7�*Nb�z/6#TxN��-��9_�b�{�5��bC]/�ؾ\}��<���������t?Sb+��T��C��{(�X���e8��>qn[i6p����2U��V1�C\�l������"΍E��w>���_��Y �����e�ͪ����t,���9�yp�p����?���|2�JZ �����(��z[����Κ�a�������Da�� L�zB�Sa7ճa12��T�l]���q�,z���ݸ�C�[���	�n���K�Z0
�>p2�p8�"CםD��>������)��Hz���iD�]��T��}�_�������*�j�;�_Q��Z
1[ۍ�f6'��i
�Y���r�پ: �2�gi�l��h+�ꌢ��k '��A2U���ݪ��9C�VJ���Z�ZJ���h��+��a���L���c�����k��O���ggb8_bK�%�����&�/6��v)���g؆Q�?�<dU�܉�_<�bsjߛ��q�������!�2�4�&��K�^�#�<��t��	���"|�O�\�c�F�O-I\�7al��&t�:�*zz@E	�l��jz>����f�����,4g� �7��2��'}� ��=&`��R[�poF�s�{���7g� ����'�����w�*��fݪp�m*�I�#5MUx�Fb4]ua�ºzfi��6�_�?[IP?->d� &��7�gA���X`U�ft�I�K����8�悼N�f3Ǳ�=��O^�|�o.�A���=���%�V�Wu_��\ȴb#jYC8#���ÁTjW9<�k,QK�4�v�刔Y���7�q��N3�H�a-��	Q=�s\��N�+����׀ӈp�bW��s�-��M��xT����ض��S8��xB8^�e��x��B_b}��ME��oN =���H��'2L��ς.�ݴ�zD���xD�� �!mwЄ��5���U�uE|ĳ���bz?mF
Ѧ�Ҭ%FG?�g��ɝB�bk @���#��l��N1���38!�����ҽ���1��0��Rkn ������%A��	���iZ���
4 ʱZ��jDI��_Pۇ0���a찏�nG[F����r��=����Ү��j��+  ��?����~M��wc�q��b}R)��A���C��h]�<HvЖj�-����}���4������v���w�zF���+\j� ��F^�M�҂D�R�x�S�����a�$8Osݴ�Uř�+��s��	k�Ú��P�K�]*�A�U����"���B�#�/���V�숊����t~/l��^,��i��z�.�xZ!�.�����}ž����g �x*>"�� h��쏸�f��փ��nYˈ2�	p���,���{�� #�#(YX�ٱAp/�/�({�V��k���1-bc�Y��aR��D8�l�E'!U�E�Ђ�i��Y�'��y���!��qH��4 >@����c�wM�9&�ʹ�Q���bт;��@r2��)�s���S�������<�I{�:4�F[�cw�w�鞽 �����l9�@hA�4q�<? �&�Lwoc����G d 1
dM�p���b>�����U>N��(
Gdl��1�ϓ�!�ᤍH/X;�~1#$a-I;X͝ �����AC��Xd�(Ð�#.w���<~�S�u�-�yikBh� W_����D���c,noS�y���X�L؋�Q�����#a: ��#�Q26����BPr�tN�>~�]�96��i��E&A8@�����]��ەЊdp�K�|MNP���<  �QIDAT����S���;q=p`�l�ݷ��g�{S��Z��D��k�������5Aw٠67�����;���]�����D1��#BK�T���]>L��k��~����>��F�H����L��[NSe�U{�-��RbbyJL��d�M�n��o�_#C�1��z�̍R��� �`�m��-��siZy�>�ZZ�3�_Y�d���փX���z�z�ƞ*�x�-����h~��':�%��?fv��b���0��/���Xf[�%b�#r��ZڲP�*��UW�����a\�[��|��J�E	��
\�;�K�W{r�؉DPV�OM�����(�?�c!�M��0�ʛZ����٥�:)�"F�M��D� -��`��V
��n�r�B��n�������Y&�93�#f��qn�8�Z�=$��އ檌��8@��,~��B�Aڴ��C�EC6O���N.�pR�y�j����J�휓(ݮ����{I"�W�8���W�;D)�ź��rCדBmV����<����#c�J%$@�8de�/4^�NfG��@+D(օ���!��P�s3�/��� ��^�VSd�&�a�8������.��v#��R;3_���� ��B�X	;�դ/r��6H�"5C����z��qc��c@��Y�l�,ܨ�_&\�qM�l���Т���	��;��Xh\��I�gDL)Lt�
`�l��� 6!�K�.�����NaD��k�BJ'�Q��C�:�[6�s�;GÂmUEZ�J�[U�i�1E����Jr*�JK2����6@+�c��e��蔛V*f��Y �]�-�ތJA �5��4�-�;��f�/��� h�cl���ؖ��3u�rl�I�CB�N>��N{L�Ĭw����X�ww <���*��u6�=��MW�֮�V4��?��Jv}�BN���V����$6(�M��$����7c�"��!˚��ݼ3ש5lE��5Pod�p;x?WI����/ӭ\��t�R��yZͯ��Ѝ�Y5^�C�E����4�>�g����2V �{eo��,U^Z+��؀��D`����~F%@V�l�-�8�$�A�P!��Wc@t����������bl�s�{1A��D�I���8l e��H׏�S�Ϝ�ۡ���#��<ܳe��H���V���&��>ll8?����p���3�ź�� �o����Mi�;�is�怋�S�yҌ%͜u����h@���vʘm���.������3N����UșK0cn�q锬J7 V���W�e\ʜ�t���ݴ� @Ș�]��O���"�SK�nѩ��أ^	��r�~�硒򤮕����32Kc�`�V)[��n�:+_���'M��Y(��Bm��A3���=�]ʨ۰~�B�{C��1��Y����è2� ^T��Lu�l��Cp��m�0�f˞��������0tlR�~��e���2l&��kQ��1} ��e��~�ᶅ5:�X\h�3�"Uka[쌀������E��eZ~O�<��֌�k�]��ND��[��Z4O',�S�`��\�pӍ7�Zo��Z��M��,��_�bͭ��k �u�צo��#�a!�F�*Nƅ�/��9�G�<s&i��-ю�z,�ӟo�I�����,�bm�ba,�)h!��n�@��PV���G�G��)��}.�R����M"tc`��|a�iV7{x+�:\��>Q(��A?����9�� d���� |��g��r Y8����7�U��75�8�g��,�ëÜ�@pN�H�9��q�~���C6�sG0c�$�&��YB˄#5]=���H/)��q(��ҢX�F���s�R�;ƒ
�V����@�i���:D��6z��� ���(�%������K`J�o���B�rʤ�{c�q���2��`>U*%�����j�9_	[� ��'d��u���l��`�	����]����`�O�8����Ш�6�� ���`%�� [�P4��0J�4�A���*e�L{)+L(v0���?�;ƛ�^�p�\�R��!c�Rsc�����:�z��G:�5�K�B`K�U���U��9�Ը��ޙ.�D����g�a�,/�j���@v#�xذJ�����ki�`���[������!��z�o�9�@A?���`w�Gm�׌�&�|Bl�A��c�"7�'�;5E����g���g�,{V^��lQ����� �>%Z�U��ږ)�L����H� �3y�������+�x�q����F�H:~w�v��K��S}cq�6�c%P�D�8+q�nF�nD�1u! j�P��"���Uh�?K�2O�aG*��6��NL���VցM�����<�ԑu��������0P�R�q��4 �3�]��1M�<���p{-F��gX ���?s�B!�"�gS+��3���sT��Cu_�����@(}�,��NZ*����*�04��΍��׌5�t�g_"p��&dc�gؗ�U�#4
�R�NF�A�K��ZN��,]��~,�^<�tE�Km³V|1�u�����`�(������З���n�#4N ��W����٫�;K�}�<4�s��K!2�?U}��5�S�i��e�}�LG�G�B��%7�j,;K��2�����Q*�#t�Z)�Y����1��[&1r�Bu�	�Dpl�?E��--9�doH���--�{�l!כZy����h�5�9j���1�k��U�m��P��ιj�
�@kvK�y
�������CG=*��Fj|f�C����S��0�?o�\��]Z+R����y��
�p!��ò�Y�2g<��FW���ߵ8��X�n,�A��<8��J;p���?�i�ҹ�G,lw~,��������p8S��:iE��Agה�6J�N�@͡^�T�U��De��QN�8m	��cD���ءm��"��_zo��S�ARdX,d�\#�!w���P�;i������:�F�XY`�Z��t]Մ��0�U��J�<۝ǝ8H(�ZسYv��:,��$�S"��\o���Y@)
G��l�I��������� �D����v�r4VO�ГbP��;+��D �k`^�%��.�N���c̈́]J+�ؔ[��|<���Z]�U)�ɔ��F�W��zp���o)�1۪l¢.Pij�3l�g��qK���1�H`dʰ7:�d=lF�kf�k�8G����	6�V���F ��Q�)�c�(�1F1�.�0aI��0��s����H
�p��I#Ľ�,�M=�`S���k�{�\����V�-ia|m�fJ�e�����?�{hnn���g�a�V��k�w�
�mٲ%<�1���
�}��{A<�F��8�J��0T�
�ͭ(���¥ R�"g�[�3�3k����������=�ݡIM�a�����+�g�s�`X�fe���������<��P}c+RT�K	 ��C:�dr����0�"V؞)�w���Dz�h�b!V[�";m����-4~�H=��6����-q�y�� �
�}�~i��X=�P�=� ia��8��pG*&�&~�%\_���l'Td�;����v�����;)}k�D�֎҄��Fr$���[Q4�ݺ%����i����ޝ���'T���8|֜���K±,�B�J0s��#�h܀��䜽f!�&��L����.��S,��-A�'��ZX��F"�gfḭ&.�����J�~P���ǰ*��3/�6����.&:&_|u}�Dৌ�����c�#n.���85�4�J���-rL,J��W輴,��/��v�&t��0��s�J�� ��؂6
���>+2*\D��CC���U����������R�Ī>sM�i9dKڜ <Q�,/�Z�;�I�XB��^��u`0:^jN�E�jĪ�q�Cr�5zOE���?�F�b��Π�%�a#��u �E�c�ߺ�j�'���:vT��1;"aJ���(<5*��3A��	�E�?%�P�F	@�XL[�����\���s�0$1m���ha;�/�1X`�*�lP�cY4 9�� 4O���<?z\L���[���v���Թ٠4��5ջ$+�B;��q����y�*K3N�q����@�F�{(�Ƚ�*nj�^c�uo��L��7�>ۣ�����p�S���/�;���#�C�ګ4�4Z�����o�!�ض-\r�B'M�0�~M�w����9�uJ�02@�n�Nئf�"xZ.Y*R�Q��_��������p�:�i� h�#N�<m��P��;M'-�=N�
}��z��G�q�WSN)�\�9P��dd?�l����J�^�0�#M��bѮ��l�L'��%�0�^Rx�=B� ����W-5���s_X��M�������خV��"x,�r���1%��z9&���%���~k/��݂37h����k����d�2�%����;����Y ��G@�'ڒ��� o��uv�ޡ�-4�ԫ�Ƞq�@0�.&鴨�bE�\x�IE%Y1r� کN�����`'l�KYU,�w�_�(ҽ�����] �(�F�0rh���&jt);2'uOh �c�����g+ ���u��gt��'����
�zd�M��5U
}(;�>b3��k|Z����po�um
�H'ҧ��5�Q�l `RN����2hl�u�d�x���0L-�=ٳFA�R��s@)�g�q4��pưڜ��a^��d#8�!U6�5�]�au�t_�H�̙)��
]-�la$�O����y[-䞻��c��a��Uw��������z���'?��p�c��B����K���a�f47p��nR�e�YE�3����fUP�P�xxX̡�dL)��_��	`�p��0^�I�X��z�YB��[:.�@ē���e`�֐�����s",H8p\:�	�|�BJ��:�������駟�ݾ-��8da�;�C_�Æ�kB�f�����2}X}]��w��>@e1V��\�o�>�o�����ϵW��|�������U
L�]'4�6l^jUe�J��<s�
#n7l�g�]��L��, M��z�)�����E�jZ� �G*Х{�>f	c�Tܑ��e�=��j��2�$��J�z��<ОD���e�(��HѴ6X	-�'��~,���a�L�jU��r���^dMw�N��r�H���lh�ĭ�|�C�!�_�1�t��@��P	9K�Q<�
,a�/�8yI������J��{m��P�:>kqoZ��:�[�sm_�,��/�b�-�'2l"�B���Ǚ#J��0�4��=t�D���√����c`����N�3@�}�����ўj�W�^	,��P-c�X&-��9������u�Q�m!L�BY7�;t0Nz�tbӡ�{Ld��ޮ~[a�5�œq�����-Cԁ��gt(?2VSad&u|��͍��;&�0(`�N�YΎ�B��%��d'shC �����tu��n�����2�-��Am�9�k��E�10�D�=��k� a\�8xĘ����N�j��#ǻ����尽�znM���ռ���	mI����nhQ}����}�u⮬�]��(U	��֕X�6����I1���i��ח1W*�  ��hp	ȢAę�/�����1�
�ls�J�h���>r���iYx�s�kl�{�Y�8�֛o
7n�{Nأ��O;=��e/�\~E��G�Z��;wZ�Z���0��")�� v�8���	BM� �E� �ROw��%�_̫V������d@`��z�C�Τ�����ݪ(s���L��S���V{
�J`I�ؖ�����U�t�2��n�N?����jB��{��.{ԣB���Ĭ��5�h|�ll�<�5�]ڗ��v��J,йp�!��{�N�b�"�Ê���5�Ņ
��[o4�����������7�M�P�PW�mf���>)�60x4,�0�Jv"����A�P��C;c�ד��ň�'S�s�����A؄S�S�l��zی������zkk��]��3x������ h�#��S*M*� ��Y����iu&���%�%йq��v ���D��ɗy22��_�����YD�c�"�Z�{^Xl��	Q $���^��A�`ט��p��k��^/}��ڥ���=+,kn	�ݷS�d��;C�~����D�sSr�bW�\k�IV.G���L��Z�r9�Z�1X�~���r�e �����b��W�P��9��|.�Y�z9�>s�k֮7��Z��ش;n�=4�n��8d��7`#X ��=a�}������!sj�C�@ȧ_�cY�L9@�p�T�"�͐�9q� ��a��p��]a@��g�6�_Z�c�n�~[0G�3:��̇��V	l��1��\�#v�c`��/�y 8��Ͽ��O��['��P�0�{F�J���V�����z�5�87�@�m�i2����k`�L:���
g�yv8���6	��۷?|�[�2f�� \z�e� ����ڷo��{��u��E�u�)ï��˃�8&43 ��Ί�0�&h�B*| AXj�j�lܸ�X�Σ��[�V���+��~�/9a͏�;�5�Ҏ]{Cs������B<G�3(=v�[��*5��wBk���燹Ch!��̢�Ȱ@��1Y�ZU�Hk�*�J��V�Bs��H!5l��{��\tX��6Tg^�y�Q"�29��^����� (���=��_ ����>�|�֍ھ��a��ճ��uKT4��(�2@�� ɨ
�b�P&@�F6���G[v`� 3����y�7��C�l/�-���Kuyz�Q���Aa���֬g��9�!�8�£��nиU��3�5b}&�u� �1(;"����0�τ�Q+Ć�͖e�R���bk3�g6���:),��h�� ��#u@�p
�-�-�O��Y ��������0[LC��V2c�g�2�,���F��!4�Xp����%Zt���qR���Hdp���5��)|V1���rv,���\9J���b�ίX"E��#���ж����E���aSxֳ�θo��0��a��[E�2�c�9Ugm�v�0
}N���ؘ�Qe�Q����U|NU����5��iѐ���Ң8A�Ah ��:��a���叺/�^�JZ�M��ۥ]�!���0���8���[o�3hT����u��I�=(m;��?�R�W�[V����^cU�3��u�&BY�6����5�''�3^�c����ȹM[��ik-�����hԅlݺU�`Y��λM\�y�^�,�m�7�:�?��#1���u�Ղ�:.���a�!99&��`��:��
�ӡ����30���E�9.��/�R�FM��2]���r�b
zĜ��|=��~�٦aa�V�6���q\��o�յ6��쐍���}y����cp�IK�ҥ9#�)���½;w�~̯<�Ҿ|�J�>j�A���jc.N:���K�3"�@И5k�.�䒰R��w�����ͷ�e�C؊�9}��v�Ç��l8"�퐀?��"�7����4i�	� 8�ň�ٻ���u�C �F�|Ps��$��n�!��U�����8?JB�5���2�����k�9#pq��C^�\���f.��� �s&02�k���{47~`s�Ea��v�Rg{��}����ٽ�F�ݶ����ф6#e:*w���ԆP�*PI&Yq��p�4Kuu56���L������������G�.t��A���^��&ˤ�?z�Ϙ*6FS#�@/�(����FZ�1���'���8E<K��@��e��$Y��?�5��@��2 �s�̀���\[!TA:A%-�/�O��Y ���O�$���x�2 īA$��,�Ǟ+�L�{ �A�ty@�����SՄ��(��<�k$�C�����������a�������#̕�%D���
����s�Ia]�3�
���6�[�m�j��B�h��Ύ��a	/�8�|���w�1��i��V	����TG�A���F
���D�����g�BA�%²F��19�m�w	���t��"�g�c�(
�>��n��l\���{��9�s�1��o�a,Y5Mqo8�;�u�0A����z��N1D�4�4Ї �H��3�OG1i�t�>���ڑ�����L����ζ�σC dCV=Ԁ�"dw����+׆}���b_Tf��MM]b[z
&íw�c �]��C���B��u�&�(��<hE�(m`)̀ ����lظ>��b��ᬷ)�r�C"��&}8�s����[íw�m��y�i{�ۨ�� �ǝw�i"�U�V���k�B�\cY��Y�ؐ�U�4xͯ��~	x<��QX�0��m>�.�ǥ�u�B�A@�5n�޺�l2�*4� �U�/0dwI�1+pU*���ez�jX ��
����O�~Ŋ�V��@P���a��<x$А��@IG:�E9,V�R�ϙ�n������@bߪ�h��YGŚm�h����%��t��F�%CxL�=(�TS�dL��X���ν��L;�߫����_~�1W��֖Ч�61[Gu�!�X�
���	�ػ���l����(�٭���"��Ex>>�g� �s�گ9ߠ�₋.6�pT��:t��z�}Nj������w&
��1a��ZK�W�Lcݦk]�r�i���s�%��O{��E��r=V���t=�ދ�d�9(�/�S�ke���qڛ�C���bz>�����g[F� ]��{����m-}4��a�Ma'�*-V�-����I.Y<^%�S� E^����bZ�H;���̨��x������V��m}��@�_,�߆��Ц��C,���n��a[\"#�W
�!���_��S�v�=֭�S�PU8��_��R�C9��fD�:3kW]� ]AAuP��̕I��'��,��_-�1��#=á��6l�zn�+�6kml3&e��_��QNF�Q��
?�Z��gF����k�n��.���yv�?��bg�sA�f�s-[*rƥ{�����5�KWQ�p�2|�����D�še��PT�kv9�X�r��1E�3���x�s�㘚B���93eSv�(�s�5�u�ݲ{}x�3�v���OX�v�-�b0��/7�A9��.=˜���L���=���G�K��&��.4}Ǩ�.�,�|Ӎ�5(F�Q�	��u�~݆aL�q�ڵ�
�QШV��Z�P+�F*:E��G=�W��;w)ԣB�
��
v�(<'`�qD r� L��@�L��a�ˠ��bպ�apX��耴-8Sl�?�6 �]����Q1OL��v�ut� �c�f\�k����<e�Be����n^�ѓ	5��� �BF�&P�60��uP�I����U �` �O]͍5������^�98[��Q�z� �v���-l�X�0c����I%psXO�4a\FuM+��5�$� �y*�{׬Xv�Mk�Wi��),x���|-����L��W k����;u�}�b�N]�]�kÖ�N���
3�ܹ�jք\6vR����#�[���\��ZM}u8��L=_�K���!o�!+o�vO,a?ƈ�@2��4��7������y�gP�X����!@���<�ﴍ��F�}��Ko$پ�n��J�-�b��D
�`�K��kB=�� ,JI/�h%#��I^V��e���K�r +����d���8�)��}�c���'�,�`I�_�;�o���]�����+yew�p�V���QQ:' �Bg�X��m@y�@-h� ���p��,a�JEY%VA�= ��uon�!Auv5��e�c1wv��١�ѭ �4*ؘ(�Q��!R�zՑ+q���`h���dVYE	�s�Y���{vW�*iք��7�>�{��fEi�?Zl�J&�܎�k��A�g۽���:���g>M���QN���hPԊM�v��Yao��>���8�so�P��mA�
��
�ᘆ到(�>�����l���"�`��g(y�e�͢l.�A�Y��u�a9�uo��4 �bd*��i�V�S�ʕX��jh��0l,Y|5�0d�Q�yR�Z�Oc��VI܋��n�<B�)[jla��b����@��4�,��u떛&�۶��]�1
�+�k8�a�3c����'A�M�V[+��D�u
gM�v�"m���3o�%�\	a�a4  ��M
Z#X�*� ����PK]�rik�J������_�����-��F �MN��
����55օF����RGH��&���1=�d����)�W�{���y����~�u\@��B�C6?4����Z�	�<����_�П��q@SE��!"̝6�l-�O�.:$ا�Ė�j�o�5�"�Ս��X��p��T]��TM�~M8����ߨ�넴V�z� ����
w���֊+�aE6mۨgz��=��	1˹Wjİ5�铮��4Rht�+��Ƭ�9��iY�|�m�����1��`�i���׹�z��x�6=�6�d�pֱZ��B$�� � +0�l�֋%f^�����j��+�k��vG ��}�����a͖���B禬'^��.׭�Q9MI/DԴ��4W5��U�]�	��L��I����V7K`��Y� �~�F���P6^9��/~�K���U�]���#����	Z�`d�"F�=[�Q6[U���Y�e}��%�r�d�L(�_B�&z,Q�M��Y�I�R�7��Ϙ!��S�b��ۙ���К/|8R�Z�9�q])�U�V!?-^V�_ ����'P�0EA�W;Qj� �����/~�j���(^s���a��i��5�R�N���Z�6¨2���T6,�*�/P�����Ĺ���A�\X?��	�
��M�eF��E�[A����'Mx@@�ki�&��7��bB���ł���Y�&IN}hd�v�V�F�#�u�N!��=��� Ŧ���9Sf��i��ک�>��m,��N�����ڲ����fA׆���9���M�Ӱs�{B��ې B�B;��\v����Dͯ��\d�a�&|���R�� ��WJ��ܱs���+6OʹZ�\�p�"��ׯ�)��p�㺗f�j�n��|V3V�����j��3Ч�V������8&V�g�^����9G�i���Ҁ/��>���{����Wz�54	 H�D���z�ă�֛^}Ku�J���Y<�y�@U]���E5�v��T� SY�`��E�i��J����A��Z� �B���̍m��;�B4M��U��e�j$.�}�����Z�V��~���O���kW��O���x8c�&�Ȇ4Lϵa�ڰR�M�"I��l�� @v\u���Vi,���*�u��5�F����ᱣ�h���=LE���	�h�M� �oVL�%)��Р�?�x����ՑB�s�������=�b�
��y��5�X� Ԛ�����5qwu�t]u5��S���TRA󦦱Ul�6{:�u��T�\�ta��k\�Ț!8Z�^�[�ƒ6(6{����36����\G���v��g��b]�q��Ϣ�%z�_܏e�Ա�s:��z���m�JՔs�|;;�Y>zo��^�a�2MU��r�*��#bK j.(�`x`�i�tw'�g��m�i��%�yq0������L ��e�-
ͱ�.���'TPS�@��Ӡ&�,6u���� �2�B�iRvI��r����!k�X����T�`�hn�U�jG� �Q�'ۤ�M�9Mٝwt�#�#��������'Ѥ��*�!�`P\P�*��8�0 @C�1.`ĊWi�g��,�3T��i��eUZ�u]�1$hDN����V)[H�#2C�D�k;V�� 'ÂM�L�0c�uV��6��s�y٭j�//w@�n�ś���Ε�5Nm%��+�}�{��#�Y���}��^��A?Á����� ����j�j^��ҁu�|P���ѪR"$�g �؄�<$���!2�f4wתHz�={�+�"p'�F��Uh���>���Z<���Zjl���,�0���u$LN�0!��i�FK�E�����H1�U���mPsKU�Ѯ()�Z�!~	XA/�m��C(���
0�ku���0q�	�Jr֑�P܏������|�:�w#b�
z�*cm�.	�3�P�!�^�{wޫ�bT���ׯh����_x�����������}��� 힎I�v��J6ќB�~@�a�&��ö<3#��+Վ���k{��(i�������W���N�  ��DZx � ��!�J�����2�؅�/�jk�Ko��󁭻��t���ʧ<%􉄜��l��xJ�~�JH�V\Y/�'�10�}�2Ϭ_���}������l]@��y5���.�&Ⱦ��q���{^R������]K�=Q{�T��?�c���8T����p��r{ ��?n�o��HhG�+�G�F�w����e�e�=S�\��xI����u��U�
�&XXܭ"6��SoV\[dy��'��%- �0'�����E��Iٶɏ_)�P:ESE����QΛz �R�Z#4J�s"7V,UV�uV�Nj����p��<Te��tl+D'�A�oJ����w�)���r����"�%*�{Wv���� ��XT�kgQ$���d��O���f�P"5�k�{9?NG�Z?���a���#�(ݚ��L$��O�]2�`%��AR��G��<f�J��q@׀�H�`�
 lX�I�B'oB�f���tK3����%���~Z�f��)O�n鼰H�^� p`��(���I�nh�-�u�����wT�r8 �L;�J��?������Ph��<){&+�d��#�
�ɆU�,Ҽ�s���b�	˫T�y38.G���b��R>��%��'���4�G�*��3�e�c��T#�����C�!�N��R�	�CS����z(1D���h4j�_�'=S��l�0��4�$n�@�+�5m�='�5���jn� 1o�^����qB��i\'Z<&��I1����m>' W�y �̧?-�ᖻC�j����u�ݖ��K]�k���c�N��j���� �ֽ���?�� ��j�6#T'W�����zF��}�z�/��n��blm��m��
mP�H���p��������~�-��}��![�ɥ�O1G>;55jʣ�r_W���bw4����Ш�$���!��K�XW�֮ߪ5CϦ�%
��>Q��8�M<�܄	%�LJ;	#&��ǵ����JI�C4�lMæ��Xu��R��V�	�]��֎n�.!��-u�@���	;�
�J�"��bI���^�OG��90>2�qΦU?ش��v���%R`rQI��R�0Y�{���M_��ܾYq�6Ux.�]����/��ɟ�"�e��"b�����Y8��[t��P�E%ڝs�T1�!ЊH����P�X+I���Cr�X\��lrH�q��!���ӄ�X�tl2�X��#��1�yL�"��U�J���Y��W�mi�qܞE�NSM� Nfwk��C�2/�F2��- h����G�HX
�E�Q�d;J9D�t�~��$���B�7YNUrB47-*��,�b��NDǮQ=�)�!�v��$~ެ̰�sq�>MM����N r�.�$A�Ϝ*@�XE�ESQ����K��
�9��z�{�w�)�:W��
z��.���µ���v`�I�19	 ֐�8��u�J9E�T��"�;TPAGR���<+��������0����7���z1d��l�սh�Z�B$��'��1):�J�Ep��
͐�gnIcf�`�d�i
jR�ܗ��F�P=lR2�q.�~C����8�3ij�=�����E�悾����� ,�����o0�:���<��݉,l ˓��ނ��M`�*Y뺭O��kա*d�
9�����n���w@�Ds	�Zk�}˄�g�_��5��CK��0��G�cD gR�B�#z_sKUhY�Y��B��W��ZB&�F�&��V��a/���J�̭cS��J	��xm� u<o,+hgh�f�|�ќAW�f�N�ذ^�v�6DX�&��q*��MU�*��-4��ڍ�	(���g,uz(�)FsF��t1����=�7�7�Ċ��k�l{h����2�jb�YI7��_�K���f�M~�탘�T�׼� h�>��s-q��H-1��Es�,�z��mV@�j�XW(U��ÃS?loj���s�n���>��o\�姉�������ǿ���m;�ٴ|͕e5Z��L �E�(y��iaqA�@t.�RMML���"@Z���vr�_�>;s-,4�{f�0Y���J-rr���ɍ[�i-A���-H�2����)�c�v��+~�K�y�`q�9�ݡ�l�53���f��U�f��Dt^Bl�׊8j�c���9���*cD�$�K�[(H�RݏhM�A=kH��^��҉t��#twxի^^������S��E����ƵXO�!6����ƨScV�=:�.:��g�u��0+S�0�����{��������D�K���Kd�XA(�p���Ӻ� b����e`K��Å���t�ւ6
hr�o�ճ��U��9�Њ�6+,R-�S �Ze�ؘV�8%�K'R�g��)Cԫ��ӷl
�}�U��k�PTqL!۱���w��бgWh_}��-6T�G�ޥ�K�X*����@۴'_�,\��a佧ަ���85i@h�`U��(Qv��h�&���7�ڛ������;?�jOBr���E�;����M�F�C{�RQ_el�lEI�j~r݄�d<J
4J�Bo��PDhXl�ب��lP���$��K�Q�����5�=�Lْ#W*oO����y�y�H��F���	�qғ�8���u��H�
0ʔ#���S�1���NN�R��Q!WD�*�sT	
Uu*� ����I�I�C������3I ��}C��������F'�͖
C*D��m8�|�R؂��f3�Q��PU�jE�oC�u�ze�q٫B���m%�U�1)�6miVv���e S=�T����"K��	�I$nl����MIC{4'������HF�%�V	 �ia��Ȅ���c ��S��:i�3�"mh}��#�-q���U�(���`B=�fT�g�E��x`����sc�u�c/��Ӯ|��_=����>�s=岭���c������W��cfr��u-�[��F�@� � vs �a����@��M��M�^DΆ;;����yfi�����C�����)ձ�-�d�@����xUW��3����(�L���0��݇�!4��ò\�?v�4�� ��1���$f�EP�2\�8�Tk��(t�29*~��w�$�	NNN^[?�`���X(��P�A�����B�����w�����Rײ��*Ԗi���n��J��,0l�n�*o�H�M��p�%熿����xs<�����W�/}ɳ�{�����w�9F�/z��Z]�j�()U8B砇�Ha�RR���5�]��%͇X�:	b�vT��������+X���H���K� �H���{��<�R�ݴ����r�aHN��da`% Δ셃�ƦgT��3������g^&��nQ�ot*�/_��+��e��-���b�z��;L�������e�H�=@�FNw��`-�A��8�R�$(�ac��$�U+���k�B�:=+�1+A�c�?=<����L+ž��o�j��� a@���q��Yh6:кh��&�JJE*��{ի҆�zN�Ū���U��V�a�Rl9��%b�F��Ј�B�z1A%
oRJ ���M�YԼ������.����A��x�l%�����%�O}��#�_�R4z�~i��`6��o��+M���i�
�XSY' 0��-S ߦ����-�P.�1�9�f�@O�0jU��,�8e{�T��\- 3(���Bx�����J������|���ZD=bY9����!�]�9��ӞeD�s
��
4�c�
E[�ѓO��4�c�=U3S���JU̚J���3�:F���pkQESc���PD�?=�\���l&YGK�U�R6�I�4�+Y~=r,�A���+�*�BHG����;�ƪ
�3e#�{�?���=�?~�O����<�����/�����>���V��u����qcqiy�АsJ�@(�"�>�yr�qk]�&���܃|P�v(eCXj�I̯'�y�#�9�BVR���N�[�$��ΒF	0d9f,���̑�?޵�K�������[~�Μv'���C v����5c�p,�
�}���6\G�"E�S�e��]��ء��w�#���O�ݥ�|�$_��ځOJ�FOW��� �i�(t�0��s�>K������3���
&�ʲ�	}��xCx��n��a�V}�j��U��M4l �Ke�v�
5��t�eM�+�k|M���u�BG3�N��&��rD
��\5u-v�8hvχ:K�T���ׇo]��p�_�u��n�fk�4%�4G(��x!Ҧn�2�LY�d �}��_�w�T ת�������7�ax�K^������v�Cb����e��)ۨI���Q#6�D�nlb0tv�W�N8C�)1#ԁjV`���!����0�K�/XIfϘ޻R)��׭Rqʃ�����^���W?W"p�ilJ��T�`ɍf��w��$"G�"�3�kc�
շY	b�W0!��ݡ]"�J��L���1?}mh����J��B �q�́tib����Ⱶ7�Vb{䔩��Nh�[!e���J6+誘�0qbfaa���my8,�${�H�^��/���H�ޞ"1.</��-�T�[��9���`=�R�S�Y��=b?�:P,ۗY�:K���ժk׈)�D,=��,�^� ��3�%J�� <�P�-7�d�A����V�}g�*�K@��U��:ZH[�3�?������#���^1�%#��h�l}���!���`�Mճ"F{��۵W{;�n�����<}Ǻ�+ƚ�jg
�`j�thd��Б�u��x륷o������Zժk��Îl�h����tI%V���W���_dd���#��A�&�G�@���Ukg��Xul�o�+�� @K=<�{�+~�����'�����ӷ�{A�J��i>�ř�rP�-�ژU�<���@�B��5[}g��8@��~9SC/�Ң�o�Zp�ny�ߊ�R|ֲ�&��6��9�nN������S<�Bv[��On� =���뷮�1��Q��l,�� �5&@h�� ��rml�7���S{���p��������K_������:>p4��e/��_���Kj���#ݾM��cd���n}T�I�X�(�N�bAtlٻC�f�s���tw�{�zo���}��t"�{�S���,5�����M�W�P�ޘ�12�{�(�?�q�j��L��.9�^9��pM���k���5��}t��{0|���+ܽ�#,_����;���y�+�o>�2}>�׮T�Φ����-pTר�r�%���O�BS�:wk�,�I@c�t�e��F�~�����o}�{��/YX�^[����s^x�ܧ����`'%����d���#*�)=�e�����Fɡ�Aŉ�.k7�v�U���K�^�r�j�	� ,i\���õ?�>l<�B�v�?��Ԧ���<�4�yv��*2��wy[m�����z1����{Ͻ�н��j[�\�Ju�UȞK1��6�}�c�)H�ݩv���K$EQ��|\�d�K-�FFƄ\��&�� Lw�ҟ������ĳ�۰ hD�ٳC+p3��	�W� e�)L*�/@SZ�vb&���bCS�1%oH�!BD��Ӂ�#A�-.�(��Q���E[�9�?�i@��2z�}?��@{C��6���Ѓ�6ǀ���y(a!HA�bk��ƈs�����Ԩi�*�R���\��ª�ƙ�#���ɡk���K>w��gw\v�9��j��W�x����7�������O߹wە�U�6����3M"IK6��^���hc���=�Uy�A������*rTZB`RMcU��*�`��o<�O8��%{��^�����������γ���G&��I��CFTK�ɢ9Xd-ƄOLc�e���2?L0��ϩ����=h �H��j-�P�T�M7�EU��E d`v�H����r�A�[=��x��p �� ���4u�jت�b�l
�pa�қ����
+�|��v�j�g�Q��y������^�!�\�.�;��r寊��	��?K�'o�hz�D�[Z7BNBK��������S.]�/�5M�>��)�Q���}�#����=?<�I��=đ�E1�hj��o5rd�x���o<���;W�(�q��_�!\����Z�p��ݱ-\pچ��J�^�7��p��#�S�F+��څ��g5G�f�^���A���w�X[x�h)LDd��l��غ�#���Ĝ�fmKh^��å}��d	a�F�O�{��Úֲ��n	o矉u��9�{�bx���+��u_h���)W�⎳r�����Ӟ���<Ӵ&�r2���uN�K�s��yW(]%݇2�i!����רΕ����CaŦ5�}o}ChR�>�@���p������a�u�	�^���7�!�s������GՒcm�R] �^�ꗨ��y�O��Ca�ڻ��٤4n�kjL� 9!_!@sF�����`�I �}h�56�,%c,)��K0�*(��ΨH`��ܻ�Sn��s5�T�.��W�iVɊ�4}b+��dJ�A2���Ђ�����ssT*�E�-�+A��K�ä���d�lލ ͮ���vRT���2�f2���:JC�ź⏰}��<�������t^��h=�ةJBj���P�6�?�v|a������v~�U/~�?�����`���u�����#���S�zǵ7������W��h�|�-@+�r�K�Jg���DN�>����B[ ���qs��b��)Lq�*��F���wΖ=�[�p��PNy�i�&?���^�����_Zװ^���5�N�e�K�-H,Ld���n9�](,p�U��C��ve�ŀ�;`�'<B�2(~���"�P�|�˜��`9v��G>��9��O1c�5���O�\�:͋,�.[4�BH�L:1i��'禦�hg��R8��&��Ii3�شY᫆�Û�rL�r�ii�� "�ٰ�4���fhZ;��=�B���%DĈ�gX�R9���_?��bk�@�-�0+A���m��a�G�Z�,�v������?+���M��кБ^a�����ó�����B��~��jG��w^>���T�G�f��?��й�@����
e5�z4��*�������+_	{o�!|���~���7��]a�ڍ��mM�PhQ zv��E�VC$_, �c,�V��B�����g�|�\}G����n�>��+_��/ޯ��2��,���3����?{G�O��^���
{��1`R&�̊u��WVK]cآjҽ݃�O�����fU��6/��������uo�sc�fH>��&��pX�U03T�T���H��W���rI���g�^�����w�W���I�t(��Ya8��"]oB]2:���V6oj�X�j��@����Ⱦ�&Ҥ�Y�M���#q��-�䖨@v�\�	���l��704h�J4?a��q	ݩ9T$FnRmHJ�a7;�J�G�
<jnQ��Q�7��A����S�1m�B�ZS��u�QE�z�}U)HE	��u��!�R�B���e �A�?�@#��A5%��U��R�r+H�͖aR�Չ�!����r�K� ��ځ�/��/��<���m������877!�^}���s��}۾��?�����W��P�M�{��+��u���_�F��z�LmE啥��zq>�\�j��@�h�z�:)�Y0��e���8��R1�.�׈�i�3G7l�r륗�G���z�c/���?��������u��P�ش:�4�r��Ce�^���T�5jk�CK��(؊d�%"4����x�hPh�rJ�؉l��C��y�9L��(������8�]������d1��Rp�5�MƋ�[�U)@��QW'7�jv(ح�e҆)������r2�^���4_xv���1|�s_
��5-mZ����~�V���C�Eg����Ec@�Hv�@�R�9��d;��ü�j�N��fF���i�bYښ�;��D@��h/.U��ȑ��O^��v5�<+\{��f�"��Ғ�>��S�WJ[���I�&&��k��?5%��]�+��T)YBmX�a�|V06�H��ck��a+|é5*xX"',�	�'����c.`����]�#1C�}��-E!�߽K镵���RS�4O��ϐ�'V�t�Y/�K��"8��S���@'�R���v�]�t15n����v����F8c��p� ]�J�ֈ��߹��T���������7���sT�5�?��7Æ5��%/}Q8����WL���px�!��t?ý�]W�.���S4@pB C�X) 6Ť�+�f��5]��U �u���,$jb�N��`d{�����������������	-��հB-?��j_x�c��s~��7��$گ��y�L?��o�Z�4�:������e�O��X����Wÿ}�;��M��J��:�ڀ8Q���ރ0�<Idt����:) co+H����R���=�&�R���x|�a���!CO�C�V�-ٚa��jp;7>|d�}7��ן�/K@i)Y�Z7u�w������~���i�RQg���峉cSS\4��ʰ����z�X ��%�Xq1ץ�5�%T_�ҎQm��W�Yu`Yk��{ʏ�7U�}�_���o���TQV(�)�<��11���G1�^��91��a�J/4z���!=X?ö�H{u^���([�f���\�cD7�H_����lV��W���#s��}�b��!}OE��(ѝ�BI ��_֗�����FJ-� �5,��Mq���}�I�AS�d@!���u�y�I��Y�Il����%�zZq��n�M� ��S�� ��E��0�.�Nm8��aSb�p*M �V��febV�D�pX;2��VP�D_��T��	���� �`Ũ�\����e:����B���H�oQ-�Q�
��+h+ֲ��M�X9s��,lC�i;�h��; �c��E�d"L��I2�>_5a�}/1.x29D��*�?e�����~�]n��Z���?��M1�%��mo���4f��*�z�����Z�P�դ��
�'i�z�=���}���&�J�2��N�uP��uj�Ю�k�u�Pxޯ>9����V�RƔ�A��3�S��x��qr:vk��m�d��jt=:K�M��@�D�d�Uڒ@���(��H�6�g"+B˦����)�<)��WTo����/{�uJKT�l����ܾM�������Nx��_�'K�Q��^��g��3GGC������hoy�o�']~a8���孍�O�������*,[���Ԍi�'toT����jn[Ɯ�uϱ��^�\�MKD;���<E�����+UpN�:�ȴ�_�Y����P��H-;�$P��Ա}����e�7^��������	�4��l;�w���|}wg�	�וh@�z\戴iM��ދ��tCsC��ʯG�2Z�PKkR�Ƿ0�o&� M��TZ<�m~Nu��5#���t�LU5.� <Q��=�-:D|��ҮN�4&����,	��D�������UY��.O
9���M5"��Z[$��ϧ�M)�FF������a�i�3�@|Y��ź�������:/���*1?v��~c��-&�,���c��Bנ�'�)�R�n\Up�
�Y��@yJ��
iy�%P%��J�E�[Wj2ߨ�LM�&�AT�nN��*9��/�<������β�.P���~�$�8{U���������:E��:z�'\t�i��xr���?�.���]7�RCQe")ck@,@��#껥�Sa��}aBmZOo
=�#�y��VZsuX�j�	iv(<�b�����!�0ƢT�kt����͊�������0pxO�~O�j��+p�c�3�x}��KU"�����sW]$2�&n���oSH�����o�|�+_����1��*e�U��BgBJ�D�N��
��ѥ��-ר�K��\�
~LvV=�9k�Fh�E��9፯xv(��K_�O�lԉ��5�ۤ{W����zj���=�r ���<)��T%cx9��N`uN�ŀ�u�91�cbR���y���۸Vۙ 0�*�N�P��(ܥ��9)���~�������d�}��Xs�"<�O�G;��V�ii g��p-/RE,U��e����j�Eg�_��p�~'���.�������/}~��u�B�X��7u���a��A�c�&�ia��,���,]�&���5��� ^܊��w�	qK�}Z�i�&�زT�Hr��@0h5U�Q�9~��_���Z��33~��Yk�>��������ǏN��Ըk�@aXm&um�V.?��+.:��Z�i��e���8�J#(U�E�]ԸjXXk	=�!��]��c�V�]�lY���љr�j��C���8$j
Y�eb���0:z�0�ؙ��E���%�U#g�y�f��v�Ľ�j�PbV
u��3�@
k��=�x��2Y6��f��˳P]�t�����ؖi���b}RA'_�-��E��m^��b *-OKS2��p\N����XTH�J���P�Be�P`pF5Z&�f�Ճ���s�*9�������.����W�vز�p��'�[�.\q�����P+��yn��I�R-�9��Ë^��p�Ĺ4�,x��g>��Y!���J��]L�\/����u�>d!��=����+����S�|�z2u�.v�j�9L���fi�:�W������<=��տ�ᣟEu�T�*�}9��B�2sEL��g��۴L�������F�Gì�R[����/�M��� �&����Z��OSGt�G�~�O�nTO29ezDU�v�W׹=��c��5k��K?�9O�T}��U��oڨ"��l:<�O]~I��ݲߐ�q�T� Z"�u֨��a�lQ;	F���U���O����7�Is}<��^����	�x�3��V�Ԥu��c�X;'�w�Yᆛn4�UӠZ:�}TF�Buu���I�D��i���U#���c�i��<&;6r8[�,��hH8���j��>$�3�;���/c������"����(|�k���P֊����@�\
�JCF����>��de:mE�Q���d��^ce�V-%�@f>Br�� ����db		��7�m��&�|N��"��֍91S0@V�ܞcv;�A�n]dU�았c��2sMdYJI֖�p���G/:s�w�ҋ=���c.;��w~���޽��%�EEm4��� ��fKssg}]Aij��H�@AKq��:�׆ʦ�*k�gkj�TA��/�^__=��ֺ�P�a:V9|���+�zm��� ��r_��:�	J��I;i����fd^Y�j��H��qzIb�x2��-zY8 ���\L�1L��"ĂZX/�q��9i,���߳xG�X� ��¥6L��3Rd��RS�0D�e�z�����/�~�^1
5U�{���a���hWh@�jU�E���\EMK�~������-��ȩ�y�
��1_�}�=�{w�{�_�W�.�<<�����G���uk%�}ax���rd�O������?�����������i��i���֨�29���%�	�� �t�}��36�7���w�o�0!�J�ݏ)3��r��ן�k�z�w�R��kTQ m�M�cs���������~�	Լ��oox�)%ۦz���o}�����Mi��¯��s����*�o\6m����o}o���[�*�*}���5/��ҹ%hWqD�ղ�5����#��'�#v+�uŪ��'>�I9e��+<R#v�4R��G�7���p�B<o{���.:;4()�C���}%|�_ ��(��������+@��p�c.�"��fX�b�U�P=�Ç�����û�����������f��w�&Ӕ£z����JV�#Z}�F����ׁC���j�F�11B	�������R��Gm�:�K�\����|�����ד��87\#���g_iMc�}����];Á��l�B�z�+��c����k�K+�*��z���$Q���дl��Fa1<�^�o�.zؘ�獴���@&(��F�'W�¨ .�iJ���H&��f���6��6��
���%�?�v�*��ѳ�I�qb|lv���г��巜���a%������?{Ƕ=�zj
�mi�g~b|�\eH�ͯG�2Z���ӍfbJ[.�?* 6Ewg�?�/d-ZY��4='�ش�m��T��vw�ۍq�А�aZh�u�R��X @I� Z�s�vr���s����i�`vX�-x�ύY%�>�=\P��q��t<�Sd��n�ɝ6?�5�=c%~o���YϺ�B�rk�x���FAԺ�d��@CtM��M�x��_��K8[���(�Bw��51���v�h�CGyRn�!T������{{�����B*^XQg���9	W5�^r�.�,|��__���TO�'�/[.�"��z�5��f�@�ֳΑ�����7��@E�ո����O�2��/��Cuk���g�-|���}�ƥFm�����װҬ��()����f��C�?a��K���/;��� �؃��1�
+��j��榛n�ÁЮ����ub+����w�{��^ۤ�}(|�[����&ց�-b�zU�X B�c۶{�U�4�z�/�N[;������תN�5WY��J�`j��À����WT{K��	��v�����ưf��[K�^�a��Χ;l�z���(V���e�[n�5����^��ɑ�*��ad�/���1<U֟y^��W��z��ޫ_.{Dz9Mx�<����QG�X��	w�)�TL�OM�A��A[�A�Rޟ�7�ĳ+?�,,�9�~����\�r;�3��_$|�o	�y�;�Y�~t���[��Q6؜�	��7����>�#ij���G�}����\����*��y_�k������� �Z�*����Z*�@;ڕ��xf�g}�.R���H� �����Ș/��� �_�|��A�H��^�O�o���Os�z�����g�����i텖����usϷ����#`�($������=(�7�i� h�#^_Y6�P]=֧�j�4����?;6��C4�B��K`�|dx����a�����j�5��,K �̞��)���Śth-T�}�Α�d8�q�\�`� cb`}e�(�u<��[w�R�?�;��$/ X�^��7�C�p�m�*��Oz��X?C�nBl�?�]-�ֳ��S�J�+`��&g	E�-��fw��h�-�L�/-9*��D�U��$Ǒ�_���:
v�����W8�P۴v���[׋��Bp#�1O��TEW�;]Yd�]3����&�+U��5�\�i�P��ມu���u��LZ�~U��g>Y����W]���:.��:��]�*�)LԤ�mZ��� ���kC��c�����H h(	4 �%�2��q�{��Δ���c��l��F���.�ތ���OA6Y�v��:��ڿ?��O>��9�P�@�r����YL�@�!������8�f;e�0-ب�Ya��Ȝ�T��C�����}Bb�~b���J�g+ugH@\������9��Q�#TӤ��B{:�*��CJ��;��3'�9!���	4�gk�ig���������m�jR�����������ܘ�}��5�	���i.��>�*Ǥ��0��I��'�M����\`K��z�)�b"h�2.�U�bm����b�fҥ�{���~�b{���5�ݰ�ĭ�Y��|�[
�Մ���{�%gn�����}�>e�	$��	�o:csht�
�\mz
'��5F3��ఴ@�J��Hi�8BN�a�_�!a_�"��6ր��=v|��+�'B�V�Й^��jc3�(V�.Ku�`KƫѵL�ό�jm�XV���"Pnjh����?:��hlvV�
���R"�o��U�w���89�#�j��/�2Z��{�����]�����OL��JX"fw��>�ǎuu������*�7B��19��ʡ��f%r��j��,
���*U�&������B��y����|�Co���K���Vq���L�$�0k�
�-�u݇W��wa2�����r��?^�� �|wy@�tG4t�b�u\�����3�SU��2`9:w�����Mz9��)P����b9�֊P�{FbVB��Q��ڵk����b��u�	��Q����я	�VA�M�k�-�	��7�7ܭ�����7�R�z5-j�9-�M�&^���_�e�!Ԫ���Aiu����0�~i?2)@7��u�)lԶA�a��l=���2S��{z-�R�h���S�mB�U�]��B= ���IP�]&��q���A�]��E��� p�a�:����B741%ӬG"�Ze�+���5b��S�eU�VH7T+�U�̪�e�Y�������F]v�槴�5T�h�
�]r�a��X�\v��Om����@Wݭ���-��ebT�x 
�~d(��e�~�A�"x0?��Ig���-m��B�5�},��W����!�z���[nW�_}x�^~빏����^��pݏo��f�AuuJ�Ƶ�ĭ��Wx�߿6|�K熧]����k���G��_c����pDU�ר��<������0����0���b�0C44�`:�ɂ���d���'2�_f�4�b���9�$���ª�MP�G���*+����Rgmъb�j-��*��..���d�b=Uך�����q���;���?_� h��1�4������̩u3�h��f�;g�O�`�4��%����������-k�X�)pg�yZ_�p��5|R�Ҥ���#���"���3I��=�~��,�'���v1�J:��?�Z#'��������I/�O6�e�&�FJ;M��=��`�F0�X"w�)��	 �杄	[_D�����|X��!��<�rR���c�G ��bu(�V.&�pwo���l}��tPՋ��qf觞���5ᴆ�IZ�T���%�ՙ���������Ђq,�c?,��m��L���c
����*^8"�  @��ƃ"��_,!D�Ǜʌ�9�^����ɏ�����r��-�s��A��cM�����l�J/�I�\Lsa���9$D:&@j"~9�r�O?�YӤ���@)IP&��/a���u���7�.���ŧ�'���4/�J� [��L���8�#��dr�r0 ��T�����b�?�"�m���T'�m���Z���+Tʡ)|熛��2�KNZ���*���r����½;�)��U�\�	��R��w���6�����m�����Vv�&1�0Q ��U��s��	6&����#,)��n�$�oP~�!�O��7��jZW�=�m�NC�R=�|�aD�Ҳ͔V��A����!�z:�yŒ=�*BMq
5%��in(����B���,�A�M=>;W������kZ�������C��8;3�y��ܾ�ˊz�x�>��xO���O�v�UujJ���!&����`!'[,^Ls&hx������S�=M�T��ɿ[����N�����µ�x�RRi�V'I�9+�e�͌=�E��3��F
���Gl1�p' ��8������c�135M�LYO�	�=hƨ�;*q0L�+�[[�=9Us&if�>�H4TXq����F)�sb>*q,mT�8%�M㚀��Z��ċ"r�`�y'�{aX�JoCe컶�-�3�j�
� tt߈��F+��a_B�T}!�����k&gJ���՘7ԥ����Ұ�`}�K_R��!�[e��{���+V�2�5OX�"L��]*�^��XE]~J΍끅�0�gO�J���{kT'��#��^�����C���7@�N�k��Z�cǔq'mz)��FCECU���Y�~���4mj���e�m��}Ki�-a�g ��;Ø�$���y����6��������-�F����Z���wu��I[5��,7
r��o�jV۫4���	���H�5�����Zs��\�7_��,n�E��L��m�aЫ�F@�Q��x��lC����y�٠c=}�Uu%��UE���T�@��U�$�O?��p,����� h��FNB��Ւ)��sF���]yþ�g_�o����羽�TJʟ�u�ۗ����D�Ji��/�~�ŗ�g��O����S/8E���I;���D�H{عO���N~�I���JN�����{9ձy�-�ѩP��0z}c�B�\�'����Y5�S\{Z��w�Ƨ��O,-�M�9�� Jhd(#�D� �D�-䆎I�!����U6�K�ȸu�:oڪ�̣c�ڦT�FO��Ƌ]:@�m �z-�e)����z���CZ��/��ԣf
p�3�c�G�"����f/@�gU��
/�*n�h7�K��JúH��c�Qա�\Sbp VU
CK�V�l2����8��a�� 3�E�sF�� ��S�j��_St��(5���EF�!��Zi�Д���j�s\�ڦ~��견�e�9�"��T�Iu��yƔv^By�$BX��c���kv�p�A��O'3�ㄝե~�y��b�1�_�6T�,7 ��$z��n�i���l�O�~e�U�5�Q�a�ƇB�ŲM����^���	��1/��Q��^,��� o����7|s�QN_O~��F����c�R�Ê&�����ޡ1��{y���utb��S_�޲���ͭ�i
�������U��|����t�0?X$�������+2��j�Wh1�~Ȅ�9���xު��g�d���_qW����v���y��5]���+˦�"쾽����%�"��؍��8EQ������ ����-��z��!�Ŕ�)��@wF�A��94�{KXQ�;�d��|�4���D��X�v�iG뇏 r��Oz2[�:��5.�����c�|o�MD-��-���� �S�@A��I~�u+.@Ct:%%ʞ�f\�WZhKT�b��nl����6�6��BK�r2���8�H8B>˸9rD=�v�:1M�UDGp�b�h��`�UPś{�5,d�����(�g�ki.�P��:T��>[� F*���%P�U�RU����(@���g(�c���|�ۤ�V1���C�C-,X���je��@H{%��q����' կ^Z��ej)�>�ܰY��2���J�6*D�^�T�A���r+�i�<[��T��
f$@m!��ܙ�J�����d�J(iA����տO_G����&��2�(���B5�J5��B��b���T��A��zp���ҿHMdQeD�ٰʘhr���fƟ֕A�+�ܘS�������σE���_Z7��
@�,��3YI )�*�ٹ�ؿ-��F����i�w��G�O�+������+!N�-�A�k���#�-q��r��xV��5<�����X�W�����?�_}��A�AK~]s��o�뾗�T�n*��.�⏓4-�8��R[N6�"Rж�Y2�RKo���=��uq+�T15>\̈$�b��Fqg7��pqX+��	h��%��x�@N;2��]C{X��E�� ����ig`�b�0�\�#7*��J�5?.,̮�Y|��}\/� �[rZ�C>�צ�p�t�^���ߌC*^�
F�B����� X!�kTA�2�H��:pM�ƪ9[m}�R�@�tw2�`pRaJ�pd���Q1t�g�3Tn����tn/iOĖ�M|�Z�H��s<�u�b�J�6��� ��8~��p<g�$p����i��븴1@�C1D�
� )�<o��V�a6�}E��;��V���YZ�G��5.Qp��r�J��r0zV�*+�3)��E�_'���
A���F5���J��lJ����?��Q+e�����r���!��l1^�emK��2��:�J-0��>�k�R6yo�C��R�q��&�gzt����W�a����xhs6!�rZ�gT�V$}��q��B�\.�Jy3����\HC�:�3mVb�.=���� �������E������JuU�3ݧ��$�[(�*��M����+����S��Cݶm��C=��O��t+9�X� uX���Ɇ�ꮆB�Úв�?���$��⟓�������DeY�$�4��b5�bv��-a��3��9�������7���]�e�ڻ�\s�ͯ8�?�����eԤAӀob���!ʴ�܂C?yN;�ű�����Ď?��ݹz���!Z6�}�69�t]���y����
5,_�w�:pց�V�-�
]��\Ӕ �|Hm�v]j��;֟�}���Y�'Υ���]k��|8H�
��~v0�},�g��y��hg���iG@9���M�wB�pjF��ӵ���~;yמ �b����n�B�;��tTa�RlK-�*�8�EH�ȗ�V,@B��¿x�Ƅ�V�/�e�8;'GSQ�����2�o�H:�)\F�M�=��<�7����n-,�{F[�Yo0�:!Qv���>I�!0X�z��dz5��U�M�I�Ka.�Dr�֞B܁k͘��;���a,QdM�AHs|�\3���X,,�Wu�|-�.S;�+f2Y�7����;e�%�MFk�ߌ��|�ar=_��B�+��T�̘=Ӎ�c,��`���){�o���F�0h鹧����ʶ�zN۹������=������{�145�Ue�L�%@�Ҩ�ǌ���������r��zY k��8حu���E3ݣE��M3څV�V��בɀJ��[ղa�����򚳮��ES]�����_���_��\�����K��x��׮PCL�+��gFxh~��>1y�b��>'�P'�5�o���'̲(�~���Y[f����CA'����̼��y^W��b���{4��k�`,�1U�D� �	 �uk��t��g!�>]�O��"0IvJ��9���^i�.FE�LG���X̒�p*骑Up~�0��'�K�!ZoDw�?�N��M/�e�gEd ��S[l�yh׶p��lҌY�Z��b�B�@��V#��j�n[;増�� :���.lLX}'}���(7�V�3���^�Z3{1�gi���EGz�v�@� ô�ƗIS5)V�O�g���x!'��<��&�h�QUSzLN�z�Emw��	�`��h�Q��a�k�u�����J����y�9�����|�,}:eFZF �$��6�`1���,;^6>���2��g(6�5���1d-<sșw\[�>��X՟��q��8�L��æ�ã�&�/.)k��~��;���3�n�rP~�ׁљ��~��'޳�೫�V��S�ƼBe�T@�ácG�7/�o�M�3\z����2Z������X��G���ytY��9��,�J�],]�K�J�^|���g�5U���������M��SG�u�����54�M55��ssǏw�t�l���笽{�?������w�l@vgM���H���h/,;)��Ӓ{�4go��W�����ŋvJ�~(L�bg��XŬ���s<�hXp�񓛵�t��Y��9�3ӑD���ȼ������o�-Td�X����T,E�8N��� �A�t�'j~ _�1�/c�����7{*�Y��Tw�.���5���޿�� Qr�&D��*�}�0^z�J��UV���5c�5�k�� �]+���X'�������?k M�VvarıכP��Ҳ����R�{
eΉ���9����P ���P��k?Q~�F���ʂ�E��ήcV!��vu�`y�4:z��A/Ay0N{�c���I{����%���Wl� �;$�n�FJ��r�%���TBB�SXbY�X��DB:�$����}~ߞO�aΙ3sf�+E�D.����^U���b�h0j�E�K}�H�dW~��Dz)� V��&�W�i�%W���D	X�����8�j'����n5Or���W��em=�l��#HD�����`��Z§�)cs����L4Ϳ�>�33zݝ�F�z�?z��^q��'��YX9��~�<�+���g��+����g-�7�?n5�յj���ZV�z���&4n	(e�.�/f46�P���;������:Z+�`�O��}���5j�a��͍���8��c�,)����=����yj��2Z�6�٫��	�S,�I��N#�`���?�Cc�k޷���c
��%5�?�)#Qy6�y%��1��ʼ��+�]�|hE���s��07r̀�v:��v�Z��Y�~M�{c�X����Q%�}��T��o�$rrs�L#"�<B�49Y[Sa�[a�J{�̾��tܖ?j�B�����v��w�4WLb���-B�ؠ��Z���8[B��7�+�W)y�O♇vE�?=x��u�SQ���wLS�����ڥ|��kK��C25���1��V�x�}$�>>��&�Y��� ���>%�t�䩪�����Bz���W?/�.U7c5�y�ꁶ����^*�Ӱ ��'�R��8%�ت`D�A4�c���jQ W)�l6V���O�=|J3mbH��J������n��}U<>����y�W��)����6�2ʃ'���K�d�'��y��y�iH��-�J�e�^K���DK���[��v����m�mAJ�jb�\����Wb�_*z�8/�/:#�C��J�>f����e��"Ҿ��4LKy��?��i���I���l�9!�q��u/�g�}����x�7�I&����w�KKjƟɴ�A��_�Ǒd?-B��BT�W�0�b�s���\=S���2dh��"�?c�ޓ���w�Ŋ�u�7k��1>�+�=�0�w�x)�g~`��Ӊ^3h@ ��#�­C(ͭN����E����p@�V�҂/�����d%�|x���Qՠ;�M��V���ff���1Nǆϐ	��L��mEѮ�}�#����s2�񿞲���X8����h�"*l��UcݽN�T~���ZwدS�柤H+���4<�4ܶ%xG�V�ݙ�9k���>�0ҙ�\���B�pS8?��3Vh��*�G&,iL���C��!��Ɉªҙ�|H���K���t�74���*�b�{2��$�&��e����[ǳ�1G�8ô9�� ϔ0F���]9��q"l��ʍ�mZ��ԥ�ta��C��3��1r����*T�Ÿ�T��3��ۮW�q�Ue��J*@�L��u@a���?�?�/�rj���y����i{>�/ڮ���q~_۠�'b칀|�-��:��v��-&��ۂ�-�'��R�4U�u�U�Y�݈�SАbI2m.��)~B3~��̰v��f~���0}��in3l��C8^�Ig����j ��
���`���7x�d��&NHdR9p��C}J'<U��4�_�O�ŴO�)����"���y�4j�P���3B="�;^�����Z}��-�г���t9�j*�@6P5$�lkrx ��e0ԡe�v0���.ݶ.��8}�&�>�k(�~u�03�=��h����e>w�����_�������L�>�8�q������k�F�G�]je/w�u���W��:����]�S�>�:�;��՝L�^\�m��'�"��E��c��Ɋ�D����UH�h���k��FGKw����$8w0޷� K��n�f���wR�*����!���M�\��o��Y�+y�=C���}����l<g�F�p2"�k )s(���ɠ'��?G����I6��O�7��*֠�3�bo����rJm����@kr ��M�-���9����jW�`��āT����.�d��UD ���Ф*�_�uW���9�3����ΒP����4�%���/7Љ���Zܤ.��C�Wk�[����TC|˥���:�6�њc�͍]����u#\c�$,��ت_�ϸ��r�����;���*������ ���cs�U�[Y1%oO1�4�� U�5n�6΄A ���Q�^�f����;U4)�y݁�\@#c�B�8�z$�H���:F6BX����#3]�/�m�A����Z{�M~j¥�|g7�߼�qqfC`[N6��}]�f_��}�$��g�\Q��n�T�d	9����&�����6z�b�V�_l���fJ���E	��ӑ9d����l���M�s�;�|���9���MY;4�-]Uo|��t���@���<��ĭr�op-�_4���1����-�ű1P
�5 ��(�\�j�W�n�>��������ۅ�eJ���2�����[cg�_��
�L^n?<�xY���� ���{�ۍb�k .�>MZ�����\:]��z:�X�%�B~fwX�
:\6���M~���m��H�������suC2j!�����`������vf�6��+��b�ū�=%J�ˑ�2DDR�����|5�㸐^Y|x��VܟL���~�&/�ˋi�����@� گ�{����K�
Vh��bDG��Ƥ�<�H��%G<*:i�Ax�0L�K��̊��_����x59�������N�?1�Z��1�$��M���{�P�x���E����RGJ��;����*{�M��lh,�ᙅA����`��)����c���1lD9q�'�+1F)�Lou$|Ø�	(s�N.�_���,�v������oh�MPT_�W
C� �oUǭ�k�Jڤ翵�ɾ�ƫ!���F��G���Dsهsc��J��Ĭ�F�!֫�L��?��Xvw�z��d�$2J�s�#4�Mc�˸g���H1�����=U��|���Ϩ�g��g��]f��=����5�!�f�FD��"M��&��_�������)�E��%��G�RO^���7p}ǽ���*���w�A���\ķr��G�Z�u�<kz3@�TjS�<�K��}�Zj��v��^�2H�Y�"٪hg��n�|�&I��^�OF������$dd���,S(q�W�f0�f����Ӗ���U����9�6Iw4vW>`�c*J�f_�g��{&��t_���]z��q���|����/��Fv�٘�r�v��9�ڄ��S8��-����y�*VV�+��f�6ᕮ��M�l��	JB�t,|Et,��Lu���$�&�}-�r��M��6 P=�G�ԏ��X]��^U��	��c�+�C!P�r��Zs�ċ!��̫ -�9�}��-�m�[�PT:cM�z��UnV%��Vs�j\$06��V�M��}��Ķ%��!�5������<
��K	�c7t������������̤�ͫ(����''�T� _P����\Ca��Y�,N�*jU�L4{��Du�Yw�'����|y�o;�`�?�,,��_ʌ�RHWb�',���֢g��=����2������34���p��'�s����F��²�'>y�ա��f�7���,.��B�����0�]�zM@��It�w�iM�u�l2ι۹����WM{H�S��Ÿɹ"��[0-׊7;}�9*|q
��y����	�|����ͤ,41��P~��z���il_�њ?u�Q���ף�9��5׼' �%p1�\��`t�����%�W���D����H���Vs#���2����dJ]���޸j{6�Y֟�ӱ�38�N�J�,�$���٩5���q5�������5 9d�I�Z~A}�m�<7v^=&���F�f-���(kMuS�O��>�yW�Eb�i��ix��W��kL�*�$`�x�ko����V��㴑����l�J�"
�X�����9B�����{o��;���b�m0��s16���+5[K��r��]�0�Y�/h,����I�q�H��-[5l_iQ;C5�����2��o/�_	`>�'o;e���|k KX����[KiB%�/���V^qX>O@.W���A~"�x� �k�4"]����N�$\������Y���<;f���^)�vh?�OΙ�0�((�O����&���*�H�=��Nw�}F�_��%���İJ�,��шw۬|3���g.�/g`9(��&&���sB��OK�q��G�k�U$A�-����ь��X�Ix�V=�cNq!���� /���gt���E0���]Ll�k���AO �R&'MyvG�Y��������ӅnR:97�o:�\�+7J�d����.���������%ϩ���sf�ԗ/��Ņ]����>I%N5z;�p��g�^#�"����dl4�C�2���[]6?Ȑ�/M"��;���!����ǉ�']hK-&@��d�V�Zt��x_K\��lΊ�%��'��m���o���8�K%��<���]���O΃��O�ϯa:�Dr����О�� ��3.�u��R��}j���	t
��^�gSD���||����c�Pi ��-E������MDF������)#Щ��'��e�ֻ3E�K�o{~� 敜TU��]�?����&<��1��g����NW%<g5��.4J��rx eX��pB̮�cl,{2j�}�6��q�b�'��n�a��� �Hc��� ��"y��>I�(�=4,i����>�>��;�&^��B�I�]����IKt �:B-�b�Q�F�@�\�Nm^�3�2�v�\��ⲵ�r�bY��L���"Ĉbc��1���a�0�J�iP��[��Y52q��
"	~��F�1fNk��v~lI�)Vc���^�~G�����3�*ԝ���&B��3���O��}��-�����"W���Ե��Sxc�d�X��X?J�my[������L���@,�_�V����QZ�Ca�n<�EM�A���1�p�k�f��� {�h*/uٲ-���v�����Y�㷫�	���ʟ������J)�s(�v1��1�8��}G�7�cs<ǎW���u4����9CC��ᓷFji��$�i	D^T�o�mx�}��٦7�-���99#�ΤN��z5�Y�D����4�E~�F�獓S������۩�#F
��.��;v�:ԓW=H7��Yç�Z���|�l���4�l�a;2���m3��tcɗ 5��I��HHE(S���eγY���Z����ji��RV�m�ZezY\��k$� �];�#z-����!!%���_���<��g4=U���<���E����;�D+F-~[��t4��u�b�0\��amַ̀���tS�2TJ�U�uehٵ�(�Kj�J'g�vlQ�}]��U�#��x��N��d,��G>�y̡(��㰞p ��4���!�2��AA������(kp2��	���ک�е�
�X��F�6Ū�_"M�
�91!�h�)�Q�hb��ph��6 !!~�Go�i��p�/�@����>�A�n�=�u:�8��pK�0W�4�n�K����q`e	wW�;��?ET�c���q���6��a,d�.CZq�/tX� ��ϼ�%J������O�Kͷ��/�Wx] j��,�MUjB���ZtV� �SLo o��11�P����fO�D6���h�i�3�b��I'	f'f���ct���������R�������N��6/O\\<nI<q����&�Xh%G�グ��z7ҁYyS<���hbcE�jû�[)i�ގ�+tusc��4	

j�+�GP��@x��a��|��eֆ)Х[oS�k~��;0j?�T�c��iy�u����xe;{��j?Z���B�-='�ɟ�!󷓯�\��ke�
er�������:յ�ňm���p� �0���i�#ڱ6��6qO�����(�X�5���C{	�n��)V���A+�Wɛ6��!D�)�u)��Y�E��/�	҉)�������a2������V�Id���5zvV:�c�.��ݵ���@��27����XK�&$m���_��/�Z�����?����[����,sN�ti�J%�OSUO�^���� PK   ]��W�a[}�  #�  /   images/d19d5e4e-12a2-4f6e-be69-d40783d16976.pngļ�WU�6JJ�4HJ���HwwIKw(!���-� �)-���͝������Zg���3�xbf���bo�񑡠��H�+BA��BAAg#�?��pOޠ������AA�@I(;��#(cM��tB�c�c]��O���(`}�F$Rg�I���@WV�~�)[Ǯ�4	Kn���g�E��M���㼶��⡴�U��ɋ���Ht'.?�8	4�\-��ү�����JO���CRp�_��0F��Gġ��u`�篾C!�&�����O eUvY��u����z1�Y}��O�@c�:����zQ�|(�
l�>A�Յ\�?7F�7�"�?������?�M@̪�G�H��Y Ӷ����v`���y������g���p_ɼ�B(�L_��,@p���ηL�ġ'ϛo���)k���O ����l�'NhPz~���o��搩���TU�g�#ɏS�74|�_�KKZFo%efV�kii���(������e&�?�=3�ӗ������u���&�B�}����h�9�LD���2oI�����wX���L�*��2��) ]*2�V��h^�"���%�Wj*�=.#C���Z��`��i~~^��Ǐ����&��3C��cҲ����}ظ�%�XX��hhhb_BCC�A^�R���'&&^�hiia�%UU뾂?��::�p*U!!�))�J��������"�zkѣ���S��,555{/ccc�


۶��DEE	�dqsk1�����g!پY/ϢB��S��{����NL��7��x�����z\������j���j�ⷀ�d��̏��))�щ����0�Hd�F:��	�n����$�4���t�4�����Tq�˵�p��|_��8�*����5$"J?YXX૩���{��� �CE^�lr�v��s��v�0rz,(�(P5���U���0ggg� 񢙼�̏�{J�II�&u�X��4�{�Jb�(��	'
c�#KX3!��-�$D9az�D5c��H��e
�̤�-s�3 ���7M�D�L?Itjl�|jJ��ӧ 6v�g}c����_�ޝj���'MMM�>�"(����A]N|.���������I��ʺ�:���p����b���_:JJP���+}BQ���Z�)�$��h��N�Y�)׿`F��B��O���Ò���+T0��Ezp��BB�|T�\��� %�GӬ1=kS)Q����0��𜙜�*�m畦~�x��7�D��p̠�z{
;q(���UUQ1�3�}J��E���͉�����!(�?���F�ܞ��||��k5jLїA��ˤ��31[/5�����bs�3��*��h��кE��hk2P1��rr�[�κ6:}����S<�/����E�)�_F���������.P�&���ೊ3��LON���۬>��rx���u�;6�	U����	����;T��A��Ϗ�'݁��������x?��\�ȍll��'m��&#�d'��K�N��M&�����|��m�M��]_Yٰ�#N���G
gMA+Gp���,!�}����)}���f������'+��� -�]\�`�R�)le����>�3lU�d2�L�H+re�K�Y.�R\\�����v2U4�bgw����n ��w^,�52�7$S+I��iP,�4������ғ����aa�w�{��O����(���y-��:�U����!�Q1���#�Ī���w���6;e\�o̔�ԙO��&$��|~l���?���qg�h��)RM.�N����렐��g�k$$�{���jV��?+��e%!��
���ǐxQ:��
���v~~N	�����~�G���q����jv!�����% ��W"5�p��^C�hDED�V�V��I%�9�fɘ��'o����s�VŬ�)����]�O�����)��uۑ�����!�I;Ǉ�3�$3�;��\�-
J��v�}𓒑S�O`� �,��*I�\�gee�@���7-�7Eu?L ��y��h�KF/9���3�t�%@/f"qV6%����Ie��m2j:��RO}:W"֩���w4h���кh~l��6כ�U��.�N����X����}�}���bDUA9��j:���;��q.�0�A���ƌA���@��X�0-���L����t��f呋�E�9km��{��ø�����t����?5���7T�����7ew�֍Cq�=Nm�#�a���@9#�2,�¸�yM�2괘���Ϳ��rD}����n_�ɢ��p�B�%uJz�Jֺ����7��`�*/�ȴB��<95U���'���6P)1!z=��d�~~p�`�- ��Bq5Z=_��$$��*^Fuܾ�(a�%hg&�p���"��D�Z�����e��%r�6�̏���j�����jc>�B���kڽ@.������d�J\Jjrtt�B$��?�2]Ld�}'�}��R�މ,�$�Q�o��B��::�|�o����Q��o3���^Er�Sv$Vg7��� ��.�Cܱ3�� �s���uj���A��Ǐ8���A�[t�� 5�*:�p�i���m�xt�Y�P�'��a���=_�������:� �O��U�\s��B���q,$(h�n�� ��czzz��X�~O��@�����ig��j�F� �3Ea�2Scƚ�6k6 ����0".�,@r����4Q�ASX���I�F��(Rss/�ߞm� z���)�|V�*,V�$��K)�y��~@�F^A��)����6�o:_�'��N�� ��a�Y͚ �(�y��������_ ���z{���!Y^C������sP^�[V�e�][���7g�=l���N����*��BD�q1����0�b/)�Qh]��N!(�zBBB���=�����o�����\��y����174�������r�wdD�y��r�򟴘��7i�^)�h�u�/��r��{#A��[b�<o�u�$�V�V9�M�h��q�)	��c��+�
��M��N�<^a�ږ���`GcF�*�� ѯ�$��H��Z�(���o�:6��U����5U�'����s��8w��e���藛oզT���)}�I��
���?�1�5�uF=�t1�$���.�L�G�lF@ꪪ�&�&P���޿T����D� ��0�ј~���ڿ��pP˟� <ׁ�����8��s��N2w�[��~�Fν���A�SK]}^�_�lF;pYe s0���0 ��wAxx�[�찰׏��Lw]]���u71������1�����u��.dڈKv�ޣ�<^�,��r��7,�,mT. Qv�Բ��z]p'3e��8y�s8QTg�Z�HF~�ы�i��w���NFFZ�n�/r[VZ�S�d�xP)�?Va�
ӳ��U�0,,�O�_�W��Z�edF������ '�0�DuE�W��̲�R���\eE ��hi�ڝ lD���j�*}Di)�¿���~`	��qp�mo���J�Ȩ������d���f�~��"<.k��A�FJKK����hHzBBB�BBC��vq����OTDk�g&6_Ֆ���8#�����5�#�U��ca�͸�'|����!�L��?��P8�x@D����p��J{��hu����"##��@k��yyY�Ѣ�S��J�`�e�Z��0�05�`7[32[�d?��"�����N����b\\܄��23�y������/�6��� H��R��x%u0���8 �0ɣ���/¦Q(o�>{�aJ|p�m�e���{�����q�t�d��y5[(�xrvv{�-��4�b8T�&yf=������g����ǚrrr^�S$7އ�~�4u={Ѥe4	�h�F���J1�J�7)9�w�ࠝ��塴���O�;�ͤ��!2�U��D��v�;E��dv@�4��y�ʊ���^��q�yyf�����%�į�Ĵ��e����YZY�}��r��I�A�d�#
�zqc}�h%�gްJ�?>ʊc���L��*�cJ|��-�2�$U ��b�����LL��b"���j ���w�� m���k����:Ym9 n�^��m����\]C#�EV6f�y>�&���o�F�b��=�R'Z������A,5�Y""��5�蝘0��W�B�z���\�9�X�VqO�*G۝d5��r�d�����H�z��������
DA��a���Mlɀ��M��1����)�������vw��t�F��S��b��h�o�b�!���b��];r�x�ȴ��Y5 �9p�V�_�g�s�( <u<E8�=3ļ]��%�[�<=�$���S�y��S�f���i��8ٗ�A��k�*Ӽ1g���`��_	��mVs�zi@�&��K	���f������8��d;���:%&&eҊ�R��Ӎ�a��&Y(I1&:������̌�9)��M�NfO��g�Eq~B�H}
���P�E�i����2��'2��>�cݡ��nY �	)姠�Kʃ�`T̺���'�����յ���z��m�_��x�j����U��c"CC'�n��cA���/�3��Xo�df
ZF	�����H��sѣз��[�E�BK)#�Xb"A���g�]�Z4������VW��_CPe;b�a�h޺:`=�|�P@�M^�*�~+�g���(�d��� �͇\a�`������7�<.S���y,��� �0��̈́{f� V�����ۙ�1Р0��IU����)]�=� ��ޓ_���1h5|2��	�Yn��-O��d�BN&���)ל��%3���!����<�w�%��`����s����(qJR�[�YC�󘰠����[����(�r���zz���t�1!j�U.�/�s�W�+>(+(D�9r�ܦ���My�C�A<�	$����$�#�=_����Vkk�rll�UR��
���Gtc�$��1�<ҁ�"���
��V���ށ -=T�o|&����$��BE��<2P?&��R�8==��|���i{;����&ۣIN�oBrr�����'5f��{{�j���b0��Oj"�"��v@�5�kԚ������=�d��6�]u�������VT�<��H
��(&DP�(�cܽ�?�E >�	�?�VY	�DA\������ai�k���m�/9��Q�)���$�/�cY��G4��N׸�m�G�ab����"I��b�aϮw�Y��8��Fj������::��*٤|�n��|�����b����b����oG�.�d��i��"^��6�@�2 bP�$���/Y�,��,b�gJ��U8��r�t���b&�e����
�7!�kғ<v�U�H�v�-.�~75-���Nf��4�x�L���C��x͍���L�Lj�P�[&���!***���[F�at�A�	�r~~���U�|�%aq�~��3���4=��h���C����<�������l�)�x���cHK��O�FCu /��]�a�yZ������`���L��Y-�᳙+W����TR�d�йҊ�$�k% 0n��$MP��ܮץ*�4ZJ$-�Aٸ�cW3��:�?$�����}�i�O��6���><v�G�;`��,�{��Cq?F���ڇ -� �D�ӯODk*�XpXw�~u{N�>�5���������o�e�D>��,nȐ@V$ �m7�
j�a4��jW�J�5�QFy�e�-f˅��-\��t|��!P�m����n�ā�E�b�(�c����qaaa��^�<��7{��E�t��)�T˦�}��3��R�d����`�^�>��2����|���V������E7����&-!��∏�:X�)���ee��������F��I4�S�| O����)���] Am�b�adll</�H����91��̶mO"��&U���Ƨ䃏�����;���N�J�źȳ��_d��@�����E`��&�����,�v����2�[9j���}�+(��=m��i����Qa��CV�®Ed�$?j5;��l���:���
�Q���s�(Gj=�J.,�ˋg������V���a�q{_�J^�GDA'����\
� 5l3�_�wNNY/��٭���g�<Y}�/t�u��*���R��A��'33st�����<��b�@7+ɀ���F��=�O�F�Ǳ�Y���Yx.���z�v6���ŀ#; ���=���/w;7Gi�}�-�.��D$^��H��Ӛ�N��L��Y׆�o1]#3�Z����s��3e֚��ڢ�"Y21�=��Zs����~Ҫ�	���R���.7���A�X����ŀ,���X����?͋ka�=cu��k}Y*���T"�6��L���7��.va a>RGEEɯY�ef�^��~c-�1�����U��@�п-eee�@��`|yg���xx��v�# �\hH�=d�!#�$�!�;-#`U�Jw�Dú��*���0��)F����ȴE�S�wwwE�l�����j[Ƽ;^�@V`�Ɣ<]�V7ʧ���Ib2�x��G���d	��Huz}��
4X
R���H�1��H�v��?�4���JrZayY��.HY"��
�[T$qfPt1�.��Ór�Ù|����?��`�bF)$��`[�5r���������s��i���\�/
°z7�<IAx�J����p��"���Ϊ�0�8ƹ�=[��U���?�w�.*�.�9��1ĥ&������7�bb?FG��`9,�c�{���樅����)� ���ba$^��\��+�����x��:FGmVFR9�'����Kcv��зЌ�RF3�;���Ɠn�U9/|I��5��}�qi�H���&�ՙ�f8��L
Jb�\��8�b���َMOO����q��?�n�	RA���q�B1DHVjx���3�J�Od�S(E��r�	�)�~a0#��3���>�c�{�һJe6� ��N.7}�J�T����k�z`pp;���<����g&��1r*����������.zn�%5x^�S��
1;";�������)���c%>���"09�@O�T�x#�����<=�ˈ�K��F�[��F�_���+K���W�//ח/�U��|�߾E��S�R��T)��V��P�")j���BZ���LN�>����,,���'8UUU���X-!85��0Z�	���#@��{�_$�H����t�����J;����4����J�!Ä�C��y�Φs�\�h�^��^�����ļ4=��#d���������+T�� 2K_��7�
�{����3�=���A���b�Ԕ2яI�_��V���QA�I^����m�k_�����&N���.����Ѿ���BL旔�$�����q��l�LPg"���*K٫������?��B�r� �z	�\��
˰�p c�����,У	����\�Ǚ���i%�f�����uN���`�ʿ?u� a����������V�G��H�����3�@[n]���r���ߵ�<T����hq@N m�	�CԊE�j4خ���u"�@[L�8)�Y�O&�}�3�8����������L;Rم�;$eo�p�ooono�G�ex�K`�5��~�����u[�2�+�%���ԍr<rIqL���,	+��|��"iAH�||�������QU�����N�ԫW�ƐU�߳ �X7l�������A8��y��&�8��7�eTڽ�~s��W�-;$#C'��!P��ذ»0����q������dj*��h����_��Ȕ��W�2dU��_�2�t��d�)�+�PA���l��� 1���ôL�v���+h�w�m������b�� �X�u�F�k���l�����qڝ%2.�c�S���3��b|QUV�s���t��su._� �s �+<��[.��z��!L	N�*��;Վ #�yx
�fO�>�f�3@<������
�v��G�d�h��`K�n�p"���v�{�N2��ٽ����Rۇ�Q�	)����
99�Ȇ��?]�Й?��:�e:=S�'}�j���p̄^w��t��� 7u���/��s����m��Y�OMCU�23%�u���O�,�o��SE���lb���i!=���NA"�Ma �̵L���$�
��?.ᒵ�N��F�����L.�]4z�J"�Sj��{4������|��V���O��}����iI�Q�P�����e	�G'�KK��_;����a8=?:���Z���7���p��$��|0V�\,t���������#�L�~�v����Jhܾ�����pY>|�������9�Z
Z/�թ|��Q�xď�UU�5��]��5�d�c�$�p���K����@R��Mfr*6�=��4�6I)C(X5���]��J�u��C.Jn�2y���Ȗ�V�� J@��4R������4�I��^<��2��4AQ?|0�F��meudY�A�D�[��P�v�/{,�+ǯ|щ��6���nR�^VM�CL>Չ��dW�2pI���GDb��`M+ש�k$3s-�8mCU��~K@���Z ��~���g�����7$���P��GK������ �2�
��f��-IȔ��BSR4�C�iU�Vvľy0�ER��`�|��WR4BBn��F���X�`=�̳�k��o\$k�jF�������S�SeUB�j8����(�h��b'���t�����M��^!@�& 1$�"�Tdy/���*v�27��e���4�
�K�٪���j�d[6��J��1�ߧ�P�g)(��:�ى@��p!��-Δ�گ���/�G�Ȏ��(K���
�{
s�b�!\���=3@! H�dy�!��l.N3:4d�E_���bh��+�����x�o�I)��/F�x�eӛ�ʱ-��26�2�v�$�!M����1�3Ó�^������V3M梢"���47 �Lh�w�y�>�˥]�|��4t����������������"�~�����@���-����2�w0<�'�$vy��h��� �����4΂ 6�utR�L6��䈄& Ĳ��8��\"�`��]�gvL��"��f��,\���q��M�	�	XhW5�Ym`ODӢ1�h�f���z�T���Zg��}�Z��*�{=�خ��K��P��,q�躺�g�����PJ��r�6$$�u��7^"!.�YX��������0�Yn0���2���7������̭K�N�u�x�m
9:�=44��S�6-��D�Y
m_-�����<�$��/��/ ��>�k<~�T�
H����%z:��	P>Q����].��v���� �=�o��=ݼ>�������h#�$T���2hpύ@br��衩���@�SO	��
	�lL�H>�n����;����ZW�i�SnU8r۝��(8tsw�����<�U���K��t�V��qt����{�a�����#�[��/�{�N����!�j^n�:�eWT�Ľ%�҂�Kč�D݉��t�u���ީ`�4�Kd�J��3�M����'�U�G����>Nr\��6�ǧ�#�f��ׯ�P2d~�����٢1��6/���m�.��q9��Цi8�c��7���>!Ea�4�2���N����2Cyy�����.dGN1���0��T��[�
4'k��l�75��+hN쌌:zz�2_ xH�i�?�^[��]�D��ZH0����	�a�^�]��E�v<Z�R�O닍⇇�J2��vlSx���b��"`�sb��W�_��e��6��y,��h��k�I�} m�	nu8�Q)�p���Ρ<	U�rK}�3i+�o&�\�x�w����Kb� ��� $|��^#�`N�@�-BBC_��C��	~������&/,))prq�����j/�+(a���_�+���)��T��:dus?�ux�hi5�ͧ��%�/�]�͑�9"B�H_)�6�'�J-��vR��_`W���	KʃJ���3-h�Z�3}�udI�Q1�.j(_�4�2�̏����"��KT�CT��kq}�d|VV��* �H333���J��T$�Մs��f�E����Z����v$-�����uM�Yg�_W�Ȟj����O���G	+���BY[�3��B-K1r�k`�EC��`_�n���$��*���:�C�ܫ�8?�큀��d�߿���EWvA�<�hcR�/�"	
@�>w ��}��].bU�)>�R40��$����(4�2�3]8o+~Нڲ�u<���-���:,d��ۗ��!��?����
h�i�M	��\��1%X[!?\�T�H����R��ܰUW�@�tQB�������'�M+)��&�
� k�D5YXXhw<�[g�^j`Q�B�a�$��R(�?���L���[����h���#n�:Y̔Η��}C@A	�)��'�������u_0��C��آ�O���_.F,�G�S��8��U�*�P�ⲋ��)�(ل�[��kL�S��i>|���,# o�N;G%����+	����O/�Z���g@퀻����a=��Qc�B���Z�2\��'`����)��JO���W!r�q� ���9)>^%�n��	_%|��FSH��u��*�v�=A9VsF$\O T)�R���%`ˇ1{X�����[d"�8������$��bC$�w�{-Ώ�s
�Љ��u9�*�X7�~)��#)�m�m�?̔i�B�^� y�#���1 d�
;t�ο�O�[�6]8u�4G��:ꖊJ���P�v}:k/�,�m� y���%~ge��p��Y>*4Iq�m�4�����8�|K%�����`�eC���t���>�T����zUj��-|U�Ό�����҅��]A���v� {SbL�?���i�l�Y�������.��� �߉
��p�[���$�r�tڠo(�d]!��&���L@"�%8
W�3+��v�����$$�d8�/��u���`]�� a[;>&�rV�A%��ї�2�8����g�y�r�!�KN���
��J�Of	��C�����s�N<@H@@@���(o\B�j�����F������55u;�c��ffF*3o�#ᢼ1�%$�~#Q�����ˌd�D�h�$\�Q�h,/�>�>���F�hZBWp���(u�'32��"�㳎�m�
Y��c�����3����BS�$�鴹�ρ�;ܛ,8Z�|����d��E7�AtT�{n'[{����)��!$f�����׬���x�.-��3H��"��n}6���W\�6�ƉA��@���2�66XncZ}����3IIIfxx�^���2���#�؊�n�cDA�	p,ena����0��b�χ��AL��a�Gd �T����AZ��2rN��� -UP�dF��"6ɽR������6���s��u����P���5H$�����j������F�3��g�BT��������h%�C�ȁFi�nmu_+Ӭ����m��}��/����n��zbGe�޷K�/��XTTT��������eV֛1�&v����y�J�h�:�r�����ӿ��01U�¡���3~���D��;a�|<Gd�x�����/���~2@;W"I�x�����W,��� c~W�����>*te�6�ܩ��P�@
I��!�����Z�-�QvJq��*��y	.�f������a�Z�v��^]�dE��-���kll����v�؃�w-��յ1��b������y��G�����=�hX��宂�n�r��������\�A��!�z<� q��yEV��T��H��ߛ�*]�*��ϝ��@�RGp�U���c�I��Z�kSC� �����\7�Y�pF�ee��hȌOM���a�A��u��1��_hh�.Ȍ;;m1,�y����������j�'S`�@,s�����_� -��������b<ڞ� 6�����e�ݳ}��h�<+y�4�^G�4}�jcS�=��pR�`}�
�&8W�1�m��z��%�� ��( ���@�����Y�@���Q�. ��Fv[[[yÃ������?�&Eޔ�ׯsh���Q��:�4�Mø�5�$&�.�Y-�����7xY� D��b6���hY���6�Q�7�&(��ciX@�P��8�+k�����8���<��͹�]�:�+�O���)���l��^G���m�Q���8��ٿhr����T�5�o�l�x�[�߾�Q�iTIh4YfWƔ��rȦ�l�u"B�B�f����@t.�"�������������Z'����8�>R���D ��zz��*:�	5K���g�Rk}7���x���W��$ɹ���jk##
n�%|)���-�1J�Ж�����.>���$JĽFC����k�����,�O���V|4폓�uu��������2(��a�%<ަ�~m����}!� )A���������9�h�ؘ�1��%��s8�;S1�ܨ���A(�y"B�111��FKL������'��@��|E>��0lF�l󒒒n�-�
y�q��������$��$Ͼ_u<W+Өuܛ�K�,fZ$���!�����\5z��B��Si��֒)� 4trvnԓ55�	3P�:��\��f���\?�<L���7	�3J|��\�*�����WGGm����%�o#!�sK��[zC�"""�aa����`8����0$��*(@X����ԋ"���v{�}�++x�Һ�.yx��K��}nRYS�A����X��h��9�N�.xZ����R��oc�9��N0��_$2��
8<����H�Ȕ�CK-��5Iĝ��ϣ466����n,���m�7�?~T[x���dH��H��e�����i����������r��xOϖL�j�����������g-�p�96�B�L^�����cp�ۼ�¥O+tm����\��!=SS��DYg�p$#�I�S:.vF5#��������tR'����B?�c���W�[F�ex�#�2].0�x��x9|��7�K�@_??/oo{k�O﹪U̞:YB||�TMmm;���%"~y�Y�n网�a�<��)��;I��I�K�#����x|2�ͧ�չ�[!Ȧ*�x�Q	}����U/��d j��{�nK�Ҁ��� ����,<Ɩ��W�o�P(��͎e��}��ɸ@�P���}� '���**.�NIM�;�����-	�M���gZN�COB���ݽo4�m���Q���[��G�j�N���x��פ�bP��Ἠ�
[i�q�.�eh�vY	bR�8>�{ �πAZ�YWs���ƱGt��)++�?\��K���KJO�
�?��X�}ߤ�7�-� \�����<�%/�iT[�T�j�p���ھ`���{������ݞS�,���� ��\�{t��B$�
GN��\�@hz��r�T}�\w`)qi*(ؙ��Tu-�]����Ȃ�����@I)� ǠƦ���
��R����F�m��!;o��0Non޳x>?����]9�u��EǾʆ�{xx(�����|�Y���,�ƭL`6����~:��W�XXq�4��]�/�PO"rǋ�'y�8���?���%\�mnl\Fr�����XHKjEa�|�<��'�W^C��b6�9����s@� ��8�vɇw�^(��&���}u۸���uX��%�y� 7R@@@Q��k�P(d�:qɆ���Jo���������H�׉Nŧ(M���:f�w~Ϯ��������B�)P1O(((�^j�������%ޜ�,ܵ�e���@��g�ihq��`I�޽�l�Y]]�%֢7a�L��ٯ߾���t�6$��*%��,�e��:�4�L*�����O��߿�cT� �[��W��R˦U*��əL����p�j�����A�v�t#@�ȉ������O��+�>"���.��4��ɕ��,oo���0�k!�������Z03�1�{���W|X�;�� \�қ�4:�m���at���K�._� K2G���m.W����ޫ?�=������k;;�Tϼ��0Y
񉈉�մ^�rq2���0�ݽXg����\﵈��3�ȑJS�2Y �4�6���8?�����)���r�a��l�_���b硠����(�K�8��6��r�ѐ�	�U����U�d��Rv�	�c�T�)v��e��qppP#���1�`�q������[!�ͽ~��?;F����A߾�&�ø�/B��[�	E�7�M?O�M���,~)�����A�@�`��:�y�o(1=�m	�H���49:6�v�ͽ� ��[ds��DKH�]��
�	�����D�"�AH����?�q%D��E�v�SUf``�1ȡqT�ZA�S~��`�.\)����7���7E�"�BV��� ��E�8n����7�Nk$����is� Sйh��Ť���W-#�d\�<��r{����?G��oD�0O$��p1P{B���m����^OlS�ҡ�wJ�V�Y�Ǌ���Á6 {W�u�l��H^I>�@������xDDO��	#�m�*�����!+J�O�U�� KW��yR��:�O�:Μ�S�w���~�22V�$�ݝ�#`OqX-lU��LKHH�_b���}��t;GX����`��/��-�ߧ�3�*?�����$.��˫�5��b�E@�wN��|N�)ǚb�`l������p�5���\�K��`
.����_���A��?������&bHԴx�>�&`��zs0���I�f@g�b$��k�Q|���o49`nn�9���^��O�u�����!!.�	��/y��X�9����n�B�	9l��PH׹i�hp~���?0P��b��x�#	��p�R�75;{�]j��4t���B����􁒒[�v,����|',��%��w�ӛ7�q���S9l2�;%�b>%)XZ�N �s$���R�~�z�(,L�DC��1��d������cC���,��sm&�{p���0�KK-ǫ�DÈy��߈<eZ�^ y��h�c-#'7K�a����	�QC�J�B,iiOE�b_B�#%%�L��2��M<�#ˊ���4�/�H^Zjj�>�tކ�u�Y�`�榦�P��a3�,4?_#��(��\���QʗFr?�
�f�������#����Pg�pp�A�(,l�9G��M���ȿ��0L��yB�E�o{U��J�6�h�����ayr�n�3�6�>�Ԅho�P��O�w3�˛���9/�UUT�$A�=f�YK��6�h�~@��s�c��5�e;{Cq+����m��_��*��wyn��"e��HR̿V�xW����<����n`ַ��z��ܠ�_��u�^a|����GQ��O0���+��{��F�x�Q:+6;�J��D:C����h����@3�,Ey8itQk�W�^UQ�e�MMb
,Fm]趹�����5kM����YM�L�RNo�G�\�ߎՁ{��͡o|�� ���z�R�v �{�֙�*ejGw *���a$ ����;N��\���S8̠�6�]�$��٧NJr�hNJ)B�t����d���<�Gs9�&�\�/d��x$����
ϲ������'l̀�Xp���h[�E��P�B� �A��,ib���>�q��*�v܃��?���?=;kbh#@�mgA9�1�4����X�=��������d(+�b&�jmn~_&�Sޙ.������� Y`���S.=�M��1����f��K��F���6���K-��_?0�I��H`n9���C�%A�$�^ٻ�E|G�Φ����Rb��Cރ���@6F��=�������[�7O��I���������d�����H9��K�*�1�)���|s��<��*&�GyM�x��/�����Gs�n��C\�����<��SY������*�a��Y-h�ޖ7�C�...�@��]U�i�Ȏ���Lfm����&����������k�f��'�����mmm�n\��MG��ǟC�����m7�G�,ϣ���:�Ka$L�ڋuV���P��J8f�y�L���^N��i�v���Xb��0;���K��a�Q$w�E��nؼυ�^y>����������=6���n^`�p2�O���>>0��\����N��11cΖk@�qY�Hy��@�� J�?@~�c�;6	��A"N0�aBwf+�(:�����rw���
��-pH?G!{c�!�Z�7�9���&�r�O������������o	*�.�:�#�%��>:��[k>���`�M�\�Iٿ#��$ r��ã���������X��vH8:::9�p�o��Ȧ�a�f|+�,�@�����G����Av�Y)(����U�$����j�&��@ti��!�sH+����L�~Q`s
8������ ^�ˆ���r>��~�Ǡ���]�m��Z�J�F��h]5?����|
�y�-���j���������qO��4>�X:��c��/�0��6��n�1�3�qZ���F��:&$^�|h��$t��ǻlK��1����&6� b��DU�f�������W�=9����rD�ڥi����Ke�ʘ_\|OȤ��]H�[Y�}cs��\��y������`������d;��5�j����SV�{�f�W�������Gђ���>m�[��Q�;��y-+��3
۝�!-����(��mfd``G��^���N���HK�jw��=!!a��3��(�R?NVZ�V�,>5�8QrX7=c�C���S��P�/,��Ne�bxo���$
Q��00�T�Գ��s�R�"��Bg�H�A`#\\]��!���o3�ז�KKK9	e�8��L}oa���-�a��W���(� � �P��J�����T ��������v�t��b�����Z6�f�ti�/�`q
�=uq��.'l�ky�����#R��Rr����x8'���:�1��Ǽ�?C���u����[*!�q?ê�D��߼��.�8\kϪ�� [YZ2T�OF�	-79��Y-nG<�:�S�8a��p9Ɵ��ljh8�������?0^?�2��m]x'��:��	e��ƝB�0`ސG �������ML��N��nV_ �= �#yyhF(�E22�W>Yd0!S�tbzV٭��!k����O�(��`N�ׁ�*�s�VC���t�s���M�%����ǧ.|G�ҭ�U��������]��Fԟy�-c��ti�)�?aE
�g$?�fJ�yA��G=�H~<�}ԘG�V��^X�b?]�"5�pxZ����Y��� YYY��H5�������`~{{�K�ׯ�+�r�dL�/��:*����tJ� !������twJwIJ7"�twww#�t���;��{�?X˵ԛ���>3{�Sr��͠*!a:���p)�D+k�b��n32��VK��O����c9!ub�S�{���+����-��wE�C�8���h����yͷo���5�����MK�U�J���|݀�P��q�5���^a<�nL{�Uq�~�ee�O��%��dݚ JlR�ՙ���[@�[�ŉ7�l���qqq��KH�@�JR����EF_hd��s�@O_ԫ��xZ��=�p�u��<2eOg�/(�5�Sf�H�r�j�zN|۩�Yd�(���Ĵ���p�Ҹ@��$NM9���8�k���������E�i9E^�N�%���S��!)Ju��V����r3����$�A��\�M��!��1A�j�R�ż��������D�C[�d���`G��J�r%@�TZ������hs��������hx�����ӳ��Me@C:���/ ������	M�$ߑ�><��?M8OӌP�C�j�o(��~k{���`������m�;v~S$Be�NԵ�)"畚�Z(�}sz�C���l1�N ��A��ķe8&
$�Imli�n0ӗ�-X�p�8
Y�T�t�W����; J�������` ���
B>-Fh�d�߯�.����	��a+��x�����pq�b�E�;�0�1I�yݎ�&���"m��>^ܐf��j3�4/��HKKK�S��Fx����u�����W#�'�)*~Э����,[r�P����9��r0�8@�{z)((��Ƴ�n��U {KpN�u�_U5@���}�,	fAM�͙ uk@��߾��vv�ۉ�[�+"�e��� 1�y�A͍}���_M�ۥ�������ohl$�����e0�B��Jc�$	A ��9�}y�����d����е���><RR\�b,��z�!)�$��R��.ヹ�����
c%z\�(b�h`bD��^n�l��ͰS�G�
���ſ�#��٢�SR������=8�H���
s��,�gG�jΩ��٤�V����	��L!��-i]P�m�����l�t����H��G���ګIxd�h� ���z���P���Xf5mI���)��Ho�yyyF�gӆ��)���JK�r;mXNsN������z��;�ҿK~��%�q�\�}8..�u/��t{@}��n�i��x�z�m�ԗ��mqC�c@	!�$!M<������<�AoV��aUݰ���t�5j�����⥺�c@h]��ò|�#D�A}�7M�V�MQY����C�����YƩ�~�¢"K�h�Khs[���y��8_
��F�oJ4!P���C\2��r����x��M����k$��^�@)��'��0���I����ޓ�̂��ǢUeb���G�:�l��
���zzk~V�o��m��@��;�O��{4�N� ωn7:��l����6����pp&L����R��>����ohh�MBJ������_�gOh#�4
����,�P�1"Rt����P8���!� �윜�$u�J���"w���� z��(}FVS��Kt_ZT�F��k$�6�D�W����|C15�-�b��300h�T�JĨ'���MP�,4�%����*�m��<p�y�R%�%�s|�Ȝ׻�����G���n�W|44�c���`{y˭�SM��` wJ��'�4��J�p�3�[I�A��k0,��-�K�C����NumMMՂ�9����)0׃��L��� ���R�=�.�� (�ʈzBS3�*?�&�fd,s���-�7"*��~;�%�S���z�n"5�B-���}d73�9ڤ��&�Tc O�^�5J4�[2�2�|����aNG�@�I������������p�e$b5��06��驩��{�wD�������8�~�K��T؇f�4Q<؇����lom=w ���,7;�ٷe- �0*:��$�50����u��fAl���Y�	��p0,�YK����T�a1��<][[[]b��
�q#O.��^+?a����;�'і�3�5��g|����N���.��\����`�2t�N��F��q��������0�b	�W�K{�5/vZ�Cc-A4�3HԘ┎dz������V1�tvvC�ٙ�ep�I��C��]xY������eJ�yur��7U����z"����x��X�%njjZa����T�|w�B&Xw��_�$T\����x�131e!#!-�y���8E����Y*
�&Б����w<W?�2uBqW[���N,&sm�H�b��@�cP��IV8�F0Y�~?n	d��F5p7�R�p)�jN�>]���9���)m��g�Gr������{D��Rv����F^��<b�T�щQ���*�$[ZZz��ǧ.�}a�5�+@�!Y�Ne?���j��5����0�ޘ
J}��!���B�ɖ3��p?��ѕ���`�t�&+"V���.��Mm�ʑ�V�������/N�Ř_��s��CI�5���|�B@Pdg�^�
��p@��_���ʫ����8���6���=Z6W.��?o�08��`5�&�u��^�� А9��[�w�U�7Ja��qr~�@E���c+������ �mGȱ�����à��w�?4GFS���C�k �� "2r�0=E�;�d��ûwJ��.� �';��6� R�Qp#���w�����%kߴ��6;��J�Z��XŲ��s�O���1ۏ�":P�hoH���)/���!|��w�I,��y�++��t8Z�x�7��hSS�٠v�W6R%�y]��v��ot��	�n�|�����݋"�c��)����R�pppx��x6Y�]﫡����#����O��A߄�k� 
C�0�]ˈ_��'V�g�t��K�� �������iG���3�����>��}�֛��%Pu�Л7I��7PY�������-A&I7������Y�����J���R����by��&���A EUeDM�o�`�*��Z<.���]��
����ᇕ�6�?���M�	}-�9��IESn�*:���k�p?��9^�U���_��:�ư��n �E�q�V��~��}�����z�M�u9����~LL-��5�bgcSʢ�-�}SA|�7CG{�z�$��q����������[Y� �j3�A��v3z�gz,� o��_�0�43{IE�I�������2̡Į;��K��q� �(b�݁WN��}ݣ*�q$SGf֬0H*(�1*,�8;k;b��7]�[��x�Hz�����?�*��'.|�g��D
�ʼ��O@�+/[���)/$-��ʄ
���qڨ�<R����ȥ��[��=6������)�ޤ��L$���=��6"���-�6 �QT��lF=(E+�G �b����تI��,r�ȼxM����ڧ��z/���z��eLٖo��L�FR��B�j�!	���.2���t�h"�NUuuB��8�����kb^�f��ߍ���{td���͍�����铰W�/_�2�tj�����g*폽S|�R^�_����,�{�# :5yO񮵵5SHP��"Ԯ/,EN�C! ��0�YͷZ�A���%?�ī���ы���1B�xc�RXX8Z�) �i��s�MT��+1KDͮf��~@e)t�l�3�>�os<.��SQR2�tҎ�Ґ�5��\JZ���Yޣ����V����ђ��7M��D ���tN�K`S~fW����%�@ғ/:����������P,��x��r��G9��>��U\�s�3�Y����z*������?C��o�)�č|OP�#4Ņ�9�?�Hg
��B����}8�?eKA3����鴵��tG�B6C��ZFF�~��̻�Y)o�,LL.i99g�%B1'�B`V��*����+Cm�ĺ9���B��ٜ��ʢ�0��Y� GJt��p	�w�~��'i���H������{x��#�n�S�9��̀46�̢�$������0��7��B�0�U�h���)#-m_"󎅊�O	��@Ōep�G�h}#�>�w_[]�.�&w�)C��A���O��C!>5zТͻWlb��	{�< ��5�%���[j{u~������-�M`���R%78z-v�ohAR���u�
>}]�,�al���)e�LL&ۯ�K���ʠ�c|h����<�]b���.l����O����q9u � �V�x �6�6~�|;�n&oҭ0��&񵡴xrg&a�Q+Q�ir޳;�\��p���yu�Ae4C(o�P�1���r��������T����D�}JY�Q��-N��TrF�JK�	C0I=�0�'�p�|�-OpQ8���$�@��B8".�-�8+�aւ�gz#	FC��t�ac��� !��S����,&&Vq{�N��
�ڨN�	�T��_�-���"?/*Ԫl���>팭��ƻ?�)���{%T����B�
|Ndl�9 ��O�j�R;�g��t �fcxq�/� �Z�i��2dm�+�����tdLX��z�ی�MX�4��.�6'�2ꖇf����3�X�wv		�P�揌�H���H<>>�IHH8��(x�o3I����n��9'P�1���yV��謞^D��M,�������8����,z-�ssu���l)Kw���ϳ���k�����=�; ��I:C���������9��l;��ש�����Z�ᡡ������a��c����4^(�}M�"�\�T60�x^ǃ�o�q~~�r{�S�(�\_��k�[c9�C&"�g#UL����# >PW ��{	�� �H�/=?~L����XxPS��|>� U��2�k`y�o7�a�_�K���:v�!:4�����EȾag��|��:�����ri!�꼄�~ojjj_KO��I�2����AAA�`;^ф���㡦�[[{�oiiA�X�'�fF�f$�
�4*5���(6��L�F����Y�����I�k�b��!�ׯ����x��`�2��tl���6V��Z\��#�~OJG�"n�]���>����]�*�Ka�R<#=� ���q\B�p���P�'z����|Ŭ�t�GZv�����GV`&���>h�V@"�b(",ۏJXD�C��U��j,���*��ll*^�9�ss�'�d���y�+����?<<�hw��#���#++[�b��տb4F�CVV�*��ͷ���S@ئfd�܊*'Ly���5S)���2	&]�h�&���Z+��DN7��e`�ݟY��J�Gi	�jz��n�/P�'���D��2z)�dadT8�e�����~��#?ߌv��C�Pa����LD%G͛1�����W�4����D�6R��I[��,V��HE��-�8�&���V `҄���xΨTT[��_t�C%-	11b;��s#�9v獶#�B��N�s,1E�p\�_�IIۉ������)�m�B��ە�?�46ޚs����1���4�q:����;1N��_
7����L9���c)$XHx:�k����E���{��>���Ѫ!����=��ͨ��5H��X�H1�چ�E�>�&�Û��D�n����
[�����5=�`����?|?�ċ��&h�%"%�%�4��}
y&UX"9�.��}���u{��I�˵�g>YY�_��[�����g��]����s�D>)C��t���<���`�}��/u���߾��*�!�����8J� �<j6����-�X�FR��u��p��v�`�����U-�35ot`���ɩ
q����~�����tt��A��E�7x�g��ik�o.�de�2X8:Z��l;5B]U<�tt	��/y��Yt1�hߦ�,V�vW���3���fx#��備���#;G�@����?�ȍ-�B�8�ځ��/b#_e��#��ݸ!��vUw9X�Kcc<D� ^��v�]����qNN���}a �0��t>��t�>C�#��R���S�ao���TjMz��:��������v��f�jړ����{���	YB�j ����`��f��{�G�e}D	��EO��"W��O�o	���^���_K�M�����[�aE�}�T �v@}�Pg���_ky�����Ng2Ԋ��r{��yɐ�ZRc�z��9�%���%~�Z%%���������D��짘]9L8����m��o��{@py�.6�S��1� .�ߦe<l��T��0��L#����tYf�o �)*++���!	Y��<;�K�;c������RȷO�$��a���w�(((eI=_I:ѐ#�'9_~��̒�V/��͈1G�{{����0qZr2�џ�!`�0�jO���S(MI\f#���I�2�)���L�>@�R���g92"�1�g,~���^,�����㣜L`��ܲ��{�D&RR�2��D�t��k܋�N�=??�:=�!�DJ��w�ۉ�:�Q mweb^�x^��b�����^
M@�i����2���`�QQQ���> ��r�0�H��	���~�M/���&�����䝝�4E�m�	�G��D����ry����%�p���ˎ��Q":�yKD�:���!A��Pf���S�j���x���2�o99g��[��<��U�u���Kg�ix�T�(��%��$�66����W�܌�u�-�z��/�?��Vt���?���>tՌ������U<��]���$�"�j�bk2�ll��N	�{�����z��=���=_��釾�a����,�:1!�! �ִ��{���ꪪ�ʙ�WN����*��ɒf�:�̨���|�O�O�vNVrrr"IIH�gArbܛ+[���j�@/5J���gapp��vS"A���E��;�����ُ]&��^���͹}�I���+��Ύ�0����h�i�Iw`?G;w2=���v�������4�`�;�au���~C*��Z�ZI���v0w�kd�+�-�S�P(�ѤõX�T�Dh~'ų�X���QC I=�nNH!���������A-'�{���9����O�>��0o�ES���tI�1���O�G�|�������o�2�;������ �ʞ�{^�^�bP��놊�wg��J�p�I/���*�ps�=�t%�g�s���,k#X�P���`b�50SM��H��"!�Go���@�|��埀j� !�5W��A�\��5��H�()֏U&�����yſ9�}��K��'94�'� Ԭ�o��+����ݥ�24�TAY�U�Hj���4������U���d��̬F�E�x��B��Eo�5���h=����i˵�Ǌ&���H����A["$%m�Y[޺���s!2ѱ�-VSb���Ҭ��"HHi���$��|��3Y!�eU��惜�8Ue���ą��ϟ;�H�+1
i{;��v`�H�&&_xxxb��]�'����z�#���_��p(SI�,uĘ�G�eb���兙���GZ�׬��В��W���5 ��̟��\ϟ��)�|"~24q�b�D2U*�h�b`�ZZ/��Mӣ&&&~`bb�q*ɖj�$���A�W��`�R��]ؑ�80
ɜ=��?��޾ͬ���-���ݛѨ��& ,�N�\D{�����59<�E�~	�w��X` F�״��K��x����Kל������o:�Z�h��3O�������a˱���u|$.���@��
���>e�ЈU������d���xߞ���M��/�~����.���la!u�)��%1__���2����Rc'XֆT��o�z��l+��*�o%$��(=�n������F��y�/.>���|�'G��?4�P�Z��0<^R:��Z[[+����Ӭ�N\\\����.�#��A,3�$�)�{����n�D�N��@����obAS��M�5$�:�/_����V.���%6]�9����Q-��ѯ_��NNN"{�<܈�5��Ƴ�Ȧ����L�M�"lO;��Ćҿ�> �|.�U��?�<�%{�<���~����pr&�k���`�Oo޼�����)z_��9[���\>[^��]mE�����{��3��;++�� ���{���ۧO�/		w�Ns���>k��\]��H��W^)���2>�Ɵ�0�����^ܖ^��jdd$�r��S��tGdZZV�^�ТR�����M3ȁ<n'kB��bn�裮?C����]��T_�����?u�ߗmH�� ���4<�������`I���5Usp� >�A���D�A8 -����h	p�uf���qdu⽰����\����ѯ��0��3b+*��`�^���j�$'�!��߫����LG�O|˄fĬ'Ult�#� %�ؽ�s�h� >�����O��b��6����"O����d�a�,lmI<.�d�o��f��ЫLѮ�>s�#E§��
n�Q#�i=E�^iv+7��[u�,�E{eDJ�ٿ��c�JD+�=���Grz�KZ|�VR�_���QGGǺT�*��\�**b�y��W�m���x�/%�QS_�R�eBZs�y��}Xz�kL�9I����"3��k	�XD��v�M��{3�u����-0Jq`�w�H���M���p�1Y���~�B��yd��贈�8�Y�E1"폤(�Ih�!yht���5��h���*��t	�S�,�5�d���jp��WS�)!��|_���AM�LX��~��������9z~^^�U�Ί���e�_>�"���j���#=��ķ�pҬg057�v;\`�!�I��~�P�z^�a�]&Fi(����}d�.|e88�R!A����2혯��Ô���) ]�9{���b�����f%ם?��q�`2=�on�U-�P��x����:������js�֭_��s�O[r-�{ߐ M���׃�Y�W�]!����}������0�>�}�B�����)����V�M�S�\��衜h��)%�m�u��D�����$�*�8\�]2��E��{�aB�*��nl��c"2+���	��\�YP�"�M����w7-�G����O����סQ����E��!�f����y�M4�@�|n�~�{i��N5���<��]��2ã���ظ����Q�J9��D�ЫprU�K��U���,ii!1���$!�Xip�x�>���;V����U��� %^��Qu/��?��޾V����g���?m�.s0�X������
��}����Ʋ˫+�5��7�+��V}j�E�IPQ^>""�͐��w[[[�P��&�.^|�fB1��icK��NX�2�l?f�T`+��Q�>XG����2���0�F�������ǌ��3�f����H�҂��D�������t������� C�v[oGq�(@� �0��0�j��r	���11�)�m��$�($�@jë˔� ;�E����pmEE���K����݀�_x��c�b�c1� "�"\$\�$̶b��)��-�|y��&����_����U�[�|X�SCN��G�84bO6*Ò��6�4xm"G��1aγIl�鞾�>z��G"#ח28-ߧ����.T�2S�_����q�����LqH۫�C�"���}�T���SE��,�e�[~=�{��םo��S{И�@L�-**����4S_�#�_�4�P$�b�7�������㽇�J�L�y��NH	{��:K�7S
6������T�D
��ܚV~�++ު��-�����m���σO�������qu����J �k]�ਙs��;[�jUw�k��a���֟US{���U833���4��������Z}6�1j���Y����43�,tt���¾k+��L�7�\"�f�܎u���貊
-�
�y�Ŵ-����������<)������6�vȬ6u}/V�6
��4~�o`�!_��aaJ�9�l�55+���F?(]4\�j�*C��/U#r��E4�v{�-�J��f�E�}(���Dǭ����������P�.�/�?XzOd��5���x��np���N�<�4�j��DG��5�4Β�qu7�Eߪ�8m�.G� ��x%x_x��a$�(���f/��g�FuQK�uB����b�JG+�}J~8�R��w�����W�@5;��;/���	������t�P�K���;���> �y�~qe��P@�m�9NU��\��Ȅl�	�t���W���v���P���ʜѭ�_�*ߕ��M����2L�����4߿/���>�@�Y�����Q#��V�'K�d=PV���+�	8�N8��+)(��(��bfM��%;+G KI��@KK+@&�>q=]�L9�K�������}�����@l�|�$����WR�W��ʁe�D�*�Էo4��Z��L�����"�?߸�]�9�w}2��\��R}�$�y����4�(䐞F=�"|ĕK\\��`*!�O�44�M!!}���C�p�({����W��%�}]�/�`b��K~��`i��z13[�HJ2A�𚦦�>uK��ȁ��`��)�����ǡ����z�z��5F	�z0�� Yb�JG+��.L���*6y�F �kV�\�^Wm�� :�I��oK��=ŗj[���A��I� ��嶍���ÕVd^�,744L���v��q����WU��#`�#�,U������/j(]\�s!f����ܓ9^k�'�j�D����T���S	HK���P�}�XM��0�66����$�uif�O��U�B�'���]\\8>'Emc���������b��=GY9�tx�
�6���2���=ډ_�fHKM�|�A����--�) ��~�^H�=��'�A_gX"��j>���i$���ߧ_�K�+p$KU��EE{Y�I�'4X ��ϛ{[z���
	�����G���}/Y�� �<�,b�����M(�)��x��0p�����LLu)II\�!��J�����Wʴ��҂��=ag𚵡�w��\)��/_#T�Nc/�>fqZN�544H��sy�+{ȵ����U�3��L�;�+�j�?�������B!p�G�o&�,`���8Z%###c $���k�G����r|/�����7Na����z����=7��Vh?�̦�{a�dG�,����MCA�)��a�T3hs{���Y�LBU)����Z�RfLeee��� �Md����Ε������mT�R@�e�	{k����Ջ?����I��U@�(���ٳǡ���^�w5�WS�%Δ�_�;���`ccS��z�p:��}�0W�e���O����*��P�)z���K���0z��	<�6m&��ճ��{�q�%�����T���_�a�ţ���a�����D�׵6�v��i#�Q5C�F4?��m000��

b̹qh�n�{;(���/�ͮ/[��VjՆ���'�2aVUU5q�ShK�y@�j	���?��*[W��=t��<�泦�8��w���՟b�E���lnn�Ad�\lS8bmn �KX�MiQ�V�4�k��DK�3���fuh��{:��B�;����65�Ȗ-ߧ��f�_��_jp?��^ޞÛ�.fptwuq�m4%"�����U���q��k���B�e!^����ZD���L&[1���̤��I�r��=���Z	+jj�,���*6��K��#����	����N��^+b��}Aq�!VB8�:7��e�P������8���Kb⓱��=YY�� B8T��,Df�2:999U��4�{piqSS�Tfdh� ������򬐓���50(0P]V�?��45i�����XY�z������uϘcz��I��W1�.TutV��zY+)%#�j�ԻC0DB?�������3N��r�v�
����b���A��ʘhk,S�����=5�����ֹ��< ��۽��4���1�:�]�Ɲi��)T�,,J~�<V���Z2��£��zki��z���~+-�id��b�5 (���ņR%�&0�/ɁFU��2�g$��v����L���O��X5��Z�z�������p�ǞP��3�0����_���@����l�����
;��-��|,�v6�𫋋�ى��½�9���S�����^4�W�h�?u� UK!tL��rC��#�U껮�x�Cs��Z,z�A�o�Z�>�X�eq��`S�R�x,���RBes(�f	���wy7x �&� ����쭥������fO6���L��u@�R $�q�����n2 ��C-�����g��;\���%��2m�p,yƟ�˞��G�
�� �f ʳ[�L�
��5?EY�0!HV��@��|���҉z+6�����***�(z7��]ز`r�����6:#�И7eT/ÖYPPPH
�8^�.+^���e�ڮ�7)��U__�KKK����Z�H]כ\JR
?Q������rCDFֶ��L��}#�))��KQ����=?9���ÇD<��
�@2��	u�5���B��x�����e`�����V�-�TZ�!��G㵼������ã�$�܍n ��7���=�P)w��R�{��h]bb��t0�P�"'~��x�0����|y:�譹�qք���f��*�@�k�1
95$I#���W/_6Z,V��e��%�UW�f�9A�����t��byބ�RJ�ڠ�1ˑ��\LՕ�o�Pq�;�J~�ũ�Y��k	5\4C�zc�ynAa���+<���N�Ҧ|qc_��ʚxl��(�CJ�w�����yQ�^�rC�y~�����4ʦ���}Z^�?>_NiTT^||��M�/I,j��45&���mml��fl�4�}�q�NLJZ����cҪ2��uF�U_^\,�.4ൗ?8���䖀�nO��������� F]�ӧ���`@kF�Of��r@�^�d�e�`&R�B��.l�F%;V\P�vt�njpD����DNw+th+��ތ��Lt��3� ����~��f��K�!�\�߿'TY�{򻌾a����r����KnKK=�qI�<��?'�G}J��+�}�9-&z�uܧ M���GUSS���YS�$�G���
�.빬�f7e*mRgr1��7����7���"�K�ڴ��):B��1�$���k͜��NF/oq�����%��^ ����7�1���:��O;J���yX�Ev�MW�aaa�UFep�P��KO�<#c���1��[=��u�'k��&��I���rU %�ۣ����4��דя%���!��8;_�32��R������贸W^Ν>��Xo��;��Ƭ)�D�������)��-������F罩(�j��H���wO(^���H�~q�2���azIH�u(�y��1� �UϺ����/롫X�ޗ/_��7W����c+���h!��@�g5�S���Yi��MT�C�\���������#G����).����US9� "\����D���o�y��H�KSJ��V1�r��" )���J���켍�6uوKQ�������Gҹh�笪E����kW��=�7��+�tG�U��'�P�5���4rs��p��l,XB���UN����
���o������-?`���Y�%�CW�>^�
"�������$�����}z��s���vuv!�4����<
�%�G�k��In��̴�E�7f�0xu햑P_84������kX	���ْS����it�BB>�Zb����z�k^�D�x��g��>3�+P2��a�RR�qq��2��=Z����1_�#�e �e�y�x�(��C]� Ogr��D���._@#�hhh�>�����T�x��M=2�����	c�Q7,�/�@�|�&��Nye)�G~�3���E��ŋ?#C?��������jsq�KQ�=��Y���"���h�]�E:���vٟ�	x����u�ꧫ�k�8H�y�\@j�ne0{n�|�T�ye���SO���ɾx�%.����o�:GZ3{{�Oɢ��=aF4l�4鹎��}�1UU���H��vw���V���|"�j�X2���A�|%�;63㬠��e=�C�Zۛ����{��+��tq{{� ��[��ぱ�9nvv��_E�X͌���C����d	y��*(d���tzf H|3;	��1d�]�
nT��M����@D��y����%Q�p5�oz�.��{����϶�h��K�	�����w��]�hA�N�"h|�(r��7�/��H%���x܀h��mr��|q��]��f�߁8�QZ��g����Tq����X�WV'�Q��%����������A����
���7�e������Wʕ����S]U�����Mg7��ݻ\\�*�����h$�sq���8߼��
Wͫted��t�٢d-�hh~�ooo���*x�Іd�|,��S�c�-��j��U[�pβRS�(�L���O�����j����L��~raA����(�w�G���S�	 �YXZbѭ��K�̂j*6�&���׭.�e�����m��#��K.U�԰;$��#����>Y6�L�g''4��1Tf�l7�Z X/�U�#c~9X�.�T��ԈH��d��;Q�ft����
����,�P��N���Е�>k\t����Of6Ҷ��D�o��.�+�g
�L�_�I�� ]R8��bFGE�v�r�}�U, ��>V'��E����4�?99		)�;�}1&�N>�� Ch'�7MΙ8Y��<��/,�rzyD�ͬV�q�ˁ:����f/:3�4����Ժ@����J�sx�x�^���C���}Ū���9B�Z .?@>-G�;!䅎�s��a�ip(��0�EA /�ol�p��	_cn��Ŏ���x����ǹ�Y*T�~��$<���P��z2:,=;{_���Zk��Fbbb>�(8�TV&U����p,��aL��9�D55S�@,���{?,��LF��HXO��-{��<-G��~�k��v��r�L�x+"t�o�.w�
M���xzjJ1�I���hTG�(��Jx&�l?��2�0u3�Kutu�D�o�IRFy�����/[��/,Q+QG�.��m ����+�Y��S��j����ee�9ܜ�bїY��^�w}�(�΄�INS�����o�^�݉�o94���f�����ۛ�lƎ�^6�(K�ˆ�Q�f��b5Qc2%�u��2��МIa�ߏ�_�vAJPtC�u� "�o�o�Ѹ�jD�`��P��������cjVI�j��RF��Nk������y^U�tb��ǹ�?�g�k\�i�c5�(��H?�%$��`b��UWGƫ�gg�ػ��g��ׯ'/�7����i89g���̾o	�6~���9j;Y�۝���6���(�K��{f�{�()����?��$(f@�Z�QBn:ͮ�0د�ѐ�ŵ����:���z�ǋ�M�CU6+�$��9�
���Z��|}����\r�MG ��@�[jd�=V����2��y5B����t0�z'�3�����!��������F��m�S46�Ŭ�T�4ƅb�mr�{�
��c����JDDDf���%��EJ�`�ɂ�0��<ö��`�6��0+���PcB��<K7���4�:u��E�۟4��5���`�Ǿ��@''�ëĹΞﺲ�&��r��--ꀞ<���r�Ѷs�������]b+#�k��C h󕒊
*>��u`#�f���켔v�+��d�?�z����I����D��cL}��C�U6ߧ��?���q�o#��KC��&M����annա�?��\c���7 B�x-��@�g�d�6��OetI�3�GCNޱ8;�B�}��ņ)%,&ؠ��^��3:Jk�l�sʐu�`x�Wa�z/�=c�T�Ƙ���ZZ��T�v޹��N܁L""����I6���T��E��Kx�ѻWw�bAH�P���rp-�BW^뭝�(�ݙ�c__j�2hM�`6f�#�'�#�)�#i����ʚ�-���9Bn�z��v���H�<��t��-�
-��d�ލ��H � ���<�l��������˅]�?���m��$�||� �/"��Bg������m@6��ȥ����tZehgy���A��U1A'��K5ݥ�1�ذ�8����L5/^� ���	�D�'M٩n���p�1Ύ=@F��f��o:S��cdll^g��hZF�@��\o�㇩��J\D�M������&�v^�r�ƅLR� !�;W0n	�Ǖ���BK+�����a�7gS�6�_y�؝�j�RSS3����.\��z�EzZ��kz�۬`��C�Fp��W�������L� m����s)/$
�����u"�tC��|T�������5-m:t����~;�,ZO�}�Z540*���3EuV�*�1�}�e���ϟ����� ����H܅�M������ �`t1��z�ƓEޏW�LL#��3E�V�2�E��y����� d����mt Jv|?3��|{��I��?:��@����T��N��yfO�/BV2��
�Jl�Z<&s�"�n�¯)�f`��P������No/v��!'�-Ց�Jg?�����t�T�z/�"BH䋦��d�����|Ŧ�,�I|�>n���߿�����B����2������b?+�Ȅ9��neM����W��H��Uy�\O\RT�����?y�����-���w}��)KT	�`�΀���d� �"���ߏ��|q=��T\9�=�4���H�<Y���\
Ț���\E�Ȩ{(�S� VV�O�d��Q��t�����iP$l�G��01Id�v0��E�eIY6�-V����x��퀥Xnu&f^�)>>�H�3�33L����Z����,/��Q������o��l��qd�����4㣦6�e4��!�s�߱��srrHIH(�%�n3݋�FE�����Rr�mR$\a�;�+�f�dl�k �Q��J�f�p��6b�1��K"��׀`Y6�S���(�'��o'+/�pr��|��fϰ�9��!JL@�"�;�)4�o�P�M��/tH�ts�[Iqǥ������ϙ��|�Å���a��(��j��5���7C21�,ϫ�c��[&���)U\��[ys�aqn�~�LMy6٭6�L(��׽�-^�.���ٗ��:P�@�}�P����Y�\�D�����*DD��+�[��wP'_� �P�~�9V��t���o������>��Gm��ϟ?�9�~e��=�ц��*���iy팑��#b|ѽ{�|?~)e�Z�5��Ū���m���x||̒@�,���/��͒�homM� l>jC�MG8�����ó��������R!�0)#,�l��~o�����l�i����wm�j�cȲʴ�TL��$�m��G$d���<�g���;�:)�Kq��������c�B�bgJ4N�.`��.���g���"�%���	eBC#�x�����߻G
��Z::`�)���ՙ`���*4������_{��O������Q��2�NƱ���-�GJ���efdY!D!{D��u}������������9�}]��|^���|��/9�0|��/7\�X_�����ݟ��v@i����y��ԲL���Ĩ�U�$\��%���)�n"�~��oUM����"�\��7qE&�E���,q?��j(�-kr!j" �ڐ#�I ��sg�d���ͣ��]YY��n/���?uo�d�[�C�@�C'�b&���8[�A��(�L��2;+�zȱScc� ��1���}�2:�������doB؊���ӵ�M:y�%#޻�)����G;�v�Vx�)^ipLqW5�a���p���J�φ���&�t��a�wvu��X8�4�E�G��5����?�,��Bv�`N���w]�
�'�9Lc;�8k%hz�����Z׋�(����fSW#�_��;:����5����������U��mRRJ�u~i��꫷q%�I@ְ�}�Zz�M�dbb2����D�ǚ���8�z�j��ӣ�+�Z�"ndTt����BBuE�G��9q��2�ܓx�����+���9`���F8�o�<���ʮ����F���\˙]�i1f�U388�pzv����[#�x��3�`A��0�I`�����o+~��E��8 �fg�9DEE�P�o!d��AX	~��]�߽AȔ��,v�"a�FMh��A�}�Q�O��6m��>!2���o�Q\��4���S �i�x㶠Ovb"/�b��|��A9�tqF�������q�͚��ux��9�����_l�Fl7i�2jР���W��f�=v^C񆻜�7"�����X$�%�9�S9����O����0Y���&�-�,D�:�&ʍ2��F?�!9N�<�.(¾����(��g�0P�H6�3���F��/��]�[i/�q$~-�5z�-'688���Jr3s��0�y�ƨ[�n���ܹc�V��������v�c�vt���.EG���ې�'�]]�]�� �nV^�yk\�?=�l�2��e���A�<�"s���T��d����	�;թ���g+_1�B��sP���O*N{�>���8����8��{)�7�;��\m_\�5�b�3��� ì��w�i[��]�&��ƨ��_og@��i�ĶV:���n^A�nׂ�Ǻۢ����rV���+�f�)ᘔ,��.ئ����B���b�1Ma��]J"�	uz��ll�==�9---������u����332�a}jn%�m��W�r���ےSR����������]֕��a/���<�EuV�H���ζ������F�$��V[t�������9�W3�w_�򐷶�r���0�.�+���rQDHX:���􀃣��Ц{��b��8�^$tt΢nK���"0 �h��*��Fm�g[x����H�m�i��c@�3�v@@����<a�(���	��M�u"�w/c����t�g���nJ?oN���*��3�E��o����3רV��7��Z��s�ZOμ��Y9��o��W���&,,,8 SL:�d�a/u^��]\||>A~~�Nkc6|b4�
�s�uLL*�_&��й�\G�o@���w��BH+z��E��k�@�sFf�#����� AWF�z�NT�~Ї~߆xt���M������ޑ׉sơ�5�h����d�E��X��Q`=�1�D�E��.i�xP�X������'�>��oc|��9�ǏgRd�+�S��v1K@�O�=b5UU��Q������ۿ��`KP`����b�I�<@o=a=	l�Hr�bS�� 4\�P�b0]',<��4V���o��iI�)ڭ���:xi�e|4���8^	�%�_amfVu՟�q��]�0�pl0�a����YJZ��>}��UhW���^8��[{u???�����9R~V��`����w?Ya���o}t�@I���G��w5�x���>�9���}a�l�"� �߰����Lc3�ն�q���'�O�&ʦ$@�^�5�C�w4��q*0#���-U]��♧��'��Ǵ�j���CT���S�r
g$��Ǟ��<�M�z��Iok�m\k(�a���u����A�ƈ�����j�rm$/ޗ�Av)��L�)�!f���R�:X�F�D���O�K���@T�eea��=���2dF���JJ+j��CH�!@�~���G����3__�L�2b��*�1�Hh$����ӛ�so��h����_i���@Ki��t@ �A��#O5A�ɷ/8�8vf��`O-����y.mT�����@-Z �i���#�D�X�ޱ<!+5�G����*zG(���"�('�n����9�OxsHHH��T&���E:�<Yy�%��������a�#-컂8��Bd恹������I���y�=ª�ԧ/g�]�>��Z� ���1L!�PM�V���^,VM�_x�ᢆUM�������4�%%�54��(��t��Ba�ɚ�������ӣ��x�/\$������,(�B���,]�!]J�d�A��D�D?��iMMM��V T1b(SV_��c����ֵ[o߾U���XyE%�G#w�E�#��'.�a���p_߈�IQ>Jz�\���_~g���C��鯥�K����^+�܃B\��$��xTR���0jK��iu�����#�-���D�%İ��������ũ�����'+o_<.����]y)uK�==H����xy���Y|7k�+��\G�����g�m#}�j�#jƀa�S]]��38�/u�9�<�E�
��d-a>����k��X'�̡#r��>&
�3����q�6���H4H�R�$�IV�
�M�E�2! ᥳ}�$����7<�h���ײ;�88P�*�&X�S	����VJ��'�����;�?X����fF5Z���ib-b���B-�b�c�kk�I���"��]�� �<�vy~Bl�kA����n�9 /g3!!�`�4f�d�S�U��[�E��q�y,�'WHJJ��.`"~�D/��ƨ/3p�_:HnE���aar��1hL��&PP��¸y���{�]Y��ٙR|ch���Ш��N����Q}yy��R��aӓ��#z?�}QTr���_����j���{a��W�7Ҥ\�B�K���:�TTv����8>,��bB��������$p����#�y���� �3IiiOG�-{|"1p���G�4NUH�: ���rm�"���w�*U#�Ӕ��邲��e�>���ʻ.�AL$���q�x�<��o�wz�~��KQ�h}������˗C;��J#�`Q��zdq�47:;;���[5�$�xvA��D�*/�-�(˸ͥh�[t�WUU�������]��h��w<�n6%��Y��®���`��9���ft��(���	�EA1������ե%�'�o8[`�t�b���C#�0Y�gf�~m�s���J����m�g�W�)aF���B��BS�@��Bo������$Ȓ�r�ړG��������y���Ys���'?�C)a^ᄳ���Ktc�����W[8]T��a����v{$$$L���D��ӲsB�L��w��$^Z�Nd��ρ�	\t(,�P����x�=#Y���]���eu'b�"��V3�Ȭ,��@L��r|~��T:VD������բ��=
oLb"r�B���W���6}^��%���K�r[^���P{�b+��˾f��q�4��2���333�b���O��0kbd lE��wL/���"к�Q:�;��s���[ ���<JR��0�p�g-58vj�L����
:�uJ�0G!�2lo;9?���(f��KK�^�s�?� ����QQ�8 ����q�v���H��F�K���Z�|�̌���T��P��=�j������QQ�	S���Ղ2h2$����th������O%{�5�U_��{z~BuBҌ�PTU �:h�h��������k@���|���Wp%��3��d�{g��4�����*�jj�P� 5�:N:��/�*�^��� �u��fBc�~����֤�$�7�c�e�z0Cs�ކRg���7�FG��פֿ��%#q(�ȑ�V����L��JV?K��f��
����[����݉�X�����4�?//)9e���dۭz���{��A��ȁӴ�牎���=qt�iC[k��������>�C�ɜ������ʬK�� 6T�����Jb�8�+�[�����ypf��HSpJGF^�;S�r$�a����m ����� ��ɳ(��#��?��J0I5��lx��;
�\�YF�c����ׯ_��O������ Y�m�v�w��<�k^s|�܏��>50H��F���U��C#��B�4>F�t��ؚ��§��WS;�韡-#`���U�qtp��	�y	�r�"�?�x���}S�'���/{-tu� 8��=�vD8;XA�>F�9�RcJUHII���y�1��E~�cו���ȾNo����.۞ӱ�B0�5��r�l�@�F�c�]w����68�8�w�����$����_XX ������x�3�[�z�E��(*�!',��S-�gz�]�
��.�-����+�pdv��c�������d�gg����D�~�N�ۄʣ�11�f���TwUK�52�B��j -Iܾu��`g=]���×B��7�s#?��P�`*|�^����D������?�Mr���.�w��RUU=BM!9���J1V=[U�x2����jO��.����./+<�^�����7�^��2����� �ccG��!gm]��9<�O)�aa���4?�蹔�������~�=��qpx%_6�A��1�	Ǆ~� ih�t�������{#�`������V�D*���M������F�`x���}F ��x�cU-}���r���LE^WU����x�=�u��g&��e{Rn�@����ʻ��v�j�k�A�^&��X�1mk���9uS{h~!�_\E-t�D`G;×C�0|�Z>}��$���N�6�2C+�ԗ�u��A�bZ��g�������mY�'�&�Eaf C�`���r�G<44tp}[bϡ�\/�v۟+M����ov֗�:�C��`���1�}��YY��8D<��?�΍���R�����]$��V�DO��ynN���4���Ȉ�~�]x7B����Ezj�.jz�9ް����R���mr���;�`b*�l��W1��]���%�V�w7�-���@�ʑ&trr򣠠�|��`b��17�59y���t-�����{�K�\u3�j�!+k.aww�ٸ��o�E0�;UvT�e;H�]�|�ųD���|�dF�5�z�i_��TLj�l����������wΎ?� .���@q��	%����f"E���$8�Y/�/؝5��M��758	l���Ӵ�|$�6�� ��)�X�>|�+ՠ�����/馎�N�+W��[�hw��f>��o�\Y\����J���o\LT���r��#��0�/�i,$~k�j��[�@S]8;BFN�;�@M�D���T�3<�vi��1+������iq׳�X��rY��xY��yBBB���p�Rc۱� /�25p����dud{�+]Y7�r��� ˞�pr^��DM��XάDB�s�K���9?��c;�È$,
t���]�M�>�䙇��.�찈P�Ǹ_ǋ������]��az�p�I,%G*�'���7i�0������pxy U�r����~�
Lz�b5y�]-ww`�<�śL�\F�Q����J�[������f.�^���S=Mtln�U�� ��^���0w����t΢y!��d���,��ǃTv��h`���?�;Z���Ц���1@�*�����2��iF7r:9��mN�G�pS=}���ޞ�� ~����Ya�q �;sr���r��!f��w�ظ��5$Ŭ�MN
߽w��'��._���u�N��>�m�����'iq��ʻ�p�����u�c��0 � ko[���1lt+H��U��A��H!�����t� 6�g=Z^^~���l/�s�݁��)?-�:��v͂�!+/_���/�@�1t�.�.t҃�(��������dO�d�����ߢ���]|cq��	`̔�ZZf�
��}^p�*�\�G$a /D_��W	�Ot1����ё�2�=K�~������q���Ҁ�߯�5B�QChԍ��-�	�&:;W ���"a%T�w8q�v�yoI���+���Y"""�?~�khks�4b#$&�G�����3U��y�H	�uk��*����oO���脷-��R����ә��}
��q��7�%CN��+�w �3vt0,���LΦz^ћ�v�]b='ߝ����FjP�ԛ�jנ��$u L#�xRd�L����R� �~M���#цP�`l8!��D+���З�(���tx�uBn���{AV��Lz5S;$c�kbbb����MYN=�
RzTG������>�.�� j���e���ӺYȑ��� �e������ŭ&s�]|��Y�6�Ny2BVފ�v!i����W��UZ*���24��eu(�������N[x|�[��K�Ǫt���8��_7NOO���+[�FL�;��y/ۄ��.vG����F���R�SP��V���J�X�_�SU�1�|�����,��4�Mi��F=dDXb�F���W7 ?< �EO�g���v���>:��*���+8��"���[������e(�"���Z�Up�'m�ڕl4L���P�����������u{���_9�ƈ$�͖��JC���8(��R�a{F�CR˾��&Ov�������$�Ӡ���v�}Z��o�z1 �-iikۀ ;��/���>HG�s�Lׇm��J���c���G�ߣ Q��'���P�"0����K��4�E=&��v��E�.0i[g�����\u���;<p��O���!U55,����ދ@��c�,s[�����Μ�o�y�4y�q�=�F�XTO9�؞���P�n�q*#��̶f>e(�!u=��vyjO�r�kݮa�g��M֨$�s�!�~hV��Ił�_��_��0�Ekp7EFF�!"&&���w4����H���[;C�!���U�З�U=�E�L)��%���\ �����JC��0h����q����ͤ�Y���t`�@�W}��1�q^އ����	w��kO��=�9��ݴ��Fm�C�n �f�T�ܚ���퇵���2��i��lllD���������U�1��<��8�zll��)�j!in�p�u}��Ƅ$�����At [���zز����=SS�ڊ
'�,��R����d�"�O������RV��U���}�|��^-�`h��n��>9=�Z��iG�bk2��U����!��}RSS��o��6�_�e�"�Io���.G���7��E(���o \\k�����z�����#�Pd��Bj��ohHIk���67���t�ֵm�69���--I���G��R����_���=��,��Ļq��/���9��I:?��h%��A�23D1H�Qh4}�I?�Ӑ�'g0
��:�;����*�L����8k�H�B:��4���k�����Q^�����`�R<��nbX-3�Q�Ԏ
��`g��OH K�r�w�޽;~��J���F���|��B%YA��5+O:0@����Ȳ���?�6y$R��e��6����z.'�����OK�[�G�l1�S�@��������lד�C�_?W ����6���;�������R��!���8��ĉ��x;����&IH�IEE5��767�wF�z���4TӇbdd5�]x��~��,��S�Ғ6���v�����KI��%���׿&b�Ea��E|���@�#K")8�{��ރ�.{���<�@� *���n�V�*�FN�h"�+��f���G�A.����b�����6�lp=lkR�=�� ��,�e����2���D3O�����`x�;�囼��X��imj¡�0���vW�L�鐮5/ X«���*vz��ڶ��ۿ���X��kZ����K�Tn�wX�M��"K��`k��=ce-�y�h��fB 2?$0�~��׮��p�����W--��ҟ�����Ȝ%Eyu3���8�Z�h�ӂ�6����n�h"W��a%�<����MЩ��#�Q�J����\ �նA
��^2���xj^��ǂ��WPRz�}uy��n߮��;�X�~��b��l��S]]]��?+Ӆ�M�D���i�Xm�|���ł�2�������|Sa�n���o��\ߎ�X�� /���P� �s�����_]U5��`M3���<�a��&��{�@�C+��%cj=�����n����K��"̻�6�^��_1������! PL�ڔ�h�(bǵ��>_γ�|*߽�k���-oB�=�vO���aߢ����ְ���"�{�#x��ٳ�H��7n�ֶif�V�[X|�7>��p�Ϛڰէ��v��|r˝����:�$QK(/C@H�5u� ݓblU_*�&���;X��i�N�o�%��.�~��6u���*�|�m�~�{z0���T��Jw��Q|�=�̱8�Fϫ�ZZZ�uuu� Q�**.~�ત�A�UޓS{a>/���/z{~��=-^�Q@�%���n;�Of���`J�Jban��D���>)�ڌX�1��3z���:��Kn9��znE��k;55%@br� _��s[�^�1��
�
ܯ�2��F|A����j�]A����ƈ���uu������->+��8��q-_+��E�%�u��VM��i������ꑋ�Jޏ���	QxC�]D�8�KV�Á[y�qW�V�w��%rt�dy�a��a����f���|�+���&�8ޱN�"Hayf��F*�d�����J}TdduTLL';��l�PoFj�R��,�sWuR�`��� �����C#�w��]�#�Aw���b��p���Ʒ?�&��I�_��5�����=�9j;����֭~q�&.J��i�����]c�5>~t�\�r-��$3E���D�Kx~���q&�/��"IY��|�2�${�B�ޘ���ԟ2����t�ይ>8�����a��?g�;-]�@���,T�ŁN �)�r���-)�k�zFŅ(��4	j�}Kk5��A��?�@���0�\�ˢ�I,�5DЖ�� A�����[�9?���S�l_�߶����O+�� ��.`���z��><І��������Smpve�����w� ���|iLB:�݅�8X���^3��Pe���2���*dr,$V\%�������?S���b���	�֓A�@n/���;/�������bMMM'!���G���'��-3���r�W��؞�'J���� gщy�76�-��^C.�ޥ�R#Z�N�	��#l��[�%�<G�����}n�T �]D'BR����9�kiHe�8��r�#ZȐr����D����=繖���De/k�� g�zH��B��y��i��^3=244,��0�1[�N��x��p �8������,�M�@ ��������#X�����y�&�;"�}�X�Ϗ]{�)y�@�l��t$Y���d�쁭�a
�Vl������i�kr�*�
�:u��������c�t��Yp$��ٶILb�V�����"�P/� �J�0ip��(�D޷�
(�޻54J��/0��f�R�?PZ����2~_+�,z-���\��8����j%�ⓓ�O�/{�R���N�\�/�H�//-�Bu�UNNN����p]]	3vMo��۰h�\�Z���-����R�lpn���(��DÉ�R�4/+�vU]� ��W�����YE��v��YK��_x@3�72:{g�$s�V���E��?>���θ��B���������e�@Ōk�F>^�(
e�H�a���Ȉ'�&Mx?#B ��#o�&� ͢W�����X��.QVgaH�e�kLъ�]Ę����7x�AZ�����\Lo��^<�y����'�t`-��o�=��|ҲU��v�
N"������� s���~�>84�GKG������`�����X&���ધf����KKK�j���p^�I\���(1Ǫ�n0qC����LLL|P'��ϟ��D_�\�$Qܕ���ž���o�o���4�X�<�J��)`,��������[z�b?FG�ރ�?o����8�a]�ɓe7ף)D�c-�܃�m�n �`���j/��9����ł��y�xwAz X�������s���
�ӶY�)��2��ո�|6Cޫ���xSvMd�z�ʽT,n��*����X�A8(kwc�TO�h_G_�����A�S ]�F<��M���
7$��Bշ�lG�de���:��WM��q��gڹ��a�I��J�Rj�k���o�����wa��DAI���oCw ((HΟPRR2�$#+JP��d��� .����D�eKj}$*er|S�j���b�F��°���x5��O��*7�}N��\N0Ei�B���u1�}�O./+;�S��H����Lj�n�j��2�@��:!��S�ș���v��Jc�%�~-�o�}�<d4y�E�y��S���Zg>�������eg�+1m����
���ˆ��-e���e���a-`��X*WhT0l">K���Q�Oô�rs띀�S��[_ �����i]�����\�=U��ו��g�� {v[u���o-��3X�l��~
���vF���+�0�c��`l��^�Kw����ʇ0Rs:q��hEe��b����.2� c��o̼�H7+?f���X���G�4�99��*?ʍ�6��6/�u��y-<�B�᪲`�F2���`�|rN�0��(8���QO+�x��Vd]յ��T �������*���zA��z��<�z$��g�=mpj��R��זa	��	�o&n��|�ĺ�l�a#�l�B�G��u?��Hv}�_����>����a��z��K��_^w�]Zܓk��g��"�0��I?��Vl� v��Ԋ_���1l �!��2�{Dg��_��^)�u���`��ґ�Il��G�nMEbccC!�]��K9�V�����Ur��f 0�z��sl���\9s����wQ٫�&Yo�nȈ{?��ct���D�7�>h��޻mt��vڮ����|]z�g�	0P��T�{��D�hH:�u�� � �s=))�����aH�(�->b�k�z>M�^��N1�-	1�ۗ��U1���`��fn�1b�Fy#���=8G�А���Qccc&H0�L�\c}���"��3m-N��PR�����k�9�ߞ�R�>��qe���cR�CwJ=��y��yPn�%c�,�Ŏ�7��-�̷
͹l�;K��b���R�(�L���E�z*�~�	�+^g�^?�)t��L|uJ!�>|���{��rz�Od��6�� ��_��|2������?g �S�W7�r],00p�a-��r������ہ�}N�~a��T҈���<�S������0��k��	�A�۟�J�u�ֺwsK��D�/�dm[-�"�T�9�U�7PW>����8>%����c̻p�Otմ��ɍ@B���M:���o� 4:��ɝ�F�(�<�ʨ{�#���=88X"����աL�E�o�����ۯVF�� ,�vW��=�A0Qop�=U���gm��~��CJ�z�m�r|477����s�̤�ه�#��E롭�]����of4�I�ڐu�ꉏɖi���j�/T����}�8�G��
��
8:��x��:��X�$����v���0'�Os?�f���<`D����N�d��S������������7��CaR�}�yNJY�6cw�ԠT��W�G8�%*������{���A��C웵���-=���ݱ��� 	��;����M��M��_'�$�#*ә�W�lBFu����W�gg�op(�2�ɋ�����d�T{"{�� �?��Z3oG�Ԫy���g�������8A�<����s�c~~^"������Zmε�&���"�.f�.3�l�O&��/[,_�<�Y[[k������b�E�wۛ4��=�j��F�ޖM��w��m�N-[[�z��'�G��?�^U���� b|��s�PHH�GO��5�%$JOwT!��?\�$Emz���44b|��>P����i�a�K"7iJ�؝W���Z�������!��*�F�����vuC�-d�%�����>�B=�M�%r"t�(��h7Q�4}������1���w!A�^>>-�T1M?~����Ew�'�/��MiMy�i���e^2�]����������S��R�b"_H"�haA���QDS��1v�7�r�*�#���;������$��M ��9�K��l
*�Ig�,ɯ�DȈH���o1��
�2�}O]���&���}csg�r��sN�N��nA�
��iee����w��Y�����y��$2d��ӷo���-#u�������S�hտn�;��]*+w��K��8�u&Ն1�3(y���/JG�u J.ojV�]����,��	S;j �FhI�b�^w�P��t&{�A�n
g�A��Iy���prpH8��Y^���Xʱ�����SCϬ�GQs�w���'x%A��Y���+�Ί�%A��A� ���2���I"��y߬h�-�ft ������}y�=aк{6����$7yy��P���75�x��h�XB�F��ga��Q�����A�T�ު�@�� k�@�ݶ��V�Os�Ϭ�_��)���]���N��@~Ƣ��)����I?�00����^�����ĈnM�H�8��	4��Qۯ��n�r>>�?/E��
T677�Qż?|v��zݷ,��_���#��x2m�Reט'�y�N�W�٫���._=�,�0�L���8�sjx�6����n���⪡�N`��K^��+���j����9�����z���_�ױ	�b$����.�>wr�̞<�9�����e����7�!{�z{��{/<])Ըn<���今6,�7�w�O�*f_��_��zF����g9�$������:Q��p $��c���m���� �ͽk��y�|([_��m�IP�ﶨ�Xw��R+<���n�߃��Ҧ���f
�s�F�: ��^^�,�~������̽L�;~����n���}V��ۇ���T�3�^ZZ�~���<��vaUg���I���M-ڸU�FO���{&o���u�De�'�oȢ;����ٿxQ�����ݕ���idm--���}�͒4Ņ����XT����2w*��������d������
�TZٛ���vNu��&>���@
5����Tc��dVm�+��5;9�V?�p7���Y0�v�y�S�˲�� ��&�~�8I�������&���ޠ���u4Z W���]���¥�m�/M�7�G1;3���;D_�N��ll�"���@�H���s������������8��if����1�KQVM�B�,�PK   �cW���/�� Z� /   images/d30bee40-a8c9-4828-86fc-eff82b5740c4.png��US� ��%�[pw� �5�;��ap� �	n��;���������}����˩���>�j*��(�(   ]^N�  �  �#!�'bh� �T�JI��KIQ��9[�:X �9i�jz�K�ct�B9�nyg`q�,�"	2�Rp����+p9$�)�-��_b)���k=�zCéy��0U�����M>���ô�Æ���;9 �I�Z>�`�^��\i�s`���1 ��Y�"��ҥ�[��#w�U׺�o�11�S� )����G.�+�9R�Z'v��.�@+�R52���x��t4N�X�i�1`{\$����S���4.G��?�b,Wg6������"�c����Y5�G���Ǝ�g�8��1�����̖�?G��kk*�K+��T~M�N�U�7�'�5.�<��>0^d�tx�V�J#��C��}�2��s��I�a}�o~1>sǞV��(~1IUQ������	j���c�����4�|}�t��v��t�X��`�p���r��{A=�%9���A�������k�
;����մ�����gH����*3�9fL�1@D�K9 N�s`)c?�9,�Q�	��l�cU.��!�/�<t	
_��va8�x"qBTֹ�h�3�䮛X]) S�������T�h��oO\�Ŏ��9�H?�d�a�L�&�xu��}dް�Xp�_>G��)��h�o�Mu�c$W�ZB���C`�9P��]�a���]D��f1�C̮��$��B����n)-�>5D�&��#�K쨑� �J��!�F.I��i"�������,�oF�~9B�%����8�C�Yu� Ef��`��-⹠�#9��.ow֑"' b��nյ�cBQ���}[P�D�$�
��h�%�֪u�C[Z��;s��Y�AQ�,��ٴ#�#:�g�Ѹ��B�&�tB~4�X��\�ߜ͙8�������~,�}Y�Fu�+L "���c=�|0a�E@9�v� fo���k�y�T[c�A[���rmd����޵�?��4+!ULA��<�/��EBWaEbE�;��-�L4���/DΔLC�jJ>,�O�[)r�aS�m���k%%$�����UZ�rE�����_���l����1��:+��F6�}�m��|*��h��eB��ͨ��˸�ͷDI�Oۚ�]sZ�MG��_�'J� KMP�ܓ�9�7�7Q藤F��ָ�^���ߘ��Z9�ѕ���j��'��b�1�r{��M�MM�M�B�N
�s�%���*�uY�YE�Mk�������b����He�6�fN�N<}�}C�Y�0��y�xÈi�㉽x��x�x�y�m��Ŗ$���O-�W7+��Z�E{F{ z%��N��.@�7�i�>�
0�ա����ht2��&�l���{A��E4+�,O�9��M��K��s�ڴ�;�������V�N]	�
1:9�'t���u����8kV�J~_S%k�2Bg��wSs�OKū����<3M��d���	��ꑳ���<���Rx��dsu+��O--�zMgY�?��4D�D��֙�+���Yfd�F��o�G��֩ʑS����-���!g(g�������K5�W2m�&�.P��Ѕۙ�/�)����������ƶȑ�~�v��_��i�#�p�s�M�����*��y��Ʌ����f�W.mN��v~d0�Eb�F�����u������k��#�+��iv��j�J��C@����ˆ ����z���'7�2P=0-P��5���-6&>u�	�ktq�_���eFޗ�������eT�TsIK�Wg��6�Y"�"e��anR��b��(/�l ��������H/�Yj���q��8�T��~��`�d���0��$��l ��V>�Y�w�w�Ֆ�m�����:&��cpx7�e���|B�
aY��칺�������'dNdD��+Iޮdi�݄!3�����o۬+Ԅ��Ha����V�3��)�����%?�Т~)�9]�[8Y��-�}����#�"B&����q�+u:H�d�.)���q�X��eAO_��ZEm0p;���0��{���}�� ����v�BQ3=*��Į���X"/:31;�8��~�n����7��6�{(ͱ
Mr2�9&^��&�x��o�4Tm˺�8�~�B��L]Bm����¾*H��Ṿq�����ӗ��o�s���OO!�ê��K^N.�:{P���]�2�o���~?��@7���K,':kb[��Xj�2t�t�H�W������Ӽ��+���_2@���Lk���ĕ���U����8ue#ť�� ���˯����v�vUK��i�u�S��'��'b3�Sy��]h�E��ʃ�b��`����1��4h��׃]l�Y��v}MF��^!���Dyp�q�_z[:$�����������sY�JU.�%»�jre������a�4}��������Y����0;�I����\8htu�<C�ȵ��ө��r.$�q�'w:W��Щiã{u���t���������w��)���Q��w1�K�}+қ�q��X�yCaF�&R*������f���������|����K�'�{
�g�|��4�#��֠@�٠��X�g�����	:ֵ	ߖ�vVvޗ�-����;?r�:[���/����O�O�}�Ke	3���2A��v��wW��D��~��A)H�����? ������ge�pY����W���yX6��<XJ.
��3���.��u:�IF�����^��w]P�CjAg� ū�����2�=u�~�^��?����  �����m|���v���q�?~��������������c\8�@���W��Tfz���I��>f���tn�X�7�sO����훠�e���APn�u��[�sT\3�s��e��s��R����o>x����?��?��?���A-��uz�I-8V�����M��U�*��/!�7/��?�B����Bsڇ*kB��S�����Bwo	�gG���6�R������C0L����/����8?��v����2��fjU�s���b���}YU�������_��3��I��`�0����fnE�,C���M�{Y�<#RSM~�����B�|��O�m�������bu����c;���x���>�[N�V���׃G볯���榰ѳOUsZ�>+���i����zn�4��F���fͮ��U��c�[7����S���y����M���RGQH���d�̱,�Ie�������ᶵ����szm������������%�����������c���A����}O���ŏ�KϚƫ��'����Z�U�p��j�P[c{s��1�y37U
>�G0Q^P�^�?�>X�(�>��V�֕h��*��!�&폹����O��ſ�K�k��tT��|����;��Ck��e<�Ҵu�A�SlF���-�����'�d$/�l���=�Z���ׁ�p�/Ϫ��ju���(jۯ/���έ��0(p� ���@��$!;�P"����^G�#w@I:gV?6!��"���_0rBFKK�`�R�e��h��+����O�p���D6$J���*�Yb�.L�vq���@X9��U��)h(bo��&�7�.���h���o��g'I �����W~�	���p������n�^�ˎ����xȅ�o;�GO��8�k��8�u"B�rC��]�o��t�A^�ܓ���e==�sXD̦�˭�G�q�o��Y`�����(��an�JiBi�~�n���-l�J1Z��'��шp�t;�@��m �R-E~Ҋ@������I]1��{2�Ñg���pB�(ٿa�+u����\�G�������_]�z*j�.ʙ�//����id|,~��X�/9�v*.����G��xױ�tC:��Qj��C���v��`Hq�Tc���8 �)�g�����X;��)9��������YzRl4N�֜&���x�t���_'���X1�!�ϟ�5gn�io�,�M�c[&b2�O W�ݬ_4��k��7�';f�s}���a�o�>�b��l�dnAW��WW�||��n7֢W��&Y�7[D�\t,�lf����ڻߺUI�H_��	M����k��͍�M;�R'��x� eV<�S1�V�׺����amE��tc[=o3&�OMIA-�s�$��,�W���?�$B^��o�5�*XH������ ��3��w�C-2
j��r#]��s�0�W�m hX�	F�'�}�]�M��U$0`+�
���l`Ϧ�W؃�	�#r�&k��En����_5�yfr�xx��Y��n����Luq5Zol,-�L� ��m����)m%�KuH��6*[_U^�F�Ñ�c�ֈ����r��E�s��s�R`�緍<w_@��ًd08�5��sp�@�V�� �8@)5����m0&�wJ6��{#��\�o�/}����9�ڝ;��n�{o���U]���(��)�d_[�&�҂��/�o�a	�m�0<�8�#��z�Y&���xW�{�ޒ�k��A����ԑ���d���R�=�����/p!v0Z�`�`�AGH-_"��H\F�pF��3��Q��d��}�ë���E�3�z�����̉�i���O�����A7� qVT��*���h�;���71�a��u����.ͽ9]'X7.Ҩ�,�sԱ!�]b�f���`v՝��Y�;~����xK��;2�@Dݠ��"�ډ'�[�Gdg�9�5#�QwZ:����#	g@���S0c=p��ƥ =�/��0�I�]]�@�/l�5-�~-,������%=aD���>3}*�#&�YYp��������X��GA�š,�1<r��K�n~a_Ȧhk�q}P���a	�^|��,�;����	j4+6z�r�~:��FG����>����}����yI'�Ŭ����}�[�rJ��4�Z���$�%.7*��P�H(T�r9	�Y�-���p����L;�&�-Ҫ0�.�5����ͯ�P���,'�>/�Opx�uHj���r����9��Žgh�-��*G|�������Rr�w�+��ɉ�����)�?���]5�1�F(�(�Tg}�$��/>�7t�'dx�|�_f#��~��ԅp�M1�����d#+E�f(ӬG�;[�@��@+?9��!�j�6��J֪�9_\��4Vl�TM�!ٗ+�[(�� �< �$����� ���@�[�.�њe~��}-�O_�`�&iN�|��x���� �+S�M��<>ᚙ�J9iF�;YY���0�F�J��.�e�Ss�t�L`����D؆z:hp
qZ[�����Yr���)��d2XI�TI�I��8815ƓY 	 �d+� u6l����s��ޞl�������%�~������f�@�~BRD�xw�\g�/�g�u���CӪ��m?Ӑb�1X���R׾�ݍ��YؼD��8�N e�����wtu9�	!  �fzT�֢nܕ�b2�\܃�kNGB�������	qu|�� ���):�����I�yX�a�͹����_�D{x%7�pV�,G�� �O�f���JɁ�o72��(��?��#�{*\��ϏHICZ7a`r��D�%�.���I#&�5}AуGgv�<����އ~������e�a]J�f���n�E{߇*��׉���(�����Bm�m����:AXs( �9Gv�-6g���7���q&�u�E�CqWk��Z=�pz��B�CHO�*wCm�s7��Gpn"X�[�F5���[�-;����pF�e�%gU��g[c"J��������Z�;���]�YN`Xr��	�l�^h�p�pt�ԧ�o����	�js{��πY��).�u�zv�o��P�I�~��=m�o���4X�:�o�T�[��W�B��Z��LΚ�ha0PS�Rp�I��7bv
��5�ʿ�@p�� ��r"��C�1�$44�)�涷Մ�ov~�?񈊞����`��/��U.��Ȅ�--Y񻄍��I2+�{rGF�K�W�G|�8���E[%��s�%T�6�(r�賟9�,_F޸X��<ja\�Ҁ��h�T *��@	�em�q8ԁb
�/�$����2�ef�O�O�>���"|�~�(�M[��緐��f��3�M���d!3��_���ȾfԌL����2�ly7'���u��� ������*�����68k�Q��]/�)�1pW[�i�/��ʻ�?2:.]wV�:�Y��H N�b;��Fh�t�м��5F?ZC
�_j>��� �6|��	��s���̄�i�j*V��q�H�:ʝF�nY����<�����+?[�|Ej����~�7�9��ax&"��<���k&4��v�x�����dO115#"2bn�w��u �t����{��8��l���:�yU �z?p�#aa���(K R:�VtLA쮤8�p�4�q`�ܺDm����`������J*=�xx�=��>��t66���B�94��N����w�S&|�9Y�]%��;�˯%�})vd�#�v��^�#��"��G�߳7ۣ��u����>����v,�����'�4��8���o�~�Px�G;�F5�[�K����z���4�K��b�Qc�:v�`58��x�rU~G��g�҂qdw�Nm�A����qX"4��`�W�m��� 8 (+{�T�%���&24�L,�J�J*\l_.���c��k�ڇW�J���'v��n����9��wN'�.08�H������{� �c�j���JQ�����V�Δv%�	m��,�=v��u-�py͟��R��/f�1���-K��W�@�Q1���㯜���4e
�gE�3�f-u�:���d�vڡM�����Ґ)�#&,#`Xu(he�@�qV��9��*�f�������!�%��}�<�gr6�E���6WA$�0ʁ��d��j��Jʮwk�a����0a�1L~�\�����`��Q� ĲA�n���G�����<Bp5��H�H
	 �r��U�v�z��8X�h^�,�m9��U=Q�0�ae��!d.��-[����	P+m(��ƶh`J��i\��m�x��ro��f6+�����ٺ�?~���|� Ks$����l���t��HP���3ݝy��^o�x�v��ǧ5��Bo<��oJҗ����< N��V�{�-V�M�6����1�5}?��$��rҖ�-���<�S��ݦ�~x��j�#�;��p�i��z��|p����V����
?,���Ԍ�N8a���uQGXD�NB�[h�x��ҞMV(������iSC1ҹ�?9dG�b��Z^��Q�?=�#�p�3��ȓ)��r8zn���1:��������K��\�^�<����U��y  ����A��{-�h�D��/��̐ڱ�N�o����CpT�H��܎Ћ��>�/E^]ܭj����.��S�x}l����i.nfj��Z_��U�'e�~;�����T�#M���А� `��"�#����b�UI�%Õr��+D��V
�[�o�� %�}�F���ź�KIӘE�FHl8��g�Q�W���I6
�mtyNӃ=�������5j��7tt-0��d����)����L�p����Z+�B�.5h���oPz�Q�Ų!�FyJ��ɦp�긣��ET*����
u�z8�	��m�3��:V-Bq��'|��4���}��R��-��nA�|[�Sd+cZ�YR��T�rT��b[]��Z�BXo�2��>�#5�)��pV�;Qs�S��t�ZEia!�Um|��I���{�g[�b���Z��t9{cZ���"�a���Cс�	 ����L(*:֝˹�����^B)}�+�G,�������V��߁�5�s�h�٤���'��"Ŝ=p�FA\V��Xw�/��[е�m�S�.�r�����pARq^rG^$[p���
�c����EG�O'G~�����;���r���T]�M��K9�hǻ�-��z��k�Fhq�˨*����~�KJ���7�_����$�-�	�K��	�F� ���&�4���Q�҉�{��쎟B�� ��Y׊��R
�o�����3�缝�e�ٲa�c��r\�u>y��~�#��㛻b��X=�B�-hol�5�u$�1vh�۝�������o��vT�Δfj��*y��@{T5M�O�O�鯰�r7w�JN��1���Ek�E��쯽��+�[{��)��$��+����h������0�f��I{���:�^<�J��L�~�Z���G�����(:�(׻���9�6�a��T��+��]���hϠ,�{� �<�p9$�Dˡ!�pzE�b�S�����z�&^�8�����o��N���߿�"�m�g!pCH��C�"�����&ЕylF@���2"�	���վ�y��<�	Ġ�&�?�;�Tm��t��c�;-UES��K�&��8� �@�;��#�N'���}�"R��CKV���h�"�6�����a�N%d�\x~�6�#��^n�tpR�z`:�a�C���n��X����f��N+��д��0��̀�� t4�b��eW�(�h=h�+�iX�`$"<n��[r� ~��[�^��Z�I�+�1:�kV���B�0��e��·�n^m~&r�G���
֥Ner\�s�W��Dl�p�|�!�fp߬Iq�z���Iw��a�2�!д3=���� a=Q93�Z4'sA=�e��0܊i~���Ȥ����np[>�rK�����a�J��M�|R*�E`� ~�ia��Jg�h�.� {Op� HٗA��a�C6Y%�`z`Q>��8��MM/����t���˞1�͎�l��u��گD���AI����z:h�J@؝�]�z�*^8:%ā�*$�`QN�k�_v�Cgr�ï����٤��{�6w� W%�ڬ��?fΟ:x�g��mW?�r�qf�i���i����%:}���ѝ��(0Q:�_�6:���y�%���������(��|;oo˪�V
�����ϒ�T��M+ϷԛS̥CtCP���}sޚ������I*��nu8>轧�}���#�?pX� \@B:G��w�:Y4�[��d^o�U��Y?�7�����u���I���y��ݽW�}����e�)R\�ꌹ,�\��"|q��S"?4������ڡ_㪂E�	Ot%N�[�� ��$-�V���B��=���ia�<sDv���Q�G���� `^Q:�Z��Pa+8�0`S��R����
��UH%&cИ�f)�ɴj�j�u��̿�f��E$��끲��\s�X���x-A#ղ6�7���F8]S�DWHt�;�� �ս-nk�)�Ԝ~^��%b�/|�!�Rt��D|1AF�z�~����PE[kk>O���`���Ւ؊��(#��u�l��ӓ��z��;*��6�(��Q� \�nX�u=��E���PZ��U����$m8�:���-x~�<����w� �ASض��x,&����ـ`�>`�fp%/��\蘊Ԟ�V����F�|�@u�4�d58�Ô�g٨mc�o��e,G��L�u>��<��V�P����t�I��8"�U�wj=�k��&�i����\����O�s.=>�����G1�K��2�Dq\ė�2$bv���I��`5��*�'���:�:��L>�� @�L.�=�"��y�4["��O!s�|��'X�� �A3������p�m����Ī��U���/�?w���W�����r!��\�뼐�H<��@u���\�qa�iD̶ڡc&,my���A��}
]�kA"y�̴Y%Y� ��5'�`�
x.9���s4yK�P�����L���N_��J���w�n��K����:Q����?�jP���Ѧ窭�X�Mnk~^����?��������]#cgYT\,�Т����ѱ��y���+�w��Sy=W���^d/�����ۏ�'E�3�g�O3�S�|	�3Ϻ��,�5:V%x�2xS@��!p	9ص���1H �M�J���Pe̔�V�e�'�9��9�,,��AJ�v���&#3��Qjy�E_�Չ�2>���`�F�����} y\�X��f���g�)VH���B�;|�mVm����͝�&��SlRc02�ez���-�J�9Vv�x�P/���6�R7�=H��쌊�gS|ggZ)���׺oe���g���!i ep�<'�o��[ ��`�j8��X"j0�2�!5�,[l��DB��^�r����%X�6o̒����л�A�-�y������Y�|zK�_o.�p�Ư2��d넧;��W#����*�H�$��je�e߲m�\���ص7�nߠ�w���
`��tS�w����Eτ������5�b��
~�w��5�i���Űb2P�w4�e�F �O.��LX#���� ����������6<�L�
�ow,A��B�#4��4�� cш+*3b|��O�h�i����	����c���o'�L �׸�݁.!��
�ώ�'ľ��k+����	�R�)�HP�JD�=?����������K�O���T�f�w�0�[��}녎rK�m���ūJ�%��l����:.�Ɏ~�}<�S���z�r޴�v���@W'ix��v�.���{޵_nA_RӾ�W���Ɩ��&O�����{a轿��Ä8���3i<���]��me�>�pP�Kq">�y%���_����wy�L�8�{�:޹��yu�ۧb�#4�x)����� P�Q)��Y��w�7��]���[�H��+���z���);�Ԯ�̚�#����J�%Sԇ��W�[�x<$&�j�a��#䁑���h�v"1�sQ[d÷�PC�^�P�n�BX��X�!��:��h;K��'ѷ֠��=�=�7\���}��wƤ�{��ʞ�G}s�����б�g3tF�_�V¦CE�!�-��`.����|Ū��P��\����ʱ���ĺa�#e�Jɗ}2a�L0�[p��C�Fr3���}UNLb���Φ��IgGg=�>9m�1���IРϮա�XK�D}�^"�=L5h`���� biWOhG��U��զ$�נl���_�6���A>�Yu/u�ꠓ��l��t������#�j���0VE����u&0��37�#�����Y cC]�-����t�9�I����}���W2�6�KB\�I��}:��R䇛S�#6RO�m�<�4)\E���͔9����ȏ�k���]���k��m�S�A�X�e�=>u/ 5�ah�i^*eAy�b��Yq��Uڿ�|����%@s�lD������;4F [=����E�1Y����J|�M��gEv�N�]����/�x	:�����W�X4���q��n𿍝�����Ӕ��:U�o���t�a�����?���7y�B��L�����I̢��]�q75s��X ���/��_O� �{M�Th��?�n�ݘ�߇�Od�z�_��-���7�b�H�� 0��=����i+x
�d����m$�aیe��hN:�H�h)��+��ʪt���ğ�fIȷo�ˤ�e����5�Պ6x��g�O�	&���V�;QM4�99
̨�Ϋ؈80c�.�U&Zt�wm�������;�bNJ!����f��Դ�� B�d��KD4�>�/١Z�*` X.Wզ�S��Ͼ�Xŉ,��i�a> �|.͹���ְ����Qʯ��,����+��gF��G��9Vb����e]&RY+l�<~CB�+bݮ�'���nǙ��ř�g�{�h��%"�&���\[J����I���.�D�M�gJ�IDৎ�L�"�G&��8B��-��\�P��b@S�.`wӊ�D�&�KHõ!%�ن]�*�c�����'-�lu+bww�E��U�V�!�-�A�EW"��&?{�x����Ռ	j�h�h���+���'$�F�r�QB+#�X���'@w����;�}w�6Afx�$��]8YY�a��QO�����P,vw�l�.�9R�b7'��K���Ӟ{���V�E�4�@� O����4=��3��)|��#O��cNN�-�"�fi9p�}b�>�i�y�g!�%�(|����3���=Z��ƥh��&�ɑ�.+KZߋ���
q��|���D���2�h"�ӣ{�_��F�~�����S0����<(S [a+%�����2��U�z�I���`�X�G�� ���1�:��L�\��^��>J	-@�i�
�U2_��y_٦�˚K� :���&)�J���������I��#:ԯۚ��>4����{F�Wm�?@�A�g��w��@+83E�Ɗ�0�&n�gG���	���6Vf�_��c�;��ho�T�Y���=t�z�ӡ���P�*��Ç1�Y|������)���T��,�-���F��͠�R�E��)+�D��x�*��}�v�|ߞU��\=�)���yÎ�w��k�{G��9N����6?����v�Q���AA���,�:�NB���,�L�]Pؘmg��4���TP�yc`?h�#e2��DS�r?��<�N�F�t���F-�:(��� u�t��jKT�����vw<s��/��߻�"��|���}��� ��҇�@/Q�9�3���z��P*� �ݧ�-�d��P�Z��a�R�])��0�}|��K�����H	��ƿu��<D6#~��*���#��Ū���
z�������R#u������^��LC#�U�S����~�����l��N!��Y�~x��>�Va_baa�?H��s��ǳccV�ЅȣǞ䩠{w���'��>܀#:�6��m��%�QS������[&Q�%��W�"�y�y��a��=T©�ѩ�`�e5X'���$� �>��Fq���0�ҳ�"op��58`��������*��2����Q�N=����t7	���\Ao��Q�
�(қ2�}	�"#oD6�_1,(���0Nv�� }=B[{��x,n�fb@JJxcn�m�ݰ�SG�f]A�g�E*�=����������p҈䵞��� L�+
A��L:�t�)��8e�B�� (��]fg��}�̔�hfzEmFuy��6�Ve�R�_1�,��OSsj�a�@lՇ,�o�5�g��S9kڂ]Y��0��B����X�>>�^��w�I����oJY�*�����6����N_�e��y޺��En�-��r>����n���̖E����U�D�w_��D�P|o� _D�nh_��y|���<5�Ji������!�7t-_O;;�e5(�@_�>���J�|����% � :��.�8M@�\��"������ja,���ڄ�����vT�*��&��o*�_�Mi����w���6�����^�q4`���"t?�b�<�ã u�m:��:�ѓT�T ��`�x����vv4;A_�}vSؿ�6�\\�%7��s��>Wr}1L�i�E�����&�ȍ�X�Е+��;�ƍa�ݧWԏ�*mh�UR��܍+~���%b�9�Ҥ�<���,�����T��,ZcuP���"ľގcO?����]�=�b��^pՆ�뿮���Wt4�Ns	�Q{T��?{e'U�H^��t`2��{��r�����fzT���D��hUm���3`i��jQ�v7����|��U��~_�� �y�������Xգ �;����s4 �k��⥄����������ӈ��ٴ��%z�4�Et��7l�O��p�n]bw�g��;_eMy�Ţ�9R��?l�Y|3i$ϝ1�.��r��q�4m�[�ʅ�����	��>xʁ�2��jo�X	��Ӻ�>)���P*���?53)���}FY�<�@��G��BF�s�p9����:d��1�[%�P[F��X��-��ך���C�uX���Ml�/�m�"BC�9�@��Yɒ aLO����E�R���}�HZ��?t�r��({2�y��\T�������� m_���q���}@����&=���Wk��2\Mަ���㓏'a�� [�=��[���;s��m��Ҵ���*p��s��a/S/<����B\��q:3��aMk���VVou���m½RB%���E�N��Å�>K,�Z%z�P���/���x(�����<k�};/�p���N�&�����*4,
���Ac$+f�5)�YG�Pn[�J2��t�F���A����6'�S��6���.���j�j܈IG�3���ʒ��Enc��Ot�gC~J���~.|���Np��C$�(��nG�0������u9ši
�.��my���u5yO��2������rul�,&���:�1uI�x���H�j�8J�붆6����Z`P��Af_Xr���98]U$�����o�`x:{�a���9C� �n��?T�iD�s�fʓ��!��yd��H7O�[e(������H>Հ�:�=mb��>s%ry��qݣna8$`��"MN~
'�tx��k"$Ǎ�x�n��8�E4�E?;<�s���&�p���E�0���='�η@��lH`��nn���E򪭗To6^����(������*��Kه{M9�Q%q�ȼ@���9��뀣[H��/]Í �{o�(�60F�w�0S������ㅦ�͑�W��i�gI�E�p�n��yA_K� �-��xW=�3��^�J^���R!#�\���R;����0�������"�H�g�B4�{�۳{��䢠q��E��8�E�cML���-s��6����~�2v��OWs<�ߨ������e�0����JH��5Ra���՚:�g��3��m���t)d�f���2'�����8W� {,� HH�`�̬��l��α�!W7n(7U�Z���L1<P�#�V��v�Y��e�e9<�j�^��A���y�B6��t6�E��
�R=#���1��;��o���3�"Iwh!V�}���_��x�C�q�m�Ex�p����#9`�.��"��F�`��?L����X�θ2MY<F/D�o�>���1��1���t1�����>�m����q��%\.����(�f��N�₆���~��ܦ�I" '�a��W�k��	iO4����3Q(@�	{ݼ4�el���c�ܦ� ��^w����[�ȕ�yZ���w�	���HԴ(���Iu�	NI*I�
PZo�R]kub�)W|f@с̉O�MTQ��%�s�ʇ�[ޫY�m3�Ŝ¤\��	����l��<����7�Yy:������j�N��~�ӓ�͵4	���C�8y����$�����;�����A��=�����ōx?���=����-����du�X�B�y����?֪&�=nӺm������f��_��M5�A��]P��~�A��G��%[]��Hi.yq���%�"��ȷТ� �;f��^��c�U+y13�_���5Ƽ��*���Z��V�,��a5�K
N�<��Vӎ5�7^�HWG&���>�%F���� �~J�f�wyP�!� B���R�H����]�taRF\�+w6`ఊh��໨yI��T��ZѬ�� ǘ��\j�.7xD\:srK��	X"x#�Bs?"*�x��.b�6Z�r�Oc�sD%#i�	������'^�t��xQC�B2	��x����%VD�Ab��X{p�L���Ԕ�R6ױa��.dvےChLj`��҅AR^QRi����p)\ό�9U����u	���G�����u�s&�lq�� qf*	(1w�pJ����!�M��T�$�~j�f8���T���Xc�hƢ���f�w{hڐs��1��OR)g
�Z��-�i.�u���$"�yS��Ɛ@�_�H�ŞnS�ƄB�&�c�f���2�r`qʍ��/�����?�v��Eh��C<u����a��Quv�݉KL����Z��a��P�M��!E����>��.K$ծ�F.o0�b59x�]�H�n�mb{H�1���<]�r�0�K��"�v�Mt�w߼���������2 �q^VO2ҍ�RƧ�������7K�|_t�{�#����!Ԃ��c�����.�4W�:� ��� 9��N�Ձr+]*N��yri��
N�:��Qq#
.$�ᝍ�Nή,Yd�E�g�!���=�Pq�K1=�ti�6��熀H���0֥��$��C��"������K�/�RO� S@��(f�  K��Dx�c�z}=\����4��5Y��T#�F3Y�mbb,ͨc������z:	d�jמw��,���Y	��6�P8��ѣ���r�AN��Bw9�H$�GH�z�m���tH����U�A�η���0&�r��o�%M؟��v�"�]sܲ�C�U&3��pcl��h�	W�(�7�K����&�200�p*�Z~e͘Ac�����ᜑ}�C~�%B��x���ԫyu��Y�S�Sa���ܪ���s'P��s!�mU��^�:���J�v�@�چ��i���z�D{~��P�pC ���Ȓ��P?�PZ����q�B���*�m�4���;U�Ǌ����i�V�5M�ѽ����T���,S��ړp�ٹȿ��f��=ը����DZ;or$}��w����w@�e��X �+�P�_�L�Y���+8������xm+���N���i�/�95��1rM�?:$˖�T��d�B�L��r-@k�t-[n���lZ3v�g5�����S�K�յ�N��险����ޡ	5#�fM�*�J�����( ��Yp����rlr&T~����<?2r�}ݏ^�xq�f}s���Ң����*�cv��N��� �.��,C�è@�~��p,d�_���]x#��h�~[T�u�^e�iq�h��߀@���u�B�k�� ����Ј��P9�)�	rV�λ�>���V��'}�W����?:2(���C��|.�x�7���&c�v�õYH����������5�t&�҇m�&7�ň'*�*�eD�,�ދ�.9�wp�^U�]I��K�����NˋjN9�������6�@ ��c��m��i���|+В�]�������8�z�f��(��6�1+�C��y������ߟ���C�����'�H��$�C��q!L��,ʹ�Y�FtU-���F�#�2y�sv��KAtiw�L��_�Y�b��^9����[oQ��D�r��Zt4wk�b h�u�ޭ
{b�e����#|^�du:7�r�P���DZ��n��GߠAH�ѪHa�����r��Ar�Tk�� i� �a5� �����|.�Y��Ω�=���n��~@����N��z\�]_\�ɛ(Z_��:p���۰(åX���sY�9ׇَwC��L��c��%���b����W���hֵ/�յO��~d������1�<׷�s��=�z1N�ғ��v�@�m�-�����},��{���O��º��}Wf��Xo�L ^h_Ϯ��4���s�yW�"�[�L:�	�9V	D�zq���P����1	�\/�����b�R�"'>15�z� ����T��jǟE��.9	�I["H����Vw��hw��pв*4�oϔٛP:�o�.K=��'�45H�r�mT�柛���ƉT�"\���S�Q,�e���9��M�U#�oʎ!���f�&#�0�Y{g찋��i���@�89�A���"	��?�7�0'r��5�������?zq!@m  �}�4�<����`@D��@�;��1kC���*T3�����&�mM�����n����i*6�ؽz�r��_���#��kf-ֱ�P��]L�l�0#S��j�:屶&�b��bB��:�p��F� 5�	�Ҭ��B��Ƚ[k�(`,�?�b�:	Vaaw<�X�pS�ʕ+�6B30ҳ��=��VK���P��>��';�>�E���5+cg�/b{��͘t�^�0@��2Qf��2��Y�u3[Uؒ���z�h��@�Z>�ܞV7��\���j��\���s��0\�Cc�5�����n!Lυ@+�m�\����U9��aO��(u���՛��{���=ۤ/�m�>{���_zq��K/�Mm�h�L�.���z�X��l��-L������j-�'u:V����ӭ��_��{WG��e��~��?�Ý��;��TU;A�/�tҋX��J,�츜�~TP�M��U/��)�[4�Wǡ�!Y>A�G�u(�ߨ���3��(�	2(ǍC�R婢���K�+,A	'�~$g�Q1w]z�^5b�)6�֌��6}�\_D��{����f]ןw�8	��.��o�-k���t���erh�����{�a�����]�=�`"���&��Qˇ�~59�m��^��^��q�+X�b���]u�˖BP����+$F�*���rzw�5�TO�j��M��O�]]CS�!�CLL���$}�n�Nni��E�D�[*��8�l��b0N�)f���U]v`���垚��r0�%���p�  ��D�f(��55�%X�}�ݪ�/���ZS
:�������ޥ�9ұ=��ݸ���q��Ņ5��ID���ؼB�#*2����#mN�7�X�� � \4��u�o���I[CM(l��q��CwܕF����}�u��m��H[lS�&��� �ꚇ<���Y��;������
�T0Gp��/τ�JЇk��r�M���.Sf��6�eKI�E�"2�2����yפq:��"���E�G
��U$���� O���"�2�X#��B��&�� �8/�H���4X�@-q�_�T�0�f9�V��>�������y�_�:?w�ڣ�;4�e2�:������0s��_I�ź�����3g���0�,.��'����/������ps[ Vs�[e ȵЦ�ǩ��&(LЍ��u��U_]�O'���ban���������g?����c7r�����]��Թw/�5ok*'��:&�H� 9�S�"_�|9֮��� ��4v��K�8��[��k�s��N����#���ɓ/{���$�fG/���Y2��$?�����̅��y��|��y���P	N�U
�J���CӢ���4 �;�c9x M��h��.u*X�����Ԃ�2iP��W�ޫU��|�L���0��昄���l��$�rS��v�B�����#�0���� ��Ҳ �A����-���u�;k�K�1��$tI���!�z)]ʘ�����nyt
�9�L1ދ��ՋWg5�,�œ��)�4�m�&�i���t���������o	��)8Y]�0[�*$o]�����{�ź !!%eb�-}]ʺ@цlD���	���3_�~�$ӏ!<q_�i���U6�@Gd�����
$ˁo�n���<���V�}m�?�oJ��U���䁽itp�
�z��#[e�86D(�ׇ���.g��8���� X:69�����!etNkP�bΰ��E�%���
@�FL��h�S�Q��� (��)+��	��gY���@� ֊���	�~���`.�a�x��t-�eNzl�NԵj���_�X��?�A��g����kg�"l�ư ��F�p��E둕�F�qr�S�\^��xy����:�Ǜ������������z}��ɩ+��4�.Y�@/�����@a�nd�叚͍���b�=u*mJq��c���w��#���{��������;�n(���O<��W��b�����C';�X�X�^�ƭ��nPQ�ОR��5����bi�r���e��t{��(r�+�)m5P��9[M�1��@&��z��!-^�@�i˰ �p��Y�s:.ՙf`��5��w�x/K�;��g��t%�hGw��A�C�R��,J0��z��l3��;\-��_W���.���~���߭��}��w��������+W�SC�oH�N�11H�qc\u?_S(�P	!:�X-9�����ѯ� � �J�d��^ W��e�^98��'�BtU�!�\��ظ������L�;���W%�S �*@�B��M9����@�K����I4����q��i~v�z)@��� ���Rd|�7WР�+ԴSW�M�]�{t��]�>7�l1�tbTsDc֣�u�&�X��\Xн"�G�Y�B�=
��Vaϡ)�ɗ�m��uX-1B0*�T�]ieiũ�| Ƹ��<�P�H�����s�q��=ڠ��F�2G�N�2����;J7F�u��X^ﳸ���H����c3Y�q�@�!Tيg�Ws�pd��fͤ�1�d�i�gf��?l�� ����s�'�rdm�g��ҳq�`��
��0e.x���v]a���J��Ԭ[S���M�c���~Td��̘7Ed�a����kЦR���
k���^�xׅ���Пnh�l��������կ���wv�ٿ�MBؗgW��mnJ<�F��[��Ȁ�[[���fkx���v�|:����8r������|�Y��çV~������K��S����������Y��U �充��_��^}3	��3��עm];�*��~fg�BN�M6�������,���Ԧ�yuo�������a�e���9��ےC��E��\#���+���8��a�[�����Ph(a
�[�.��|�t���t���ZT�;9Mv��zۡ�q�P�$lA�X��H%g�L�$r-�-�{U }E?a,]�>90 �-��:.ߛ	r�O�&��� ��J�._��hٙZ�匨��y��ŕ�:Ir�j�*� Xrw�B:h|�1��:9��uσ�L��{o�����43;�ώ��4oս��3���t�%靖�c�СC�J
�ș^�$�K�s�2�]^Msr�;	-Q���uC�c"����0R��u��J-=�ȣ֌�`�ˈtS[�FM4�!�]��bb�����!����T��.�mb`� պX%��M�T�����S{(�B���u�8ӼsQ ��f0]�z���u�
ѷ@���eؒG�!B�U�	ז�(��G�L�u�G/��@����C,��h�4�7U��9�s���4{��_'9Aǆ��x�N��F��:��C�/����#����t��c,xh\BA�D�i�����8�`#�fԵb�<ﳚ���]�_p��!9���-6O��ļnT,������H��F_X"�%�7`��`S%$��o�N�(h�����ϼtjߛ	�}��M��߰�1t`�>���Ƴ.�*Ҫ�R�gYi�P>�{k��nľf%j������zm�t[k[�\��z��z�:z��ܥ�?�����W_|���/����c/����=�5Ϝ��]�+��.IMH,�ey��A��0�p�+v�!y�n��&�푢�ȱ*��{��5��%@�KA7�;����.��pMN�`Y5 !�
A�5��QU�M1D�[q��) <��������9B\�1q�d�hX�1��O�:)Ჾ?}�Y4���1�(��% ��sx7�Ε,)�'v��!2��˸Z����juP�g?���H��+�p�E!��PKH`gPi��r7$�~��w�xG��G?am����L���A`}��ƦT�&�%9ܤ{��Y���k����>1}n^sO������
48�k�SH�G@qU�G�����2Kb�����ۗ����3��+�=�t�ݪ��e���#��cD�C>8��b'fu{U�0 �yhj�$2�z �-�E�ی <x�kl{)��sN��7���-�m�2�p��b}:� �T	�����vauU�"}��`"�ȨD�>"�&Р� ���+��d��F�a�*��ӛ 0a47�uȁ:�0��6�Tz�/ ǈ  ���Q5���`�(��ЗXBh�� N4i�/�{��y�#,u���͓Mh�gw�و��� U�
GP���:��<+;
�}�a�^�f\[X`�8�`������*$�s:�ԋ�.�����9�������S����m�{��w���/_��n]�ҕ���ͳ��_����^n�ru}���nÊ|m�(���
����\�E���( ��Ya�����`s��ٱ)�ܯm�v����ty���qG{��]_�¥��w^ݜy���w���G�?�y�܅����/�����R���I�������{�7�Kޗ�A��! i�Ԃ(�Eتg�H�4� I~/�6�P���}n��Խ�&�8]vt .^���6��FM٧��V 28#��������3�Q��R��Q0�U�Ē(\��eP�s\�����k!ޯ:;_���Sȭ�Μ9��^�p�@�;W��v�G����c���n�W[���c��iF�߄�6u~��%�!?|?�,5v��ջ�p�k�ȹYD�#T�lU ����4AZ���mͫ�Z� ��_[�2��Z ��x��쓘�k�:0b:>E
�)`�莾����*���9T0׻���m��B���o�٫�g��x�,Հسř�tE 
!�18�3�O�����I�ti �^a���؉q���Z��I}��3�
p
��oِ&��~t��I�L�&���� ���d�l�<=����Q�n��,�� u�4�\t�&�)`��qm6�O�1���4(0D�!�!�nB�͜D<LY�Ua�k���)�Ɵ��^Ը2["�d���˳�>���^��#�/ؾi��\HT���	����*i@S{��ƭfh�C��٭B�yJ�g�}�-/�EU�� |�wb�`�)�1��B?_ ��B�CH-�������[q�g�o���k䦘�Im>�?�*���}� qQ˥3xv	��xΜ�|�	��LP~���H0�`���b
�CO�r�;�xF�p� ����Ͼx��l���t�*KG�i]͎U#hKu�J8���[����i�Z]Z�������DOtO8�٥i튺����~�l�볏�|�q��~�ѳ������_fYZZZuy��ѡօK���]��/<{��^���/��k}w�M��C�.�q}�&C�#9;z9�G综��"�[ٕݫ���� zQe�@���ȠK��H��%���[HѸ��DÄ�/�n�]���^9]8%�';J�"Z�I9:�t�v�rh}��~#��! ��}"�$J���/�O�iT���H�Z��HM����U-�����^�i��q�)�%�)�(����n�����{t��n�)]���0�ːj�cg�V��|I iXί��7Ȁ�C�+#j�H��>�����Ki��ai�4
`Ɏ���}���<k [r��REZ��@sd�Bx.�h1�@Oy2�hbz���� ��YW������[�#%d��Vh��2� Y�
�"<�S���� �`�cj"t@-R��rB�~疛oI/>�\:������ �/;���Y6�FTǘQH��a�%�f,cM�l
1�j,�լh6$���x�)(�j��a���-
X�	�.�C�HE&]�lb�r������ƻ쬪�{�S�R�{����u85^ǣ��xW�I ���B��7tx�kI�^P\���� �M�W}ֆ$PG4Ӧ�C��l��#G��e������GR?�TU�1��EB�+��f���8�D�+�a����P���0�{��E���[@v�,�̋�Cb 8�72��[�!<��<4E����9B�6���nȎc#���S�>�G��~~�G���/�n��Ͻtf�?|�_s���w5}��m���'���P��(��߭�߂�+ ���Rc��T��K쌲�Y��ؐvt�[Z��n�觟�˟�L��mǧ�>�w�5�SF����։ڶ��陹��/^�������zsO�k|O��d���� ��j��UP�r��71��U��k!�p
y��f�m+䑛��Fm/�G�&�jȚ{
qy�J���q�uQ��.b)�ʢ��ށ@uJ hM�A�4���ё|���8~v�%4h��uEQ���Y��an�Vt�9�1�o��Κ�rD�����m��:<!G?R�3꠷������i��&�_�u�`�E8eP4�ژ��E��;8��r> �6a�q��M�kn��F�K�c7�<S;�P�����*��4.���^��ka�t�ԅꧾJ�o	��6:1�9��0�Ì:/����(dCas Nw'�;1!�e�\������c0 [b��*7�`�j��1,ئ܂�Ԑ�9wu�B��������P%����!L �J����K�|"s�7��8�2<O�c�l�y4�7sbì��h�^��,ӳAq�,%�ܚ��{�
����*�H^�bUz�74n��1�j�W��P���~O�<�8�p�N�����s�Ⱥ9�j�*���bߩ�f}U�D�N��c��}�{ҧ��P����κ���[N����t��e�ߓRާ9�����s�L(�[�d��q��% hvthɠrU��}#��w��Uq~}ܫ�C1ǝ$;�ݐV��. ��y�r����[Ͳ���	�[-(F+��C����ە�^���0SS�T�y���g���_���+������B��S_8���#z╙?��8ᢝ�h�	�������S)�Kw���z�X���j��;;]���E��F�9��ӶfqqV@H����������j/��Т��Š)jޑ����-��Ԋ��58���%� �j
���&��P��m��HD&)�A��a��Uy[���k�%��r���&rm���Br���h�A��� �ɉP���n�2T��Q��sreI�Bv�#�ͦBAJ�v�m�1�PMyU}���Qe�W`lP����)M�:��!���p=rN�>�.��e8s	8ӱ"<"����@�uK��#��R�ՄuPE�n�*F�������j�s�V�, �F
��a�
 ���X$ݶa�1���k�JӃ�"����;�Cwݞ�z� �<�=�E�V8X�`n�0;�����#P����f�r�NQ4��!c�0����Q[F�l��d¹Ѯ��R��[�@86:��t�����{��w���S< 7bu�"3��[�ǚ�քlҒ�V�E���b!��B��v0Sݺ~����=W�/���s�p��!�?SefFsJ��� ���M���t��8;K?��ֶ��*L8�1fR�Uf����0�!�ߖ>��f
O�H�����mVl�����
��N����4���.��l��i:ΨB�\�^�fk��!��C��u{�G���{�������<�������r9Z���|�'���`\� �>����P�wܮ�E+��f�B\<����d��b�=�^��YQ���@�l�Z�3N�s��f��0&`��lP�/��4F�W��'^�x�;��~}�G�#��?�'��f���o26�?�4��ǟ8�����詗�}{mp�N�bִP�����G���Z�y6ހw(}�X���)�5��r��[E���%�a��K�,!#i�H	��V=.4yZ���%���$,�&���f!�3�����"�ϩK�{ׄ͟7�;l��D%H�LU��͒��0 �M-��*T�ӭ����N�u��3`$X>��I��#�MιWkLNAj�H�k�f�,�d=ձw���a�v�vؤ6k���ظ���`���B`4 �F�@�M���h���qU��-��5���V5"�W$2ݡB0�b�&��BK�8i���8�
68�jEa4(�=����)��J��nK���+M˖2�`H�����G�gj<�똿��O؉q��xU��;�X�ʳ��a��L�
�-�w�
K�J�C!T��p���7t.����W%�������0g�*���T��R�]�>X��]>sN�D��N�c��)|6�N�>�fp����P7�y����׮^1���1H :a:�������b� �d�g:5?��F�
MY5�PtR$����p��;��M�kM�)�Z��6�j��{*+S�ѷ~٥q#��0#�6��'�ӽ^R��3ʜ���U"aX�V�X>3$ 5,�CB���Çһ��٧n�'MپG�}Rs����<M����o�`���H�H��]ߕ�x���_��N�Ȟ{4������\���10�^/`��/� �� �Z��n�� �C��Ue�e�b]���C'hh�z�^O�iM�D�
�D�z�y(|i�yLs]2�pK]$�<�~q�q��*H �������\���c7]��<���w?����}�C���=~�������Z��v}�5;7ףJ��Y�/mn���|���ϝ���k���&w��u��7��Hg�iS��R��Em^Ƈ`E��z��|���
����I�qy�v�n���3�I��V]��V��P���������ve��q �}����M����dQVl��4����ܪ	!�v{<�tp{R�go���oC]cqvb�@�5�aW�_�>f͌Ő,|�k�R���?�A��{�43��F�ێ�:;��SS|8�G��h;�$T��}����#��	-�	c�1��)��1��BȶbJH;v�\��y]�������_\�ty	R)�뱨[�G��'G�PkR�	��F���!�#骄��W�l�!՟+�r���v����ߚ&GG������@�,�ft\ q�@Ì����u1(4UȆ�
C�B!AtXb>.���Zz�q�'����!������ 4E�CU 0���uT������ �#��"m�����(Ao����F1r+��G��Se����6��/=�������'���~���/������c4�� ���#K0|&e�kT7�J̰_[�W��E9�TB��}6"TC��ǳ��>KU��Й75=#�<0O��L뺄�u�fkn�q�m��<d/ ܟּb<�~ �s
�ql@���SW�?��e���GD�K���ӫ
�1v�.�"S�Mڿ@1��*[����;��/��/x��]<{&=~<�sN��tt�y�7��Ok���ؕP+��
�m�؆ ���d�w�D3Ã5`-yV*@��5<���E?<�4�!�}kg������f��3�C������F=У��Aj]`N��P���t�ۆ6?C�#i�������S_x���/���-�/��412tq��{Y�9����_�z'ֶ���Ӂ���}�jh���z���#�$�k�	mh�ԡ���D�ʁpP���&( �Zi���ROR�OU���kI��שJwۢ|����C8��5i"�{G;"��m����+���C�Bq((*����wMo����r�G2
���
���o��D;��r-��a�X��q��íBYd-���m�[8M�O|��r�E;W��]� ��)8�7��ǽ��̈́$h�J�⊲�S����a@��~-R�?�,�*2']��3�tk��.**6��!W!�>��7xw��w��ܣ�e>|"���:k���+N�)$��g`�X|7$&}��5�4�b!	�j��.!�gD��ij��E�����+ 37�=w:���}����dﺄϑ^/!��:�ώ����ү�c8ɵ�p��38vv�%�Q�6$�: F�R���z\����)a=L#U�	˸E���w�}Pņ ���MM-a�:���/_��&�����ߚV�i��x<}�[ά;�����C�/�ȏ�����#?����F�3?�����E�#G���cH�N�-8�m�7Y�{�x��x���"�QsDv�w���;xPUR��v��_`��KEl�w� @U���_��@}v��"g����qL��[��[�G>��Qi�n��v���<ux[����fc,u�[�X��皀Q��306�Ω8�ɓ'U�aX!�=b�V�z@�$�x�4���j�K�ږt�9����b%���P��N�E]T���$JB,�� ����#�N�R��Q`���j����5�c����F�����
��i-���Xd͹w��+�Ω�Lm%�{t,6	�kZ'���|���0�59�n�=�|�Qe?^M���B����g��B�H `e_X#4}5٤wd�Ca�	i�&^��|�٫˭������JmyeY����>mV$$�JkN$jt�Q�:��^'ew�?��zV�=�hú(OZ^ot#͂е���"ւc$�H�|l��x�q�#W�_�B3�3���C�(Zv����{U�3���K����U-�v��?{{#��k�v�.MO�X	=��}��4,r�Ҥ� �]8Q� �%V�N�]ZP��H�eEK�jA�#�\���fP\0�q��:� �/����pֺ��%���Dz4U������^�h9��JA�-?f���%'ֽ�/�(|�0v@�uZ�F���������4������+�@v���e�N�;�I��.9����O_xQѓ�%���чK�+�k*[`��x��=���`�	�jQ��`�l] �
��(T�ۨ�6�����)���q�Ua��0�d[�Z�7&a��b�L������.�z���~]3�$�x�%���]L5Zq��E�� �%��:9�}�t�=b�v��4�THqD�[N=�E�tB�k���Ŵg`8���黾�}� ��!]�~?�J�����k�腆^��6#�J���6��e�>��O�6�L�qe���Z?�����eS�aCs�2�C�أp4Yd[ꃖ�����:�������O�TZ@޻oOz�;H�z���=\!m>�˦�����Q���i�� �L�Z�RqC2g��Tl�@tՇbp�;�p�E�n[s�3�(���X��e�>U����U��=`ʤ��D��}#iVlO��-�-�_�L�{�i.~���(ݕ~��~>�]��z�[��a�UϘ#�$5T���Yj��㽺�a*u˾+*�@B����J����P@����г��u��1Ӝ��<E碤�;v�q�7�<���s 3��\e7j?����M�r[4����ξ��eK!C4H	81���X��.k��jy��e38D�����w+���
���fCыSr'��@� +��C>G�H�"!��}����^��ya����L���E��>UhF�H� ��P�충�B��.�DMi���E�"�#�^;n QU�gE�2炄�iȜ�E�:�j�ǖ���X������g�B��ٖSǗ�P�`p&�ۡ�{�q�B �b���Ҏ[�ƃ�ɠ01���؀��%�h�9%V�N�^ՠ�Q��bǉ����t;r,��K��{����Mkr@�I��U��Bs�!<�0r4��I��~{�h��-?ܣ�
b�X!&uF֍4m��uL
�c<�w3U���3��y'��svZ7�
 �<R�`���&�T�|���E��c�P� W��a.IɆ��r//9�m�GCW�W��2FT$tb�;]Z��{�x�B�b�ݿ��i�����8�#��7Zp�۟hr�O����������N�jc
�mi<z�:�g�L���!�	l��k,��@8�K�<�P*Y}.PIͪN�	1v8{ݛ��%�:>�%��M y�,p<59��7�g>���#{'�J�2�X�M�f�3�M��9��@V U��}�7ڒݩ15,�熼0pKR�́/Bl��X�O�n��MR��w]����V��l�;�i��P�ĸ�i��yN/��y~/S� �K���w��xK��ŕF����*}�S�R�	���)h�A��c]``�& Ê�:F�\x]@�j
�\��i��g_Nt�Kk�N�"��=�&[�����7?���g�b�ٺ�P����s9��W26v��
c���ye�:�#z��n�_�k��$����d��i�ƌ���
�Q�b�����釼	����|��b��nl�x��2����??���y�����o�V�����{/ �;_-��Z��+����E�aBX�nm�`�i)��8�/g��"�$c��=j!�p���.�n�m�(bs�WHyMC8?t1>����]�'��ӭ�#������I��c����Uw�!jȁEJ>�M����)�]� �4�u}�
S���܄ T���rP��#
mP�fa���Y38�#���gt@0`��I�p:q�z5���w��G����\Y��i1�7���P��>ir�q�r�b�?�}������,ׄ�c  ����\ǖ��9u�:��}�^��Ħ]�9��Y�#��#�˂e��|~Ga&*�l�س3-\&4�ݵƆ������bm����;Q&d�x�b���>�������7�QZYh.�Kߠ��(g�/�G7�����t*�l2j!Q`@� Ӳ�#��S��^B[:6��v���(j���&�F�} f4w�/%��w�l:]���ۤ� R�歃�w���0c��������A�Ic@}*� �0�#mK�#ѿ ���u�z���N�G����QL���^�/��M�$<�-����Fu\���U���316,����;��)����lBD�����tTz��Ӣ����?�>�ɏ��S	
6�\�L��B�� �QK	^�ƽM�'�L ��Xy�����+:<�]
�څo��*9����VʆjfQ���t�ٞ�^?�̎����Y��τ�d�pi^*ɀ���b����#�5Bˇ�lS5t���P8���Z��	������[��`��nly�ՒC�a�[���A���f���倝׻��R<�;Y�p�|�ز[N�L"hkJ��f��7��� S��K���X�U�5�q��r�0Idn�c�y{���GU�%~X���-��8�馐��:ęjERA_ b��� d����s��zA>x���Y̨��ҏ�M��z;UdN�	���X����A��eǣ��K���R}���p�8�9���hx\���k�I�%ݚݤ[�Ȧ��I��9��֨�ZOVZ��Bf�<�v�q?ts�4��l�����y���i��ElN���zE�����ލ��Y�T���@`ѕ�->W�E4%�#(<�����;��u����l���q����9�9����	4�]��;��[bs@eS
����%6^iu��#!��N��^�@�}[ N)����]I��@ˉ	[��iga�,���$���c�-��"��P�pC�7�
0�!�o����fz�;ߙ^y�e^��, Y�g��S8x~i͟!�kR�9��4f�}��J�M'z&X3�l�
�~�7ؕ��W�Ƚ����k%T��.y��h��j������[k�n�1D�E���*�`K �B���*�wHn�>{D���[
�1v��`t�[b~�._��a�nI`�{c�cG��(��x��q;�*����|�Nic0�q �![�HO�K	�I�@�'p��Jr����*�S�T��:6��C]A�Va�j��F�.�X6a~����:���g�}�h[!8��"zD@�((�c�JB���ࣜ>�ETscΡ|��a��n`�x�[��(	-tR��H��ubb�U&^���o��Ui�o�_����@�Y9Z�W� ��	ƁE}YRT��U�R]�(�n#O��$h.efh׫�&�+2��1�|�j����S�0 IH���/�,�\C�
�[ab�u#J��AP��Y_	�H\�
��n \�cO�p_C�+�{�= �Hq�����PX�;�M*���ZG�Цt���Bg~��qũ��Td��g����0 �r�M5�DD�����Q�ٴ*��C�K�(Ш
F��@�)�+�}c]�D�;�ޏ`�����j��F��p�a��ơ.P�!;8=Z�min5��� ݒ��k��Xֽ����n�д���f���}�I��ݷBH�
ڮ/�����~^�O>��3lV6�R��tVs�c�=�
��J˲��y	ʛ��(F��9���ngGV�;�H�B����s-Oy�7rO��+��ԔTP�¬�����9�9�p!��t�^��9��QAS��W��{������v��X-TY\ ���KU�E���k4��(��(H�z�'m��XƁ}ҙgt-l(�R�#��F��~�S�%����Q��4x��y���[o�5�^�v�i�y}?41(���A�*�y�D�$-�E��F4�������WU-}%�}�-�c?�yN "|�%@��z�E�hj�Q������2u�^(e����j[�c��L�U�9��u��Ɲf����Dk8�B5�X'�>�M���r]2�����~2�i�b�Cm)�3F�\N�Gn��9����,�fэ��.��_��\����r( ��L���'�;';0����:���[9735~h_���9u4�Ĺ�|8��_�f�����I�����d1h�;|X��g��q	)������i����y2�^:yF�W#�w��2rX(�q�,��	���>-p�C� U@����&V$�)�J"v߱������\�h$�T]9���hT4Qѝ���v�P�M�����ٻ���	fڥK�)�,5sQ�O��qF̎mRlqbXH��C�0�ZC�~i4?��f�uV�BϙE�	��}JQ�`��� �����hPz�����%F!��=F�B;���Z+-�{!��G��HN���f)�,�j�G�Ύ�GST��T��˺:g������p��h{!' {��ձF^�C�3}e:X���zo�[Il.��P���+�J_C�x]�Ϩ�)#����}>��گ{XT��`o�B��:.���zY���E�D�X��QhJ�X~��b����'�dv�veM��h�� ��=-�\ �����:����Ջ��2тD��>�o�8�,V�l��V �[���X"|ZS�.	{Ra ���b��w̯FK����E�(����^fP!�G>�Y�T�)���c��^kҢ��_(��P����,ρF� ��B���/C
ա�!4��� m\a��jt[�q����׻G�	�5��f�N�p�rR=��P�˧^I�/��>���N�������a*�ܰ��Bx$i�%Hff�M"�Z@lN%!K���yC�َR���^��"A���z6�W�n6ȜU!O���zl&X�Fp$�nj�p0m��l${t�x +���C�\iz�����6�Uڿ�6���%]���X,cc`Pz'/�:.���jَd��z�X���i=\�8(:-z�`�����Qv���ľ�K_�3?�b��8��x��xe ���gr�_��o��~�NO�oC��[S���b�~��φ*�6�ׄ�dKd<�
�\X�0r�����#ZMW�5��F�E��3�`bKء�|��6;�j�=j���ʙ�RR;�4��������t��iD�r��I�J횮Y�4 eX�7��H�s-9�%u�v%[3�g�~���\������F9$�ա,�.e��G�P`�N��G��um����vP�4�������P	Z�B�F7�D���!���"0��Cg2+��sl�tc]�C�
֜V�v����BX{@��
���K0U�:~}C-h��r;��t��R���řn�@_-�X 4@�Js�{�17P=th_ԩ�(��}�۰�]-N_L���)>��;ӿ�W?����ȭ7��'�����g���c����n�Mb���W����~�sk���H�0�Jc�!��/�x�޷���.�)�R��^ENjQN|D�έ֪�?����	9������/�ZtK�Ʊ�nN�}�{�3�>#��B|�=��r	f]��Wl^=�x.��.��S���j0"�`�X��å�CU�yA�ې0VB��ѯ�ބ�O� ���8b<�oT�R�w��DH���5�,��Y!קIbM�dW~�:|D=�&�?�ph�����ds�p��t{b�t�>��e�����C�.��N���-1���ZP�[���ҽ�1@��3��W�L�%��q{���z�"�I�ް��E-"���6I��\e��	�	���K�>ܣ���wަ>{W�yղSA��=jƫg��6/��0I'��
6�)u>K�}��ҹ��������^���4�T�u�g6�޺Fo3��Z�!�\E���6( ��:�ڠN]i�".���F����x�}�� h��(�ֻw����Ϙ�@���(�3(����;1eCF@�d�@�*��ЎJ(4s��������:�g�P���pگ]�ჇҔ� ��A|K3O0#Y����kYRk*a�tb���*�J(��E��ǟ4a�FH]F�����RD�4��n��M]�95����S��L�K)�aѯJ4���]�6x����Wt�,J�k_���}��Tm*%�n�t)�4 �=	u�I��룏�P�8� |��\����B� x�~&pJr��V��ϝ9�{YO���S�6i�;륅(r������΁�\���=�r�83eI�αp�##��������P!�5e��f��8T��fB�a�=.� {l��:sE�PHK�������O�
ǜ>uQz��t)��Z�VbU��ȳg��s��O�����l��?���;�Eao��&eK�N�
=-̥�g.lq�Wԏ�:�11M�.N��Z]S8S��Bt��9b��q��iR��Qm?4�hR�o��؈�P��9��4�=�"�S����H0��i�M
\�m(��*��²6�Y!�%$yYU�����^	ꕄ �2/'���z/}9ds�շ��	9�t�U�L9���m��/�=Q�0V�b=[ڌ�h�VUoHa�>��}�d��ҸB�=�I��C#b�$���;���	ٗ.MO�g$=���\�/ϧ�E �4z�>����~���vl�\b ���1�e�:֣^�l��kda기pu�n-�8�<��A������!{Ϩ��d:02�f4ޫ�
e�l°��t�Z(�Zm"/`��N�l�;����E��d���� g 5�z�a���5��[E��6/�z�>?�\D��[��� ���7,��Ǘ���r���bވP:���p���rwx��h��Q��#.�0b�F-vBQz��lsUU�U_�S���u"��-�K_u�A/�dU�_�@C�gT���B�w�P��޻����f�M���-�d']�4m�r��-�v
΍�+�t����2��I�:��`2x��㢯SM;�&Y`�nX���K�d^�t���wɡ8Ӱ��nBB���{C�u��]w�)0�ߡ��.�/�2�A�Q:�~L�k����8 ���[^ZM���:m�nxV����r��K��F�J'r�a"�����	�
�d��3ϼ�z�Ś��MKk3>��@�m�S�e���h����h$�}�b����h��:�S���M_��Uꢎ��f9�G%Խ��;��
ƅs� =v,-�Yx�;НJ?�o~A�ߢA]��]~ŀuB�=��p����ӓ�=i������L���#�>m}՘��q�(�p�4#����cj9|p��Ƣp�2�>��OHܮ�Ld+"���#5{fTaN��������/��
s�.�|��~0���gĨ��kr9]�f�P�=#�R>e��!E��;Op� �7h�ک{�O]]ivA���ae]Q��܅�tN)���Ǐ
�H#4��ZLoem1oǾ��t��^����(=����E9�p�knf���H����`��O��X@� �p�0k�#*k1��Ź�E�a�-��+��vҾã
U��[WAL�^"ʔ,����cK�c���H�g��/h�#�G�<7��Ph�������@��A��OD�K������0��D�^ �na��:���֠��1�5r�*���ޢ���&�6���������#�{%tJC�H�<�Z	������D�ȶ�r�4C�E�#�lT�Hk���=K�k�ֹh�����r��p壿�,P@�F<@�gAU�d��Bp_Ʊ_��ˡ��;�, �d]�f��Iņ�q�j�FqCv�0A�/H�7
�,k�S��_�?�wT���	C*����D�������Ϲ�z���W���Tz�v�6~`���4�����3j��k��t�X��'o9�:6{���%-����s�������EU�~��e1H7Yw�͏�8�p�L��{:�"�,�02�����4���~����s���R�ȣ��tn�ً>�1tQ@��^vcО��t,]����M���߸�w�r�O<��Ğ#i�7|cz��g�g?�i�3�^y�q�#��t��K�������5��ܼx�T�]ɬ0�=#\��yF�����B@�鲪2�t�tD�L�������ω�9cVbJ�Y��G��/�w:�!�c��^��s/������t��=�2�����f���y��xN��}D��ų���}Ea�i�/�A����R�d��������О��r�Mi����w�!1�z���B�U�>���d�x洳�p����E��MX\�C=؃�n�%�& H��9�6����^v��;n�-=��/:����':�%�)���L�n���˳��|N��a�����/�1O�
����3k����f�&^��"�C�����l$H�Ǟ�<��Э�{�=i���mب�)wl�pZ�|:���K��t%M(kk|r��g�{�!��=궮�K�#���i�BGp����_5�Tn`c����^���A=?bFHP���͇��ҵ��ɢ.fߖ�[1/��"/�~A��A�N�鬧[�H�|����
��.�
�c_���
dV!@�"���PԪ� yV��1�.����iI�NՉ�;��Wl��7����~��P���0�a_O���^��o~2���s*Cp ��_��tEl�O��_�5ϊ�����5�E�{�	��b��l�h� �p]n�C=0�I#���%� ��>;�^1�N���3��V���md��n`���S�Tw�U;34���5/��
��G��i���5?�o��'S�|u= b��b�9K�
�� !�"���ҀH,�t
$�@���-���E��&h$�j
�I��"6��wh��u(Ty^��KD[v���oI�	� ��$<ݯŐ��+�O�a��{q^�刾�;����R<N��u�����=��x�&�b�Ω�����E�>,�1�rp���M��=�,��
q�X�3�+xS���<:��?�ԓi��@���ǟ��q�^ph뀴)�NZru1$'t��% a�}��z<--	<������$��F���*�'i��Y�.�M�4&�O�u�E"�[��_T��lE��K�EM��7J_��w� J}^���M��)ܢ�0N	��ē\�	� M��(d��4�N9��Ys������{���B}���뜯�������ޔ���ߓ����#E/=�����KgӃ�zH�t:=��z�	��,���|L�����Oֶh���?>6��҂f��#��^z�Lz�����{�I�&) Im@L�зʾ�� w]�gK"�=���8}����:A\oKs��ԁ�'����Fk���M�y�"�*6���oV�W�ןx�	����u�l��E���z�g��5V��ٯy�{ҷ��o���!fQ��=w�cG�X�{I`��[�������Yb��@�P�r�T�Am�W�bH�H�t��+�/
|_����y��&ѵ X������{U�u��%e�Ix|e;�����ྃ���~�����z Ι�jl+P��x(�T�|QdZ����X� 6(�9��Ԁ6{Լ������d�� ��l)L!�:J�k�k��Z�s+�,V@cq]�IkG��{S���7L�����A��][���7���tif%�z�X��_������MiN�8�7���̃>�G.'K���zk")��^]fCKZw����%�ޛ�'�笣s�X���G�/g�z�|����x��@���<����?sq���к}N��0�X� ��`gۭ�����X���k����
Դ��J���u��3 +�[2,���X,*� {)6C �-X �C�'�'W��J��)����	�
�����f�mA(uSD�;kI��H�GT�b� �!`�*�Ǌ�-�0 X��[p�O�$�J��q�|�^�/��iPo���d����Pz3�\!��܀վJs����B#B��S�-�T�L97�|��
���Թ��[n5�N�����51���̬��ȴ�q�Ȱ8�U7s�"�%SL��$ȥ��Rck�g [��sCL�\^Ĥ5�	i��&��p:�>��1�'�h���U��qF�����N�O��.�� RJ@��t~�{�������(���'u]׃͇�A���$1�£�O�M8�= M�!l
�a@
��pP��4X�;�R E�h��~��#bY:�A&G��hs��ü��d	*�$�̈́X,� ���y[TH���Ɗs2g��% 
�}2oI�� ��ӽ�48�h&.!3�}L�1�E���Ze6�c�Ӣ������ �5 ]ծ�ܫY(��W���*��XX�1'��r����W0S
�!���(�,�h�0����#-�΂ަ�cQO�63���h�*։g�J�$,�=��Ç�:;�)�Af�������~�5)��6�������F��-x.�A���(�U��֔	�-��.��>e�W=�K
�]R�փ�'�50�����pz��l;v{ZQ�vM=�ԯ�W �=�JenlS�T�K�7n	�4:��LN��|HSE&b��6S��T�-(�"B�h�A�.�G�\��l���~����w��W߼��/Y`�/�"-P��V=JJ��nzU
�I������5�X$���N�H�]'���!� j���G��q��Wquj��?ґ������ήyJU{7��j(KpP�Z8K�}�C�IB��]�WBM�	@�{Se��:r�z��'c����h9�ye��j�cG:�P���j�Cs���E�Ľ��㡗�8�4m�USC����*�=t=� 5 (�;]�G��ͅs��TwF �].Α1bf��d��%��>�R9$����*��3���X-�
sىj���^`by�,����.07����G�u]8+z]�k��߇4M����5��P�5��@���&��Vz2�g����d���q)�&mz @aCYt��~9:@��3���2���bAp|� hB�3/�
��>����Y�V4�Ԉ!(D�B�W4PfJ䬸���H�<*�ɹ&'��"��ӂ�H��r����x�{���\fI���!���U/�<'�,'�y��]��͙�*HO��
�ҏJ8Y�9�{�-�<[��.Q6s����+�1"��Rr�l�"��%���w!�F #6K�_�a5�j��u�;����=D]�R󆐧�kc�,�HB��ss邴L�c��X
⹠�<E�E�Q�s\�)�rN���Đr�%�N@+E4؉��g�j�T�����E��zT!_����/���3x�-7y�_��r2bn/=ۢ�a3�ߜH�x�8���$s�RS�uv��w�s�ΦǵY |`J"k={�A1����0X=�=H��"�Z��� 5�Q�Blܧ~i�-������³���uI��ģt��d36'nz���d�u�=��(�s"�$E��u��%���o��nh����5�Ru=��SHVC�u�q�Y��P;�b�z���\�z=��n����k��:vCi0G�u�U,��s5�pL,Ξ�b<7;�n��f�E��iр��'�o��(��B[
���84�����/j� ���^br"B#cM	;�U�[b �  3N[6�D������j���M�N��jĹ&N������u�5 �Zd��ڽnlj��v�8V���b���%�?(x�Seg�u�z<UW�~��j�p~*2�^����k��rVїL�t��`g��Dqj�Ú����s��C������%q��(x^�*o*M��
�/ؤ7��)�77��@�_!A��4d�K�ӗ�h2���;�
z��jΰ.�۬a��6�+T6n�gB>���:2�)2�65\��N�*I/8.��QR!�|d��~p�0^+�WUÈZ38������cӓO|1���,�	]�4�#zb�Rd�E��q8kw���n@�ٶ��r��|�A��amqO���唙� B 5�{�5�b��I@��۹��k��3�g������و\��nXlд�ܑ5$[�9�֘qm�AF&�}U�Y�ߙ0Y'�k��V���3�ƥ�5��c���y���^_08�����F�>��%���c� �\7��;��.�#��( )J7Q��f�.������H���<?��ۯЩ2��i�;�7휺���J������Q��6�k�Ц������w?���z�K�2�6kß�=H�H�Ɩ�	�S8K6��P+�_iB8�En��Nھ�>�mK��7�I�!�Q>����#�]�@(@��=HdAٵ���J
;���/����z- ��D�e͐�	�U'Q��SL��ڑi7��L2���[>$'ؗ�y�Q��A��X�q �ä́�`Q\��d���珤WG5ޖ�a���������$`ҙZ��DNH[�B��V�Q̉B���a^�Z2cƂ���s����%�:}�;yt( *v�,�d��&{x���C	9B(-�2�U�F��>id�h��u�}��1' �� �Ь*d�]1eq�>�#��ġ�f�a�wT���'�	$��qЄW`��,���Z�G���7���ȱ	�^��ΰ5��`\�b��Þ,�A c��sƑ!� B�(s������CA�fg� �)I�
�ܙBUצ��D��=��l�������� e|希@����A��6�bh�{EY�̗��G�&�K�R�>v�(2n�έc �"+}Γ0�YR���ӿC��z:�(vP���ؒl  S����y`��f`Ђ�3;S=�9k���w�A0��ha�x~�!<�k�S�٦�X��J��mA�����u�6��L4 �eF�7���y݇�m
T���f�yX!69�dZ�w����?�ĵҎ�1䙀�@�M������6�>��������#?��Nec>��S����騴Y���`�$��iG$`��y��jp��Vm���WS=��{%�oJ�7�.�xg׺Z�4������1؀RQ������d�$����҉ae�a���7H���x���?tCc���ʊic磇hQ'�r(��H�%&O��x�Bȷ#�u�+3>�l^\�7�&s�����7��W�>9���w3ͯ��X�̈́��[�ܜ�������`Q� -���E��y3+��,�T��  p�cڱ���n�q���08ZO.�c�G,vktt�U�-��s�\�8ֲ�3�np����b�~��m�3�d{];� c��"���'c
_紨�j�A�;X�i�1qr:|o�O_�<�n�N���	sPtܫ[R躩��#ॶ��q�f� v�d�P�'�;y*�g
j Y��a�4+�Ыv�W�/�X �F��?)��+*�R���+'��������x�2�F�궉5g0R�S�0���/�̎R�N�ת�UP}0y����̬����U�!��9�j �K	[��+V�-j4�C��9���#����w '�^�!�M��q�{�h�mL���"�\���bg~�+�]tXp߯q> �μ��y��īR}��a��* �"�����5�r|7�����j	�2 �*�� d�L]*2�(�9�{��WWdI-W�{L�o�0�:6v�=���]��N��p2��Q����n�c@u9���]~�=�=�닁�d�	�ӭ�R�{.3/XS��X�U�h�O�&N�?��:#P��c�Z#�*��ܓ���V��ꏤ�nR�Z�^����������ߦ����tǝ7�����?}����G?�x���KE8�K7�h"�������9�Q��VsK�dӅ	�!��V�pA76b
�G����	$@��+�iS�±cǵ��*��x��M����3�^㕙�b^/t�+�8�6V�4p�m ���jw^���+��c�#vY=���P��agG؁c�T>Ο1+�F�솾_�BgQ"�%��?��MJ8�4#*��3���tt�'�=l�Q7��iA�,B�葚�G�Z�?����Q�/�!���\�J\K]L��������/�+Ph�B�	¢>! ��o��@��GE��ﷃ4��=�^P�'H���6��K�$v�f��w�jnݑ��� �S��\4��e�_,0�}#�� T?!0$��rxF��,�N�x�8Yvv�hR(9 ͔� ���$���,�Q\]�;h�0!(������"�=�e��0ЉƵnJ* [��D��J��s�� Pv��JC���*�n�j{Q9F(jOMN��q��z�|�"d@+�\\�6���95{W]3����A �h�g#�	q�Ց-�h��]�K`�hx*�K���ߖ�Դ~�V*� ��|g��+��QX��#�+𰪐@��I���_�5,篪�E��xƢ��������S��%�ı���9L]��-�mk^Q7,6��B(���(�#(��ϛ�̦�d� ��,n��4�k�1��CL}�=w�.�*z���1Ӝ��ZWVY?���--�)�S5��Lz�R�隵�.�|6�\:�nW�����?��u�Bjz��~,uJ5e�R��Ǜ�6��P�V��c���ּ����zMO�����n`l���ŮhH���[S[�!	�P�����E���z��k]J���g���Z�͋�w�U/���$�Ź��+��� ��+fح�||��F��g?����A��x�t�
H�����������u���ɱ�@�� 
���P�&��#�w�-��:���v�,�#����ET�p0-���x���]��+��A���z�+'S�;N��@�G��7������ٹh�\u;u��@}��)�������8 �1˃�z��~�M��N��2��Զ3mZ�XlQ�~�����A�
Y�*V��XTڥҰ�V�ɚA�c��]�X� Ж�{t3V�	���o�Oq /�J4��热a�Xo�{��Cv��¯u(g����fe;��`Ć��p��ꡕ�>�$����ju��^ )Y[��ҍ��U�ul;4H+4Q���|�!�Lc��ap͜ �	���������!?�=�3b��J� ��Y�=, ҂�zc�D-��
���Ǣ7�5��f"օ`� ��(�K�M7f��q�~���C����Y��<0��c"��7@�P�x1�
�m�S����W��k��䚂��S�j�bv5� �lx�n�!|�W���	T�q�/M����Z����	������2��z-�l�����c�k����CN���������/�L��o�]��u	��u�G=(h�K���"@�7�?�&]����<�dW�9�~ۊY��J�@A78�0�0r�������i���.,X,t���Z�a�|���ko�៵H�]�N0Cw`�������^	v��r�,�>�#�G�
����y�s*�����*�\M�k�A�׊���y���-�=/�i���H��=! I]Ǧx\�?��ԎI�w�R}�H�IKa40�:��]@�ԘZH��n>3`>2�B 	c;B�#Q��O�\*�G �:Cs'kl������gsp�B �
�Q��{�SޡFgm�h�ն�v�| '����3���}�Ҷّ�N��q���A9<Q1����_.�� ��k����>��b�pr�8i�� ��{:��񘹪X9dj� b�]dvˬA ��u-���GpK�,�������� %w��V�����ED�ss������O����~��p�\E��z��� ���sP1u�^��E�Г��A��9��\Va�G��?[��쮬!�Uq(v�z$2�"�	&�KZ�(y�&�Nr+v�Z�R:�8��(�����T]�5���h�|�+���y��_0D=fNSd{�06}�{%2�h��<>K���U�L��<����>���я}ʡ?qQb�g��魴Gw�T������ J��-F�v�*!�������O�gU��&���M��GT?죿�;��q���߭�PF�J�+s1�ɘ �h�<|M������x���me��nd���(4���ŋ�2�!�ƙ~ܴ8�v��A�������노�P�{ ��ڭ�Ʊ����N>����Ԏ�ÅAT������@����A(���S�����<D<�f��Wny7�Y��%�G��G���S���ZVZaG�%�oD���6X�lĪ���R��cf�q�;p�P��� ��[��"؃{qxR��wQ���M��C��w7�Y�>e�Iu��"�ܣ���Z�T�!�?����^�Vs֢�Nٙ16��|���<&U���T̀5` ��sTg'����a��Y�| 33 X�n���  ��z�TL�� ������!�Xv��(^HM_�O�
���J�gF�V�Tw�ze��	��� i�zs�߮��_�q�X<��N��
'�ōT��ܩ<O�;��d��
�
�G�*�/�\��/!t�W�' ��F!�T�*_`{��{蘢�+�J�(��1~�z��y>�t�O�; +%�9u��J�3Ĝ @Y=��-���~4h����۠���J�8�z@/�&��z�G��WNk�@�OT�����+�!�z�;�zS��U�?�$��
MN�ێ�ǀj)��gYa�Q��P������>����[|�*M�j�0�ޠ��[���0k�ϸW����6�Z@��]�<R'�X$a%H&D�߰��@8���ӗ��uA�70�ޟuA�y�^0���9B]��Z�w8����_��_C�gRi�CC���=�]��� �%�Cw�����iŅ�$�`�Wy�_�8�� ��.����E2ĴСu��:�ߡ�!�-����L��n!D���J����Z��S�A�����Y��G�T��E�AF 	E�2�tH
A0�S�T�=^L+����b ��lv�E��札�?��Q�$�+�fj��)�r:_ճnU>�!�D80�f�{��v��X��g��X� �h;�*܆�B� �@��b��k-�BQ�i�b��D����C�D��vE�b��e�+0��ư 3%iM������"C��P�u`� ���eJ4�\�.T04�˜EU���r��.���2���s�9�s��=8�����B۳��V�b=e{�tm%��m��.��Z�e`�Ƈ����&�/�b{i��Fu�j�dMZ:zg��s���1�L ���5ޤnU�N��<�z0 k��;����NY];��@g�l�P�]���$�� ���Kz��Ҡ �Z�l	,�m8:qo��{D�ɶ��k����B�ϧ�S5x���ծi����U�W;�餸·����Q�����̛�py^�y��o��/]���/_�( �؋�!2���B�]$R42��EeYB��y�*������^��}���b$�~��, }���xy� �+����G�%a"�s�^�ݳ�=�N�<�+�ʎ�k�I�C`_�E�(.����G�+R��y�v��u��B֖�MD��OX�z��5g��������&v���8\�0C*��r/5] �!���6-�Գa�cLO,Bh�q���w�Z����=��� �/�Ѱ?/��_ΒB��3����1��rbLpN�3��	ge���˘`[�2��?-��d���F��x�tXW�<�Z)������� ���p�<
��$������b���b-64Nd�p��A8ƃu3kU7�Jg�)L�k���N�ah�jNȆ��\ȦZ�c����+c�0��	�� �^�����<���_Fx2XK^����'ol�� ���*8����d�t)Y�_� һ�`P=���`�u���pb��K<`���W��+�Ɵ뭴B�����D8�Ў�an� }M���e<�ޔ��1Q��W��-��ੲ��"��V�2
*R� �=��	���8���e�9w�!�qe��U���ǞH��P�cbxb|(��-����H/����S���S/��o>���C_������>�ZHL��6�VT�r�[����~G��U6!Ɨ�[��D��jm�`�aH��Q�!�X�</�_�m[��[����i�� VO��m�, �Sv���wd����j��m8vw���/;�|��s��p���X���Ñc�X��ي)�n�b�u�e�}^8��[c�(!���R�O���ϸ�Zv�A���Rz,��w��L�7��y�ov"�ʐ5�� �0�=@���~pB��PΪWY0�I���3�Y0�/�uX�96�C��q�슲m��W��h�����0��E��"/��ٮ��������[#�6��m��Y
E�"�j�E8�T�(�3�xy̮MR'���}.��Dx�q1;���yFc[�	Pv�!���c l�K�ܰ��b�]���w������}��	��}f����a/��P�X�����7�RM-;6�X8)D�����z��쒾���ܬj1e�n�f8�e������+>����󳗻��>��: �V�h�0�+Д7j�� &���&Ѻ�HK��?�"�0����{� ��� ,��9�ˡ�T֨ut*���me�u�!�ҭ���[���M �b۹:{<[�R���������Y�Ϛ��;�����U*����~�JSx�Jh�=c%��ܯ�aSz^�g{�e�5������Hz��ϥ�O~:}�7|M�����a���H{հ��3�%��]�.��R!͖�9,&p}��:��fgws"�Ҟ�Ǒ��H�`m8J޾�B��sX��ʱ@A70�b����Dvj�Z����a�-��wC$��\�rm����1�	�8FZq ��^t	����T?
����?���~B�wv�~���8ip�[�H���8q(htU$�2��}�Z�n��v#(��"Ev��v��P����C ��DQ�������0A�; �$=s��$�uW @�6,�؂�3EϢ��rc����^��1��L��rj�r/&>��w��ϬL���AH����$C�0����c�do� ��Z5Մ��Ɍ
JUx�c�6�� ���@P��F�}��0�ò�uS���!b  DYU�dν���`#B�l�g� %g��T��|UP�خWc�]hQ���d���ۊX�E�b�6���w8Xq��ae���E,����2��L!Ć�'Bd�x�0hy���Q<S{fs�У��`�w 
~2�J�Y`@ ��I�7X&lN8��"��r�ޡ8��f��ɫ����3�A�k2Us�S�����}���� ]�@��F���흡��`5�2��a���\���w9����L����o���BXqe���>�5+�k�I816����>�9��:Y{�y�"���|.�-�N�S�ĥt����g��;�D�f��?���o������f␒��*G/ϜK��b���F�[�'�֮\H�c{t�z��.�a��"k��(�bW���W%z�yh�vTF*_�b-P@��ŏ<�dh J�	*'��v�*Ȉ����ݰ׫v����Z Y8��)_c	�q\,v��+����q|���� T��w�����[hГi3(oiX�F�����p}�(�F�`��:)8�\Z�EH�+�O�Km�N�#3X(�ƚ[.�7�X2L �K�$9/@����r�1�i���p9��a�pX��ݱh�� ��w���"��n ���g���}1_BZ%
*������b_Z�-��:��C�N���T@�V�?�F�v6�Af��5�}p�v�w9ę���T�-�����z����P������s��c��k�=�dܶ�4���O�;�!y��kO�ϟ�kf^��:6a�<g�O֥�����G����,����JDϥ~O�c���}سhIr���PT1�c]��d���|��+��L���W���b�}����^��m���@�ȿ�� �s�H" D��</�^�r9P��cG��)�R�'��&�k�Јjw��r����<���ȁ��?�G�?���N3ϥ��qO�'�׿M�<���J��a��?�W�w}�itl ��?�'����ӿ��O�ob'�y�0 쫠S���bp�h	�fr�Z#:{<vz��T������`{�(�D�t�~��ơ琉����k��ݹ�ﳳΟ�#m[���*��j��gX��
��� ��r�.�c�]���w����e;ӌt�l�VxD����P�:BN���v3�!>^��d���Ǜ�V�� �;��8qt2���؟�+ʎfTUfI��E����p�.������l����B}|6���x;�g&%t!�_ΔȎ#�K�4ؖ\K��f%8��#��]����jg�vME��]xv��:wY�G��+g���h�dp��(�;��2 �Ƥ�g�\�C���w��/�J�l�>��=gJ�����אs{j?���y��8��j��5@�F���z�����"���=,WU@�kʡ8�*Ӕ���ڀT�������̸0N��lg��}�5__�e{g`���������E;j�����Ξ�s��l���pc�?2��!�&������_�m|:�o��� e@���N
$I�S�V&m� g�ZS�U�`e�R���iY�g�sګ�?��%�ӟ�����1Z�<t�	�W�Fu�T���w�'��o<�Z�
wB�-��-��Ԑ�󘯊�Lj7�v��IL`�T^o't��J{vA<M�2��Ȉ��o2{�z:���Ũ}Qs���][��]�S9*��8F6���'��Ŕ��"w�vh!X��c�A�+07$�Uj{%.�h������o��̠�㤚v���q,.��G����ݮ#*\��z���i!��P��δ�W�q�bprd��{r�C���uBUZyδ���`�||��Z�ɋ5�t��l�v��N���%������w����PSe;Gb��[W����k	&��fdG�=��U�ZT�_;��E,�|F0*`G�q�]�3���<U�I�f���������Y>O�_��8�R�#! DnF�_�u4g28�X�@(_K���}�2@����S��X��A���b�2C����Ӟ�9ڵ�ϣ��lH-^yN_Ϩ������Ή9a�G���r+�/�|�0��$V���σY����v��k�6kg��!���:!d�M%.P��[k˅��s�=�z�^_�������g{C�������:�����ӿ�qi���&������'T}],r�v������Ks��JX=�������C��2�$��5����C5h�:)��Z�X*��<n�ύ俜�\��ֶ@A72~A�����9[&��*QB8a��^h�䅟�U%��`�'c&S�m`(�C;�l�Cw�M��~[do4�k�9��z��%RdQ��d&�_�bݍ�F��c#lT�Z10?�?�^~���o��2�,/n�}�rF�C3�"���]�v�R9;Z�M�?���I�Z��G�\��3���(h1(B٠��vod�j�Ɓ���z�B�%��0L�E��#L��:��x��y��k9~�w�\��Z&���Aq���ö{p�w2kD�̙j�Ai�σо=\z�p��<�# �����^�Η�v������D/�-�>\{�厪0bv��[(_��<��9���<��͈9H��k)��X��t���ܱ����g(�_���/^��l��L�#D������u�^ZZh.�Bׄ��Y�L?>ü�=��B�و��q���<����t2E����'5����T���ֈ��u\}����\��x3��{��
���q��3�m ���y��I�;����F6�j�#Y�Z�\1Zz.jt����>Uվ�������m��Tk�.��첢=-%V4	�S�[H������2�������FLY�U�jC6��Bz�����+�o@��c��m5\��I|�u�[��~t��ŤK����k�p��GJB� (ov���W�
����Â
�o�U�Z�^��B�Pe�x�Ks���f��n*�S�+;$��m�bU$�XY�I�]�r��S�ISo�MB	I�0� �Z J�8e�ә��
0�:��}����N�N�v�`n�L-�Ut<"�q= �@tnc�����Z�Wɤ�D��T �k�K�CF|Ζ>5ObQgA��C�s0]�fL��*������<q�0-v8h��69��w���|�<��� ��?�Ϻ��w�9�9W��1��2���l��=J�'�M��EA� f�c�(�r�^�P�'Ӎ+�˅�48���C��*�s�,�\1��%���Y���=�Q���{?�a��!� �U�r����~�#��Ρ�0�ưC��{f&�~)��s�a����i��$����ɽ����0!p^��z��g���x��hZT�΃�79y��ƢP�։f�yn���������-gp�pf�8e�9�Ky����P�'�J,\o7�ٶ�p��z6���*�]�-7I�Xi)�>��j��GL<���QC\���^HT8q�ѩ�óʜ��3�uakD�qT}�Ⱥ՚5��GBt�Ue�=�S�(����t�5�e뮫���O��ށ�jk���w8�O�(=���ɖS�j&��Y�[%$���+���n`�]�ǆ�k�����(�H�|�6�v��� '�ȖKl�5�E'�>߂c�,����V������E�`/��m;�H9��7�ќi��E�ؙ��,k�1�	zE�Z���@h���Z�����,�)�NV��q�
}��#b^Rh�3�H	A�.�3�T
�vyv�0/f�9pO�~P�BdS�ɺ��j�}�
��8�e ̡4X��D���9;��1�L�흮�ag�C��}�踕���5�Y�p8��r�j.U�7U���^P�Y��"2Aa�.�@s�Kۡb��r�9���a�k�s���qf�<�"�ʫ}��Gȶ���|��jKgǜ�'��u�T���sw���9��������'�S\��!�LŜsH���Ffo�D�&나��ޓ0D��������2�k�z�.��'<����&F�!�x|���U�W�Wf�4��a1��W����g��EMK��rTѮ�:�Cy|�����ꁹ'�Γ���S�и��y�WZ�.�p�4D���IG��sZhc9����t�-��w���H���w&z�҈��h[@gG5�:`�7�錊*>��K�"�]N�lߧ�iSi�0b�Cc�1h�S�=S�il�xz������ϦgN�u�X�޳���T5��̺��(���.�{k[���7a��QTl����Z֑uBժ�~j����WC�k�}9���p�_z��Uq��S��^G�{�� bfF��A�!����bC|H;��z@�j�T�e�"x��H�%����Uub�wC��)�hc�ʵ ����)��������q/tg!5��������n��Z��* H؂]7bk������>�� Qt���\s�F�q����O����-[��i9sث,"��q�륪a�Չl1��}~�C���4v.�K�&�F�0'��Y�g��cG�8�qW��A��r&`u|�o.֗{da�-�6�"/�@�C��p�赢�|�+��'�z����}�2�j���Ɏ�g�7 �����p�k���R�Y�� 6!�e*�ﶁc��
��T�����v=� GNq���s��0&��k 6�箻����64�７1�S\=��)�8߻Ǩ2fhŘ/h�\�gו��"�.������g�eXf)��.�s�{Ό_imx������	��4��>3Fn��zAhv�ldd�R����{��w��Kcb~'�G�g>�4��8��ݷ�P��B��?���@��;n��J�h�߫jLs����ڊ�"��-b����)qف�o=��<pO�V���z��ОT�<��*F�n��Q�^I��Q��L���җ;���ߺ( �Ʈ*W�nC���\U�#�A��pp��_�I�]���>�ŧ�3�_z������9�+رR?d@�b�z'Nx,RU:&��Ml��X�@�]g��=��Mqo8�\���a(m�o��֕��w�(`Ȃ�N�0:W��"o�&G�K΢��PW(�E�ir�ܢ!gj�� ��\�k�εJy�ޓC/�/U�%۸��iw�v�m8�ރ�u�����3��]!�������{J��3��H[ �H��z|e0�GȩЕ�Y��,Jf0��FA��dQy��sD��1��= $1��C|��P���7�q�dV�}����Ο2
��$�2�k	�G"�n����:v~&rh�lY�2�[b�۪ @�_>��� �
=y|�^�N�2�`;x��O���z-���1���ܔ׹6�s���2��#h�V�l�2l�5�����٬ |���Ҟe�{ܪ��̲I{)�6k62��*�)*�,H�M��N��4�d�	eq�x�c#B��U���J��������������[��c�	ZO����l����c�~���4�sZ�۫�Ѭ}+�J�P��m����|z����<�zǦҠjK�=��(�ZE*�RFj�;���@�'��r�7:�����( �F�O���B�YO�cY@�v'V�W��|j��������}�K'r�{a9pZ�:i�.�� �P�MgW�R,��e��*�2�X0�㇓��[A��{v�xQ�)�B�+�Ąi���=����1S�uX�Va�c5w�X�V�u=���g̰T:��H�����0��]����sv�����dX<�:���F��s1��5r��U����_�{�ﱑa��6���3 �nt�4j�1!R�:,���u��s��Y'�Ӳ3����mƞ{��'9��E�@In3(əKo��ɶk�d�o2X��Dv�y12ۘá\C�c���� +�7�<�.g����A�k-��p��e������&&��Ŗe]U~�x��_<_�����E¼)�]/b\�}3v�;�v��J���%�N���y�SE�����}��h����)���WM�c�!���Ǽ���y: Kd�*³k�K�Ra�(w�7~�7�G�|z��j�XYW�c�;x츲��B�W��W���z	JX}uz.]�zE��H����耲�.��J��M������SuX5�:h����u�ֺ�O#{���7�ڕ����5�u��|m��"ݽ�8�v��7:����R( �F�+�UZ7"��A��c�nn���r !^�lMv濙bQ�V��d���vГ�z�nU��k�Ϡ�pJ(�Cג��P��Q�:@HN��*���k��YK���ѫbuz�e������ ZZU�C�C���Ř�1@:O���l�
��b�?��_�)��4��(�2m0m�����g�9��V%
#U��2�$P
��@�1��l�G�uL^��W�OֺXoD(���haQ1��i;3��З��~\��v-�ru�.1f�S��,ZdD(��{[,֎��l��Q���؄��qrϙ!�N,��tݙ�����t0�E�K�������dp�>gہ��\{fX��8Ute9�
�GO� ���=5�9R1{yNy>W��^��*t8١�����C�]f��v͂��3�����e�����+vK.�Y]���sߖ��+���D'�1DCG������wD��vf�k6���=�f*��5�#z~�Ħ�V��M)7�}������V2Ӫt`���0o�UC��)���3�H���=��`�V���Yg�޿_��GF�����)ė���H���P���� i�N?��G��.���f.+D��^c{�hyM�ohCﶦ�w��M}���3�����z^���K+�*�^O/]M��t�����J/]�����*2��Z��9!;2;k�}9�[���� �aN�5���o�X�5��� ���,��_,�uA
>X�W�|�ICT��w���0܂�n�z�1gMƓ9�}u;yb�ľ"L[N=R��.�܎@Y,��.ޘEW^P;����N��.40hk���ڷ$h��`�6��4�ۢ��@߀T�uD���Jݷ�:fcv[nha�q�d�H�����Pz'*튮��#z����7Ů�zk3hԩ���0�*���Ԕ+W/,/�!���+]�#���]�Ȣ�` �	
p��]{$�CE��*�X�~��B��{tMjsВ&�~R��DcXgV��z��"�2��l�a�3�3�<]3��z�U���U�� Ե`�B�0A=�n����XON)�#����[ti���!1.ن���Fֱ�@����=NլW>6,��� K��m�����X�e��я�{U#&o:ܚª�pfܲ3Bbͭ`W*��ff�����!\�V�0=λ����j:�k�ޖ�\�Z'�K�]���*��#�HQ���W�&l2�l&�,�Ě<3���	P8BH�gW6Y�Ƃ�����a��h}⢄�jγQ	p�}^��YD٢�����CG<�n��k!�ݛ�{�Ζ�86���ٳiAa*lb��6��N�s�Z�� ���OC��;�Ÿ���~!}�?(1�������[Jm_]ZI'�I��#��4���"-@�o�^�G�.S)�kLU�WӲR�;d�~��U�&�t�N��.i�&�>m+����t�i�؉4<�H=�;;�Щ%�m���j��64M_�������߿( ��F��j�"�ˡ����*ڛ�k�D�|i
����.9Ț/yw�����ô!~�.f�PJ�-�C�Y^"f �FD@�B���om���ڵ#���{Mяǎ6j�X�]�`bWkڞ���-C#ғ�G��r�ⅴ�^Qd���S;�ɀ(�y1%_�o�T��*�d�Z�oto�>�y׍#��[�NO_M�OO�Kt��f@,���
5�A��W��i7U9\�!�ٱ�rQ�и����-̾H�	p��.���dG����U�0��"k9�ʑr<7��f�SV�O��S�Ք�&FN�ά���Q��?YKE=ܜ=Vμ7?~\;�%i9f� az{w,v��7�������-s0��x�Y����"kX+^�|��)��}�Cfb�#�fM������;�
��53K��c��RT��[i��l���0�1cn�&��܎ۣ��}��F�sW ؙ��]0���A6+A��˕7��g�:\�bZ�d{J���o��oN��}�e* ��S�BsY�o����#���du;�������PGJ�%}sm�w����!B���g>�~��~L�X�;��-�++���]bnв� ��U]��ŋ�
�t�]w�!�η��ѣJ�2�h�+0pb̯^�I�
���t�7Ž���I �/�=[N��,�7{媎����oJLx�*fh+�6WӰ�*����Ӓ�ua^=��6Ԭ�G��Rw��N%�KȤ^���j��_�( �6H�G�	�uo�3��W��p$�<�ηS�E���T�8�����رq�0"��8j�IU�Tv����~��ZY�0�k4y�1�D�����p�Nd@�ܢ#}d�D��Z:�w��}�{M�gMC79��>���*�߶��u�Z7�f"B[����2 bAǙ�����Kit��n��Q�`Ɉ!,{�`��c��m�h��-����XiQ�r�]���p�r0R�11]��zk��?�i���Ύˎ�� Ӗ�qe9V�l+����`��М����9��q����}�;#�l��r�^�Wr�^9J�J���6�`�^�ۀ�'6�T`C�0&�	.���������w}�w�f.Qp3�$���x��y�����[;k?,Snw���7O��7�?���@����-k�r�0�١!�6�fi&�o`H����|�ؘ�ߎ�̡!9���]�zw�_��#�ߛ�������Ӯ+�&��0<W��|N�@a�{��y�	��ʛ��}��;p�������7]����d�Ǌ���/\�ܿ�[��Z�%^�银"@G6�#�<bM�7~�7��h���F��6Ŷ��ы�@E�]�1�7���@����<��X_z������ϷZu�s�lR�gGzƁt�������l35S���k�4���}�0S&Zss���#�z-���
����Ro,lD���� ������]`!p2���%��xs�+ǥE��ͺ(m�U^��3�P�:����'ӷc��p���Jt�'�� �����Q�P�����*������_U;��x�0A�D��13@q���bސCw:���[�
{ 3+� 9N��`�^N��|_z���ipX;X����	�  D���3�K�Twg�!��,�`uwm���[������p����O��?V��;����Ä�e��9),�x3*�ŎW;`6��a����lH�2��-�}��O���O|"=��fw4��w!ʪ��+S@�-�P���z5���$�sc�X�C7,&l���[^I�|�C��sߟ��m�e�t�^�K�.�^���Ei���xv�j�|�v�L�g*>*��� �(4CX	���ރӥ�p���59�V��|��Z����`�ٜ���PS�I��n���tp~�#j��mzF��[��*�6(M�$W� d�E��^���t |]\T���(�������.\Z�3����y �����?K��P�z����=�q���}�������[f��U�bC�u���[�w�T:~􀚪Ω% L:����sS�;b�-���v�jg�3@���
�i�6]��i��1b�R�C����s�!����O�m���"	z��"L�X��?)���Fmg���e�&( ���sx,ZZxs�=m�<���X�_ ���_Z���𲣮��)�8s.�~o�A�'4 $x�i1����t�}�Iԧ�⊳�ܺ0����u�2*}�'\�g�ӒRsYH��k�&}��|�ŨgN��uf�s��ώawW�P��a��w��E�ŕ��
[9�xo��ᵤ]h��[T}��j��#_��`P�KQ�:��[�ȶ𢻦ٮ��@C{K
��`����w����ZD�otIPuݙ��3ϺFM�N��0 ˵e�c���,h��xe�;��4r
�y���4�GB6�����O�9��^�v(���뤩˞.Pɼ�ޭ�i>l���}�]�/�~&��9�g
�����Р+L3';|�?���	q'+mJ�-� �}���+S���#�vɀ"_weF��Ie4gR����	��^I�o��t����ҬCG�����R9�����ML���8o���f�w�����;q�Ҵ�9c��c_L���Z��=����^ �J���m��	�X�j'Qu�LP�Q���V:
�nT�G ���s��F� A�U6��r������~��ނi�c<K04 �?�?��t�w�Y��B^u�J��K���+.����w>��i�Q������1�����Κ[[k�q!�F����W�]��ӽ�ݫPۢBi���Z¨�ز:�SChyI�[5^�R��rZi����v���ꍸ����i�ʹ��`G������6�@A70��o��;^���ڳ���k�������@�|c�^��^��W��y�� afK���%6[a��dĳ�8(T�D#�LiC�9���#��8d' "L��P�3�d}rT�m8kI.i���l��_x����w�ig�vf�lvh��?v���v��b{��bQw�����By�f��[o�9����w���?��:s�t��N=�}=�B���4��Q23���W�A.��5y�����,�n}���Jw�f�SO=���������-�����x�w�a7�Q�{"ٌ�Bt|m9D�ٛMi �4+�O'�˯�z����OX��cv���-G�� �f���B�U"V�-ɺ9A�+��)\�:�^�������ΨH�%�|~����������wλ�T�F���v�0f�=Ö��"ff�~ה�h�Wd]99A�0ٺ"�b�������x���?o��o����!�=}���������ܸ&���A�������Y���Z���a�?�����J����t��)����+�����HO�8��`�t� �&�@�wg<JϷ�Y/�\�~��Y�K�B!����N�^�2x�Գ�6�����Q����|������~o���|�����=�d��u�h�Lv�6<���(�}4�TK�Ad��]��Z�أM���\�j@!+͛˗.Z�`FC����-��r\ӈ ك>�гt��	����t{��J��Wl���}�/}ʎ�@�0�G������� Ͳ��?�cwUu�ӓs��f�����` Ex�
�$�$A	��������a209�ι�+����}v�3=��L��?�z�����>��{ιg����{7��L޲�o�6z�����p�?���ge����A����w�r�P�Ŗ]��r�{sq5��X�@po� ��c�GcPŤ��®ҡ� e�Z�>�b�2`������V���92@ۖ�\c���gE��ػ��U��H.�}j1���pQPv�ZV�n�x��y������c��򒗾�|�/?PN:�$-��eb�ds�w� �����iP���Ge��
������Զ�2�~q˽���QI���>o)�׭.�~��ʕ߻���������m`0��7>���?���n)��0�O�� �ņ��н��/�+amy�{��0����1~ի^��o�fRk�L���njdD�8����$�7�f_�%C��Epޣ�>�;�O|��C�Pٹ{Yѷ�<��*O�姗/}�?�"Qe�"jǟQ�Z�+�i�Z�iD���dL9b   �)�	l#��)a�Qrý�o����7��|�ӟ.�wn� �����Cҙ(�7ŵ<���܌$Өsdcj�`	�yWb�v2�;���c��s�5ה���_�˯�ܺ��=����xy9�Q甯~��:z���M���;٧|~���9_y����F��������]��� ���\nP����9��{��_'v�!EG�	L7`��)�x���"WW ����ϻ�ȕ�AkƆ�,R���}�|�ӟ�u��Fz�ﾠ<��Ow�����7�7e�r�0��D���Sc���zѧl�\�c����G<L����>�պ<~�[�^�֐pѹ�46���ͼ�����K����� �� }`|o���r�-7�1=�]j����A1��{U�LݲO����eU��H���vn)�z:Z��̝�7�y��̎�_�;�7�{�䁡Ѯ�ˇ%؞�Q�f�=oko�
��sV?3�9G�-]:%	�)X斞1�0���w���90H)L/k��ŶM�)E�Y�ҠiV��g�:N�d�8��uP�]_V	��	}�ލ��ض���.����ꁀk����	�%s^�{��u�гkqqH��N��Hj��EhQ�"����"�� -�]��yR���{`��q:Hn��kWy�w�o�;^�6n����@�>�z�a�)����_�0u@�1Io{��yQ��<X�_��xg�n�7�,߁�O��l���^w�,�\�벀��q���AC��7)eㆍ�������(�Ʋa���w���q�Y忾�������Y�%�'��,0g��yِ�����aCW't��܉��-�|�3��@ h��QY]^����a�;��������]u�gZ3sZ��l`�6퓼��5���6�ȵw���iW�x���'?Y>�5 Z�r���}�s�)g�,W�x����]�I�s�2����R�8#\�b�9���k�d�E5~fA�
�x?�)O)'�|�������s����r������=w�`՗�a#R��1�Q� ����O�>i��G�t�l�pls����B��G?Z����ҫ�9��򲗽��Y��ܦ�y��u��J��2A���P S&l���.��VKP�X�:>�3=�.��2��8���EP���-��|}���?���=��e��NLC�O�A��M�^}f�(�`�������:���7K/����/��^�yĜ����ny�����#�K.SD뀑��<9�)���a0u��H,{�'�sĦ-t���Z�tTEs�ca�����j^S,��DX%�L�����i��l����,��T��2�	X�j�-+�^zi�v���7/����S��KK˃�z�X�����o,]-�=m������ۚ������ͱ��M�M*tR"r��5���ԾwF�ш��P��wN F�;��թZcg�'iV��h�פ���r�c6����bKZ)4;�ci�d*��tV�lLl�>�ߴ����;{P}�P���5�����/}�.��9m�O=�ԫ�>�+�CM�O�� �0F|^c��P��{���;�{[$�������TM{��6<F_#�K�Az�F�(!��wP�n6��,�?�9q}.=��d}�Q�%�d�|��֮�B�{���Pn��E�*���b�0�0�$��A���ǜ��^_��W� |�_2��7������/g�u��$cs��+|<�m���*�n���
��ݥ@VÈ��}�{o�R%���N?�m8]�������=H�y�\ ��B�Y�@Ȼw� b�Ƅ�h��~���XM�U�N�K��q���x/��r�]���w�׼��e���2�������=�l:rS��5�h�骰��1}���_C����#�������� ����rĚM�w����W�W�9��[�̦��B���d���_A(�EEe���qM\n��	�(��E��42Z�bæ��S$�P�z��c�)���3�]��������UX�𕯲�Ρ����sA�O2��u��'P������%[c'훘+�͜���`�MoWoy����x�+���!O���;�0� etW^�=�9��w��R䍉�B����R��Ѳ}�v��?��﷼�-n��뿖e�׫4Ĕ��p	�O�*�n�p�gA�y�Щ�c�o4\qfv�ϸ����>H��s�����?��.�eT��]��qDs�R%���r���[��5��h�y% �V���4����l����vq$t$�����:�`��� �y��Kӽ��%���=9W�"͇k������H9B�չ�>�\s�5嚫�����	
��9X�%�����꯾�%e�e�ms��g'$�l���kmk�`M�RL�S�}�\��w��v��ܬƱ�t ���Ҝ�̜�g3��3���xN�����]�6s:fN� �&m���� ~��zf6�75����Nj=��'=��#6m�������}����_���0��O�WA�����4�zḿ������{�EŬp�n�mz���U�'��~�py�cD�G!�3J�7I�0��X8-R�y��6Q6��߹u[��p�)'I��;|��K��c��I�T ̤�\nZ�"��6U�W~ �R�u�7:��Moz�싾s�������򗿼l�$���3wև��7�\�<9ћ�w�t/,��;L�������_e@.��2kN8����w���r�)�[n1xs^��%8d�%�^�}#�<������#�wja�'랓j�;��)*m� F��IO~�ټ?}�[zv���ۿ+W_}MY�c��$C��z��  z/rN�d�</ݤЁ`����X�p��6Q^�◖���۠n��b`y����o�9���.J
�6�~�H�9	�i/��ߓl�e�&��dKg�FRu  !*�2�j0D�/zы��A�>=��o~.�k�xq>�~>�^.�&��ZTXs Dx6�,=n(��M7��{�� u��@�s�����?ݶZ�x�]�����Q_�:"��$ &z$\���G���Qn��A.B���.�`�φ�we��|�Ϲ01�_jX��g{k�2�9�b������?�s��t3[��J�2(`@j~�8�21;�l�]J�1w���r����+���kָ3��v�~�DKp3N��]e�`�p�"�_��֖Ve��͑
�Dݢ����u��?��;-&�r�U�/�vl-S�=*��?���x�1eǖ������\d��Hͷ��+��ڿoN�[D�4�uv��u�x_��5I{47�bE3A�<��rF��Ts*�ɵk����Ӥ��\��m�C}l��S�6# #��J7��A���o��U���9�E!��a}4�N=����O>�G�����M��}[�]uǌ�ϯEt���b��$R�i���@X�{|)��=�?tq�/&�����y��ު���3㢡��"��t�@����9+��E�J���&"�N��f��M�s�N�u4����B��%���+F�W�1;��2��A��-R�<8(��}v�K����b`q��U�Vڨ:^�җ�=����n���VLǰ��a�%uR��
��I��2(S�!l&[�������Z�I�v�j����K��h7.B،FÖ�+�q��V�)�b�������q)��(�1�hX��*_ Ӥ�\y��~����������f�?.P������UF�j(3p����M�V8���r�/�vW ~"j�E��v�1�KUy�촓N���V~�)?�]+n8�"���v��A��L���E�6��(q��\��]��=�E��Ι�X� �8յ�y����c0 ��8|p��)T�&���|�����=��]�Q�t��oZ��
�ݤ�C�D� �I��a���]�l��K�� �
���ҿ}�u� �,�Ò��}Fs�%�����W��k�q^��g>�:\��I~�(l).j�W!�i@��"e$N����=�صx�:�X��|�7��ՏU~ƅg�1Kw�-��O�y>��~����3�>\+F��c�ZX��o��\|��z�������[>���T����v���� �Ѯ'] �_����_�)%q"����g��eҰ��,k�u�c�*M��u��zB�����ȁ��n.����̌�<�]��jͪ=�㝽KF���)Bv���D����.���葇wfF �S@��j.��y����O��aN�O����j�Ӧ�jQ?�h l���6������S��K��i�jW�~�7B���u-�7u�c{����ƢYk���'�x�>�G�C>_A����Ԣb'��HZ���V�k�w��K;쵨�'l�yy�3�d�}�B_Y,��1��,..@FwZ6e!�H�ء�|� ���916�ZX���.�k���Yvn�M#����2
{��uJ�=H��=��`�5F�6�rqӈ_��|���[�������W;] z�$�|�+^)V���;���ZL34=��Gu�%=J�z�;^���Y��$��P2�#T=�"�9]E{���4>��L��駞Vv��N�pT�۬E���Q��ɇD?�ֱ��q�ӎ(��;Z�,�d���C��:��(Na�P�N )��s����/~�\w�JMp��ĥm�;�6� ���5+�8�>B�N�U�)�Q�"/�� y��Uv/<��s˳�9��7+�x�4'\����-ޠ��2D���u�"MIv��ġԎ
�t���pM�t���U9dd�	E9�.�j"�RL��0�-�H2��n�Zz�'sSOh�`	8/._�`�hDJ2/ �f�@̙�#�U>W�'�Ͽ͞�?\�������D�x�1��nW����=
�)U�9�Gf̘/5h 3fG�e \���ah�������@߀;���/������1�^_�� �+�J�ad��H��G�gua����U
@���ث�ӹ}t�۴� W��MG��Qcܛ&j�m�_yy�=�q���//;u7����/~�<���v����F$�)�x��6�M_̨� �{Cr[�M*��k_��ǋ��㞻�a[���w�܄�Q���t��^m�Vo(�.�:x�ƳM9�V�9;E9��^��ѳN:�?����(|�U?���" ����M݊xY�U�����?Z4O��m�{V{}$j\��q�G�9�$�����uz_O�^b�[�<�]�ڪ睷c�B��	��t����3N?}��������v���zFv���s&�� �0�}fl�yv�%U�>G�y!0v�'�C2<
cB�{�X�Bg�lR��o��g���qP"1��5! D(�X�v��e}�on�
	���U�hQY"��Gn�v�
�2d����d�D?��*C{����yO��3	�z�����S�l]���b�^E	�
�/���N퐹=���TbqB�D�!S�j+�vьLkGv���)c�F`��J�j	i�c�B���U��->�]e^�CTvC���
mN R�����R���qF�x5F�y���	'�\�ؼ���k"��KYF({��([�f٣�b�����Nډ
Q���ݸ�?�o�S?Kd;.W���$�,�BH)0�62:]� �}h��N\��1�2!��\;� �qjfL�$ˮR���Q_H��p�EA��aZLaP���M��'�~X7��Ssc��fRV�=�ɣ��!�9� ���9�&�H�<e@?�L�o:e������H��µ���� w��g&L}�.��ф-"c8O��;�z,���h��sB�"�:�(1f�`1e�f��Ä[sR��V !Q6�9v�Sa�sN��P����=�r�F�۸360"f��'�`:��J���� �=K��$������4�:":;4�y�?�9�[ fV����/�^��%�sP��nX�	���+��,�˗��;f���@��Hխ�b�zB��2���˩��#�]�����Ĥ�}l�tܚ�G���{��}s��f���G>�a�B��G�{���|ƕ�׷�I0���$�mry��R�h�	x�J��lE�~Vλ 1@ο"�?�&��n��N����bug=r��X[��i�*]☞�Y1���G��L��ڴ�����O>�������=��7��b��������)?^-YA�1^^2XP�����Q�ÀN��W�1L��s��/��4�\�ݻA=�*��퇗`J[��(p�\Om66M��o,���&Y�� !�J��z��`D�$�!�2�C^����.�X����)�9���_��UO��ya� ��;��^v�S C-� @�!@�����F[ �@��	T�TT�����DG��3U -�a#�r�ɲ���� T��-�U9zB��1�b� ��w �����e7
cD?��r]-X�H*�:�_Z��ႁ^p�jk���伄�ʘ�=hH��ف�� ��9�)�׮8�(J+A�����
v����+�������zFet8*�WfmWh�  D�*��E�� �)��U��#�{D(2��
�{ڗ����uyk0b�Y�䅋C��G;�1Ր��k� ��<�Y/�$�!�7��Wj�RK�|������Wf��]�ʢ�p/�V�x�`�`���5�HVI?��D*��j��!��z1�R�!��}	ۅp F4}����   IDAT��ȵ�fdTc�ry��^�Fw75��;�^|��fLp]Პ���؈�pw	�;j�6=[`3@��*��ȥuwII0{�x� �������oܚ�����C�neEV�!s2Q�R��{��r�uוg��3�G�9c]���[F�}���z��o�V�'��6�<��1�	�A_f c��g���z�-��OQ��Xtm*�ڶL�H��jF�R��n��!�<5*���1a���i�Etx#�U��^��=T�G]懂 ���R[��yJ������E�l��ܦj�]~�wV�)���#6�n-ڰB M)9�0�x*fԙ��EӋ��<��lU4ǔ.�#�٥Wy7n� � ?���v���Z���(E�C��%,~x3Aj'T>fT�����1�H��X�7���N�|LA�����Ź2C�d� �%͈@�%b���n��ϫ>�4��
X��31��}UgЇ;���9S�l`-�/t1$�P�bIg�Mqo� '/ra��]a\&e�ڕ�������(s�.��.�5��V��)��T���R�R�i4[�5�Co�9nڴ��OZ�� ]�I`ڄqI��1��:��=�r�`g�y7*��W5����$�Б��"q��N@���L����H6��*�M�V���H<����R�c�oW�����3��W��6e"C� �k 3�U~��7��|j��<Q(4�5;v&x��^��C&f�I\p��H�5�H�hw����(N+�c ٤��+M���:�MJ��1��pa�6�9?�q����%֣9��(5��`���q� (�sb�`�j�i�	��}=����c�z%�~X�� t@-�l��w��]J�U�n��W�������t��+N@�7�c0��'c\����>mtT�L�$���TG��A����kS�T=�btG���J�g����e��yj�Ij���OM,���j-bɵ�xY�
�K��E�*@��,�;w3���šY�F�A�;QS��y~AeaܿOy~n+�u�(�E��P�w�X�(P�!dmv��2;�V�,U�V���O>E.�=1E���hTK
Cc�g �A���Ls�?�7���QUH!$!�Љs��
c���*C�>��]O(|��a� ��!w��\*A��E�AuX��̈́l+���#�#��� h��4t&n[�l/ ��$zYl�(t<�Fz������b��B�;�\�Ղ�̑7	%V����>�63ЙUԞ .
>�0��;-s�p-'�������꓈`���j�"��7s�[�#�����p��]�� 5��	7i?�����\�Quj+F��r�F��5�| /�4��0KT�Q������)�Me0��Y.����l���{����@��!��Z[p;�!#^�e�
j�>cd�Q ��WtM�7�3_�$��"b�dY�|f�L9��g��.�M8�s3�d�Ft� HZG�;ˀ8����O!h��2ĳ��sTm�L]�w��q)~��D��h����?�Dg¨�Zֿ������� �c��.f�6>KNe,Cbg�����Tʊ6��ڷ3j���S�	��d�O!�׵a�xx8��vɅ78>��\*�*h�
$�+^�_�u�-R�6&�Z��:���e\l�"tv������q�����kA��f�\��esa?�74.��vM,SdC��creQ��u�Xt`г���c��8+�* 
�NMg["��O��R�^��[�k�+�߫Eh���Ұ��=h�u�9稀��f�>��ăJ�ȇ��A~�[:'׶�cgk�1-h�0��@�C$D\��B�6j]�����6���X ���@]�C@�I�&��aq��Q�X8�}b����:�� ���rn��	�<�\) *
�E�)�^�kdHh;fG���j�7Y��?�`?3�*�dd��R`P7b ��\]]h��>��U�dUG�2uR<��G�*v�$���4�e `#��耘r�2�H�QD�ъ�Bn>�3�A�̆���`4��0�#� ����s�|_�W @����>G5�97z1oH�0����{�KLFS-����V&��x�f�)���B�X��G�D<�9�ZN�5���=��,�|F�6�XW,ܶw������y�{N��?�Y�{P��������w ��abn;5�cF�����dA�J��/D��f���{����u�y��p]���B�+��&r��e��AT�;����R��]�g�7�j�w:ˠt�����:�+q���zmJ_"
�+w�A�?T����D�Vvw�9�GA�)#���K����+�vPE�>|%gT��4qm��p�)��@��Y���1���>��䨀��T!¬a�5�t��C�էr����&�Ώ�Ո>��\�~����%�5��X��֯3� �T��������o{AA����'ѲY9Q���^(fT�͊�K%]eր�c�*�B��pW~1�e����W
���CJDYͫ�r,�a�c���M�UBs#���Y��f��h	��]Vƙ"�0S,�Q:� ��6�8\�"�òTwE�؏�&7�Nh 2���F��;�9��DD�XlЂ5�}(�/�~`b��Uf��>c��3|u��ZO,�5���n��*��
`��]:O�Y�	��F�[&C�.2��0H����E5��w�h"b'Jm��2iWe� ��qz9��3ˊ��cB�	��,�;�GbS׃�Ǻ�`�t~�R0K�S��߰-�:�T�h���b^h� ��Ɣ�w����s�έ��;�,Y�����TjT��L��k�z1@����{�,�k��u�P���4T�/A�YT���Wd��te?�3yz�h9j�6� F�8���|�M��S��A �% �ov��� I��c����Iͅ~�����0��d�&!��ilzڴ9SZU�P��߿ҥY~��^~�!g�~����ʐ���t������3XfO<�w�QX XZ+'�p�O�jo&ꆫ]s�����<�S%�n-��8P�$����UR�A�16V^+�v�6�U$E-Tg�⯟�Xd�k��(�4�^D2�p����#ռ&�����s����RP9�p��h2�щlB����p��Y��Q�'D����17& �b�M����hvh��ѰvSc��Y��.����0#����d��n�ܒÆ���;�&+D�c�Xܜ,��A�~���H_�F��04�F��"�J���X��ŁB4	�#r	��H!]�*@Ӏ>B��Z7��ɴXڸUMNFq��#D@�T�
#�9Bۓ!��Vm�����̔tOji mD�0�� Ȇڠ��6�\+�0����`E¥6_c*��0q��<��"�3�^1��O�������Tc0�G��864-�� �/ے�@#�A�����s��xL9�3����>�le�~Fy�C����U?i������T̃|��$t?��C���@�ܟ�j�`��B�7 �v��X���>��H�s��{v� ��EϺc����-:3��x�8�ɂ�
��8s-���v�����Z� �lW^��R���&fs�Ϗ�Ž��e�ÏY<~��&�<�w��9�!�ϱ������:�(��1��h��hk���+�?#GV@�k�G�o"��3?�ĉk��g��qY'�ED�w�����Qf�E����ٷ�������;���u�l��)�o�6_o|���:q���8yS��tp�6 ��LoZ�|�e�����L�a��x=�aXb������8w~���Q�>3���nl�1%�z>�By0��ڧ���V%�ӂG">rgP_jRB�Equi7�����o��"0�]��(�� Ǯ�X6(�F�v\�Z�o��z�v{gժ����B��?FA�\_�x+��	�ɢ�D͠q��i��+� �=.*�S�W�V��G"�(��ϵ1 DFQ*��M�@;<B��u>tA��tYv�Zxq1�y?.���ʈ�CV[:I #J�ȱ����R�&������ �Q��������Y���dd�]�lPB|�g�Sʝ_ù)�}3�>�������B�թ���i�7Qpɮ.�M0.�����W��>�AAה��]�����zֳ~����,b\��w��u���!ȍ��z��8��O��&��n�lG��1C7S7<��TG��P`w�\qI�-0I��}�߸�E8`ڭӍ�g����� �pfu.�gw\F<��������آ�0���>������3�{0u@�����y���n��'� �����%��Ч�b�f����V�*.aAz94��/��Y�k��~�Ck�9�O�������2�3W����H-3_�a�Q�eY���UB�%��-�il��6��P��1m@
֗���kZ��r��c{H!m�Q��� s[�lw�@g�"�(����\�a�"Y�@�M;��9]D�G���6"5FԮc�0W��4��^b���|���{`��k`Nq����@���b�F(F.�C_���[s�t��V"�&_�Bx�|�$��M��ain��cnZ��2	͠ȅ�G���ŤO��֞�t�r�vlDfj��L���)�� �����=u�[P�t�M.�� �*��;��f�%��,S�� 
��_��`���C��CaF-zYu>Y��1��`\P�D��ygN�&Ј����Ε���{\gXf�}14�:�$?���'hS�IjuyY3#k��P-R�a>�)�A�[<Z��v*�Q�� �\��ţ��0�f}%&�ς��"�P���ݔx��i#��(n�d�<O�6܀�­���|r�Ufʺ��J�=/>�9��tuw���v)�����#�OI1o���S`d�4B{��ا�s�
��
Q
�΃ԃ
�-yoЏ1ga��p.ړ�&YϜ����VkV���=�7P{0R2�
6�l���n* �Ne!87mc|<_*���������]&���\6 0}�{0Fzܰ�A�����}Ŀ*�K�i������K<O�����[���Rq����sM�z~��YtA�o4a�Hh��F�繃:G�;< �ni�@�P$U�zFѤ������y�7��DGح�oʬ0����QE�H�P��ܪ5���*��D�_�jj"�Q��ŵVe5V(G���Q��K\>*P�u�H:ʆ�/��/����7�+[��i��%߽����o�{Ri֯�:�M�XO��i��W�C����*�a�ܤ�aQ}v�����1- A�e�� -��� �v~7��hr�]j��3z�[Z���%!����Eƿ�#L2)� �uƴS�P��
hav��ܖk1�x�á��	�C+��P�
�w�$�h+��VX�a+X�X �QHS��I��|x�f �Sp D�2�J�n ���)��^�2�.����<�!F��;zYӣv��.ڋ� ��v�2�b}l�|�X��F�9ޠe�����6���S���8C��vH/T�C�R���'��5�@�u2:!���]dc�v��v#�R����W��V@�q�0�w=2�����K�M5p�u,�Uw	}�c<N:�de�]Qv��D����]|��v?Ў�ڑu�	�� c0y�P3�O�bi�Z����4� ��(���/�G��e��p�Et!�������-���i�) �{>T&	pD3}ܾvӆ��� ���{jk��h,�1�m�S���(8�+��s��]������'�#}���XF�`P�%�\�VnB�c\��0��i��&ɜ���(L�$S(�n����9ah}F)�C9�K�tTnz��s�A\�����q�K���,]��c��1\��F�"��S��q�>p����׿Z�UY��N;�l���T��%�sܹ���i��^�U���O���L�a�q�5��� E9��ٛr�vd��§�"3k,����-������x7It�Q*�w��%&C;+�o&�9a0��D5ô`Hud��9�X�z%T�i/w���we��~ة�q����)@C��Ek�Q�0 �s$���8"Q5��Е�!A!��@N��j�$����ذ�"^�%�r�Ο���~5�DSm�"���5��zA��1pVae�G'��)�$?�#�H��@*�^�:� ���Hq��pof�zlӳ�Ny�r�]��iGc���d�0Zb�� ��
�ŘQ��A�<'l�j�=���l�LP9'����f9S��	��5D�q"b�\;M�י�f����nL�<"�&�t�:A���fX�2�Y�9�h�6B�q�!$W��.H���V�l�����0ٖԝ��rm.�O�ie��N@)Z�Y�ҍ�&���!A��鈢�3�A�L-�j�+H�K ��� s�9�9�kOc��G��(?�ju'1ޞ�l"
�MTٚ�g��-D��Cn
��� �|��7� ��,��q����.���l^���*�F��1�ٲl�
�A�td���SD��t0��g�Dmt�I��XJ1�&���k#�W�r�맽m�#M��`&���k��}��R^��=_p�M�h}p��&r�0�~���%�������YH��]�J����ig�����+����v�ª�h^ZK��pZ�V�H���a؊ů���E&�0�F��)[f�O�燩i�y�#�8~��3��E�B-����4�;X��y�aт]�8Y��!�E�L�^%�;���S�-��z=y����%�G�U%|J(�(�)e�V��q��9-�,�$-���c�,7�~��ګ쪚�a��Mq���ʡ3*�t��˪�8����C����ۨ[c�����;..m�\���~�G$� ��(2@��( j`��(į�J�\2M�H�@6�ӂG��nh4?`Q��2��ԧt #�UvY�!M�DٷG�?���M(d<ht��"�,�unZ蝹�z�wg�� �@�v�wы �e7�O���@?�B;y�t�l�1�'��L�5\�������%�:ҏQ�+`-�#�*s�DԺ�i�S�ש����<4c���n[�'��v�C6t��k\3�i�	�+D��oGQ�ڙ�M=*�:)f���9�+�U� cءy1�Q�n��Ʋ�e�-�b]��"�0���,�Mt8bdGj&��Y��"�
(Q���p�.�9���'�v
�G���sűT6Oc�k ��ѩ�J[�9�v��<L@�����^�Q���%U*kn)��`��fʣ*Κ��'z�ρ3��(g���]?N����O���eY�̺����$e|u�V��c���p2ʇ�Ϙ���B�iPX��SJUt)��ʜ�ɉ,%$G�?���hS[ft!^̥p�(#���J��C��5Qɞ�1�?�3{����h���m�:u`�6�"����J��m��l��2��5��'@:�cg4���!��Y [[7ͭ����|�\u�b�����_�6cZ;�` (km��_��Y����"tCV��E@���?�U0UmKLK��;6N��#_�C�r�U?P�5���~�g	mfW�,�+���G�0���"����
p�����Z '�e�t��n�#�Ԃr��7�uJ*�y�rb˦ҹTQC��3��j���阘����K:X��]��!ؙ��c
�5Ô���Z$���J���~"�0Y�#�lZ����!J�~��+�r���iX߹��ۜ�xRmb�O
5�+���:"a0�>oU��
��a�yj-MK/��|���$Qi�y8F��mD-���o��5�G4�!�˱*.�<�.�ta��m"W���2ڴ���:�0����M��sN"�y�R��GT�D��n���@�N���� V`킄�r�^���p�`�Cfw������b`���΃��o��C��}2�d�$ÈA�~����w�v���2�����$%�c�G:_��sϹA �	p�n�f樒.��� 0Y\���e����؍�)"qxչf�,�� T��b
R��V��0����"�>�aD]�T��}f� �75�-܄o������=�F`z(ܘ��� 70��bԩs�c��)� E����1"!b���#�$��fb�?'��6�a�**l�u~�tJ�]֯f�Y�X�)G�+�B��Y	��~��)(�"�̳�<��q����5�;�s�u�63\K��`�d��%�p�;E�zLl�n@{�Y?�_��j^Sό�%A��V#p`�D��s&n͉�Q����R?K�D����W6)O�*�ؤ��ގ �M��B�wsm���(h~%���c�	:�1�3#;y����W��`��Q�O���7z�ͺ ��]
A%[-�r���~�������}2R}�\Љs�9����ZDHH�S��]8:%Hm/va��٨v�-Zغ�1jo��Of'�5���c�pQ�R��	W
����h6�� �R!D4$�cwR��ZA��'�oF}
r]2��q�m�U�Ͳ蜔1��i�\d�-΄u��w�[��1�\����PV�n�͆���2l�!���C��mAj��e���F�s��`��ϺG�H�?`� u^q5���9��K�>Ǖ�¡�J̙�Kb��7��Z^vu9^Cc�t
_��YֿRI�-~��r���hǽB�O1FU�ù87�����Uv#���Q�*���^���hG�D�	�F����ŋc�$���7�ol��/�����4�8'ғq�ֲ�o��׫,�$�L�0hjeUw>�oS��: ��L�yO�$Μ?���炙+��6��q��w�¬ߕ�t�'��o��a���8�tK�� Y���f�D�	�����2�ų�3�s1�VZ�铑�9��r��Mб�]����7��-�ɑ�~�j����y�`N@��qk	lV��2�Z7XwAX��[��U�ݴ��a%�lW(�D�P�sb���P�VT�'��7a�gt�ܖ���ƤGnᙩQ�h�V��Ea�K?I�/2A�9��_����B{����c4�@?\��b�w��6��8��&����v�h2��[�c0<c#���|����q�������.D�*1�*��ev(�<�m2�=�ϙ*kǏDQ����NeO��!�Ɯ� ��ؑ�1�Ckbwn��(�Y:���	$�c�ć��!��.��n)D�S���`���Ϙ�b���kW{!&Q����H���е �Z�b`�I����ar���6�3vd��+i��7̂� $�7bC���V���^h�Bf#�P�0İY�*�>���@PlND�D��S<�� �=Mh������P�fڕ ���Q?��q=-�3FCͱ�/m4�P8� 6�2�YS��ͰX�O|�S2t�˙g��q�`]�F�Nن>���_���__��A�KD^��y�J`\���Y$.`ˏ50���lT�K�1O(����)F�c�`~������ �1�.�u�p�dɌ��m�=�����`3�#�ŋc�K	x������fD���/!��l�*��|��
�׮B=���	�b�G!Z�3�!��������f���g��V��
��=d~,�h�c��	�0����M�RIV�ڼY�;����;����kw,2'{%wW;ωj}�/W��и���ݽ{�ֺA1A�c	 զhQ���>fX���k��}7��Gsp\�3&'��5�m�f(`�����LA*!_��fz���ô�?N__A�1Zf��Ө��;��!��Y����.���d���`E0������� ||
q/>{��T�&tW �?�y��=Щ�1�z�c��\+K���zbRt��9LRE!����{q�`gE$E
���aXj9f^K%�D�aw@	V�
NG��&��Ν;j�
n�������85�k\<�d��AY*&��0`���P\���4BZ�%6(�@�f��U��f����axj���z�[�b\޳b�M�{�mF���B�@�����d����f�N��$YG8�C2���O�+������t.�U�Q���w7m:� j����O��Qd�>��m��r�^hI���Hc���b@с�������v�3��_?��5;ˉ'��H��va�����_P.���EJ��d�0� (���(ے��1��6�$�\x(sܦf`����F0����� ~�H���W���g]��B>�f;��2��(E�W�l�D�)�yN6���^�J���Pdr���X��8�0���SG��:^v[R)����xڗ��X��AU|��x��x���/�LF0�d��O�!^v���s3��֘O5����� ��iLp�nX��������v߶us$U���L�p�w�֛#�?AA�r�o���mykY&`�k�N�X>;wl0"g�)�	F����C!�Z/n���#�;�t��*�PE���M�UǬך��K;��ZF�g�^Z�ha�-����� �0F��@̻��U���pe��ra�nd�~D�LQ��ع�aU8�w�,��4f%6���tT�a��$N9�$�49d�����1-ڰA��Ds�o(�t�	acH�?�4�-�u�^M�E���������H{���E��5F7��Q���lD*����k���(^ ����Ȫ���8��r�"=n���؝�;�fi��C�Kc �DY�m:`W�V�?��0$�hX�A|�E`���l�F1� X�FM��-��LP����3:#��t�ѩn��=�
���a�aÅ[�蜚Lcc������ ��A�v$� ���[т�v����c���0IR��40�N���H;}w�2�M �����@����2 @s�1G� ���6�%������ng� �x�%�:�&��Am�~1������S�=.�v�İ�蚍N�h��g(�*�G�j��6�5����'��s5A(׶��n�p�;����`'��c��t���PS���<uT�"�)�Xe�d���A��s�l��Ǽ�儕�5�8��)� *���R�d��zew�څ�'A9}i$���c'X{�C�ļa$r^�Z�������T�cWy�~�ERٶL�5B�Ӷ��,��~q��ݿ�ŠI2J1f�W딈� ڷ�?����b��G�ZE1�Kz`\;˩*�A$�)�?�P�m��i��P�}p/Y#���5�G.i-Ǯ��9�w��������1�R2Z�p�I-��2�����I��6v��H�\�x�d����3���f�hڑ:�X˔4+��yZk=h���mo�)�16�JTeG�-�Z|=�XA���=1*]����c�z/��K�g irw�;��|jw;�C��T��z$VHB(��+�biƴ�_����vl���A��أůM�m]F�A�G���"�:�g��:�����xr�6(X�K
v��� *��`!"�pDu��TE�1^,���p��0�G�t-\$��A���f��CFXt���p������]e��E6��G�#����/Ԧ"��s�P�^�:$'~� ���b`�:)��7	���"�j"�`b)��u�L��1�zd�%��#<�e#Su?K����n0|��.�6}�����~w�fԚ�k$�^m��F&�>1��lOʴ��O����=.�V��ރU=�#�M��NY�!�0"��D�B��;!󸬔jA�s���P;T+����|���g?cƈ]��@nT�(���f��<��d����H��A��F�FȆ��S�Ǧc�4ޅ���'�H���0�0S0-��z�=����?�S��_��Ѱ]Q��=���>�	>b�N��%v�Sj���\2/`�h��`#�F��Zs��0w]?�nu��V�9�?��V�<Rޘ��lD"�/N�~$� �2����j���J�ϊ�JPB��W}v��7x.;i�j�Q��<@S���scT�a�'�Q{f��8֪	=�۴6�yםe�j">���]�Їx�B�i��ε���厛n�i�\\Z.W���e1���%�	�����*�k>v����t��������w������+���O6�v�i�seF�	���l�(�/�mr�wv�	,�"�mY�'T�ar��XAr���4>��&̓f~���Y>���Gσ�x�]c�c�g���{��}��o�����֭�d^����� �~u��Ul?	����#b�Ch}Z�%�����
��)�a���������
W/ǠePv�Q�c��=ZHY��g�zQT�o���`��!!�a�٘�*\S�pSC��#ZN�-��i�/f@~y"� V�(Wr3Sn�sk�Ff���~��s�30 ���9կ[��«bf2��{�1�1!�U��Y�M��m��b���A[%��~�p�e�9�pBٲ9�P��!D�AQe�]��KE�R8?��2��"3!p3.� �B�Y�S�M���4Q�ÌX�1 aͬ��B����r!V]?��Q��R��z�Ȯ�B��Ex����,.y�ZPyU���]96�D��0$��o� `�r�`��A#����NY�% ���� ���q��N���`�y�8 5]3~����`e!�yIC���V�]��KU����>Q޲Q$�E�����E��C�Ir��W�Y�]M sZڝe8\�������k��I-�󽸿��u�M��Zus�A�6Kj�(Λz�dar�Hp���\K���������;�eo�<j~iMp��3��6����q�Yֹ������i��u��Rx�`a�5��gրSN9�<��/�w��U\�c=��m[��%dr�W?j��������v�˹��;�,�.mH!��zV>RRPv���=�ts9r��r��e׶���պ{�{�FĊ��,K�Ԭ���=hfp����c�h����ޣ'��7�L�U��Y=�3��Csʍ�����*Ay3�Lx���G�,D�KӐ{5�cѤy֤1֣��$���ޜ����={����Ϫ_��w )~�f�,I�65~��'m�z>�l�_8��f&����>��"��]u��\/z�S,�7ҷߎ�	��B�O#͟W�$o�z���C�ª�	B93�;�,%�Wj+%ج��>�� ��-��"*p�,�"3SA����uN�6Rj{*+�ع��_�����2���Xpt�R-�i���f��1��f�,��z�����[,�D�X�����YaW��1I���Bx����$��}��� �FQ�@�o�����^�牭@ŉu����|�
�=����BM�v��lw�r!�}��P�`" ��11�6�Du�1BN��� T����'�e��$�~YЭ��^s�ϕ�GqU��2�`!Gƿ�E�P��M���.�9�׀ň���;Ŀّ�&'�����R�D���ۣb�0�g���/���̂�-R$��c��]��H1q>\;ˢ����e?A	2+�r������FC (uX�^����0@�1���C���&56��ʟD���\k�v�k�7B1�	�l����&�~��Sl�\�lB�>}�k�Pju!�Ʃ����P����5`�{���}�K�Sܢl|�'�և$������։�p�`���7�0�r��R��ti�_��ؠy���� j����G�
0��}���O)+=v@i��ե���NI����σ "���=��rm*_�2cM_H��d����K�W���Q�|����="�}w�"#�X`����y�⒋ڛ�g&2�r��֞��&1�M]��M�+�^��ѓ�4{��=8�wL ͏3��pe�9��p�)������G�L��#[��FS5��_/�����f桞�qM�s���J����qۭ�/���(���g��u�f���/����a��/�C��t3���|�&��\��F��ޚc���F��{�`�Y�u�A�6еt�YQ�����:�墎@TWg!.\52f$�`���.}����(a��u�)\��+n\/,�s�Y	�'��s*H#) P���.��[jw0���B?אav�XO��'g�K�8��4B/���}�'���X`�ѽ �F�3�E�.�<D�D�9�cT�m�FF��-bp!C�^(\�c�Y?��Tʂ�:.h�n֒�~�J=����J
��!�r����.���X3WN��3��1�;�bX1Xb��Y6�G��5����D�״��%1n* n.j�9�Jk���LW5��/��a|q��( Ee}��c�x�`7"�Hԧ��*��ME����p���ۈ�ͱC7������y�Դ�{��(ߒ�X5�O�p#s�n�6y��K�K�r�{�m�λȜ5����j;��b��n#���4�bt�����I-Tc!�!';�s�g�kTc�yl����U�]�I������ Hce��ƀ��������r��m�hǈX��{:'�"Ƙ��X#��n $�6z�	��� ���?��'	�<�"v�g��-w�&��z
��C[����+&Y� ֨\����9�bgר�R�!ˀ�9��(�P�d�t�4u�@U���_�H���%�*��'��Si���9�3���:��έ���ۮ�٥�V�k��Sv�I���MN���ܵ�u��AaE]��)L� ���.lV}������B����:�c:^�j����푘�q=�Sz�E�D^�0�@�yi���;F����~}w1��=-�|g��.�o� �maG�'=}d��}�5�Q���6�7��ޮ�e6���L��
U�d��UB�̭Z�z��wꁇ�=��	n1�Z��5Ǳ�ڙ�j1bW�}Xa���԰U��={mb��r�E~xv���홁"���퓗�<gb72���� ��z*���"�3N\';�q�lk9�\1��`��$������N>k+�ǎH��������a�N�a'�Ӡe��Ha4���o�v�<��Q�� q�
����oټ��`B�/.���93\O�E�#���)�5�S��`��C�		L���i��2X܇� i	*���Ǚ�TB����@;>cl�MCBԣh�+C�D~�Pr�(�6�1!��=C�����K�6��+C�>8�5�T��f3� ��lP���lq4nf����_�T���p�nC��
���6�Oj��d�0ܩ�q��\�w��$��ݩ��ڎ����01 ��`�]�{x.�������nV�}Οs#�,E�K� �1�q�<E0�� 7�	2��W/����-2�G���B�|_��7'j/�6H�� ��{N�����au3 H����sJ�Jn(x� H����n\w�u�r9N5�X3wn��4}(�n���\)�Ї��J�z����2>]e�r�9�h�z�X-���;��N�/����v�TT\�+�������=�����ԧ����
�Ö���3E����+����7I�<973���;��ؽkjnJ��-sJ͡�unJ����a\hf���gi���&����I����Lͨ/g J9_�r�j����������֏�j�����o�����9a�ZE�k�$�W���6���X|ݯXA����~06[p>�L/$$C�������].@(��=�P�} y@��s�ߴ3�eJ-��ј@�`"@!��,�$�Nh�&wZ���+�ɕ�_c����q��[sd٥R#2J���r��
dAC{���l烵Ц�2���0�m�ŝ]L�o6Վ�F>B����#�}�_�����dOfv�9%E�А
�R40�	Q~ ؎�Y	��b������ט�H9�Ō�W��Ϊ�W�-P�����-��e�M�?I�a� ��0Ҥ�m���x��٭51"Q6%
Fm�ۅ{1��Q�o�k�K_S�=��,��� I�/,�+�{�[_�83'�YƽKF��3�x���#r�!�U�^�~��JȺݮ�*�~�x�T���D���1�0��)!:�������Y@�P��p#��9�Lח�ߐ�j�H��Y����g�* ����w�սH f\��_�9�>s�~E�߭�c%v��;D��{�Q�CT�^������ʫ��G� �'�`���� ���d���@HX���7솎c~����T`�L4��cC����1��殻'�c�����q���zp��6か
�>����q�2��]��M��ǅ���.Q%�J�m
9g�F�C���w�Q��r��ǔ����9��E����g�"
/����ȇ?̌���|���\����5�����u޲m�J���1�u�Mײ���s��A�o�jW\7Qg}+�	ýLAc�U��nrwu�M<἟Y��'������,<4��$��":��S>����fB1:а9� �)�
4��Ր���~Q]]#���q�b�a�Ij����:�~,H����
�1� ���u1��B�;jn}L��2-�r�Ѧ&��E��vO_iV��Z�Ě��TVˈ�|�lA��sfL_Yx]hSL��3�mj�A��Ȁ�9�+�	�O�vU����u���I-XD�E]'j*!vh��D]+��V�}ø�q���(�5,����]�!#�Ga�,�d�&�G�#A���V������t�,��RV�l������ʡ�Ӹ�^ppզz��p[-ފ�!���&Ѓ�i��A-��qR�^�@LYgF��`ȴ�ӏ\5���|� *��%6Z�kN�^�H�[Q��lR��4�}��ic��(T�%*QQN��Ui�=�ZT\��0�  �*���;lZ8�I��
t8t(�]�� �»���C�NX׬Y��
�Rd$%DՏ@�����A�&�W�~&f�E-�UUH�&%����xRbě��41�S$z��ʳ1*���KpB��!'�=�n�~|��������Ăp�ԝ�I)`�S���6�H��:a�HE�KʸØ)���A��u݇Kd�H�; p�x�Rp���\�t\�,���g�t-�U�m��~��z���l�K�賌R$�r��o�И!�Í�����E�1m::�ĭ�`C=;�	�]�vX)7��ğu���+�+�W~��5ɥ@5�t�i�]�$���zr�S��q����&���oH��Q�Q�'�Y+0:��6���|Q��6+}��q�'��=JܸO)%��?�׊��|߫2+������Xq����>sfa�?f=��c�`�����0vQ怄�5ח_w�D"�Ljb�������kMGDJ�Gi�)����M\�n�a�N��:�DD��'�/v�Ӕ�Htu�_���9�\0EW,��n�^�@����Yg��Zv�~k^B���O9�!�VL	�����������3,�2 z��MU�.1�� `<�����ȒL��
�߸�|@�̌��9�c ���E8j������]�ڟ��G>�����C�=h?F��	�� 1_V��>�Q�Z�ЖK{aם�qGya����Z��@�{H����t�߰CZ��2�P�#���Wax��& �5A$�Xq�Ї��1"�����g4Rf���
E�	Ɩݻ�zڭY�GQ(Ww�"���N�dR�#3sɂE(��EF4�I|02�P_����_]`��o�Y��RG8�b���`��U_9c��F�!�$���EuUq���{��%���E��WIW?X�ԉٍˆ�^;�,��byX�5��(:*�7�6D'���(��� �\�Mmh�6q���l\[|ϕ\p��&
���7�G�/���2�\��]��s���I�s��y��#�<�d��*��sr̅��۔;�_�zy�c'O]2%�F	���=��~M9Qn3���A�(��:\����l��������ԍs���wͳ^�Kl�Z׺tyYջ��a]����~�Fk��Vj�[������ڴ�(�G؝���A�a��>o.������:_��`-���O���K�Ԩݸ����{6�6(bL�v(�ho�arp� �D״Kǔ_�{��`d+F��/F%� ��xY �s`$Fw�28:b�F�\2�-b�L���.WH*�3��	�ЧqC�Q82�W�E��^~|'��oY���� �ES��i���}A�햱�z�V*�M��.-�,��p
�-[��]L��1��R���H`��؀\��j�wؘ %��������~ZY�Vn �-b��  /e��D��ukו�����F��U
9'pH��h�uN��܊�:���Y�	�	�3��X�aX�$A�C�RM�5�W+��6��$EH�q�ܮ����'@^�fK���lW�p���� v�G����-P�AtD�\���t	q�4M�lٲ�Y�!��=Dy�`�l�a��7fNqU����(�q��,��������"�4 $bޜ�hY�)�1	�8��B�s��:i���2z>ȭcM.��}�縌��hb���G)�|�]�'�t�57��O����7�G{�8W�����z)VOV�k��Eغu@zq�s�y�Hj^g�!�v�]E���'=ɹ�`u�%�&�'?����}�s3B�^��NP�O#��vn�J�0��y�c�Z��CNi���	�X�Ʋ\�7�>�hi�FU��*/�p����5��s�v�_��aΝ�Z�@th��>�&6isb�F�r6��CG�蔫�˕(�p����C{*�Y������������":���0��� �&�ҹC�Q�0a4�`�{a��`PhVh$���h���g#;������jË� ����b�NI�(�H�^,"Z�v���z��N9�e(�,�L
,��+{��R�
_��\��ػgo���z��"���oVE��N���)2;���4v���i�^�pQ]�u̴��v%��8l	��Z��KeX�1N�j߰n�����fu����`Y��;`����wA땺�F��]:G�y@L�.19�(Wʄ���=���˥�^"�q�r�l��a���%C�>%��6k/8 n����]��'�- 7�d�#�7eIb�)� |���"@��"^E�Q��?�A���?g]F���^1Ǔ}��T��cN�D��<ĺv[yΔ�n��|�_,����A�~�ܮ�����+��a������fƷ�A���̂�+�3^�:EZ \Dοd�� Ap�@��O|�Jhy����^6K���c��?��r��T��ps3��ݬ8�[�·���ߩuJ��<�/�^F�e�E�
ox����k�i����v��/��G�N�� I&��s&�I�'�w�K���s��O��f�*�F;H~�3˜��۽|��_��_����s~ٺm����g�ē�v�aa�z��`� (h�8n��-c�$�6�.�d��{+Uje�uڨ(7�zs٣5g��b,��y-�94�[�}�=I�Dz�a) OWeOO�<H�����vP+n;�oFa�d\_�D	�3�6���G��Y����=����M%�I!,��tdT��C���x%�t(����cTS�T�ֺ�蛵p�x� B�(M~xP����~Ƞ
���W�\CcZ�����@a D%r�m!+@P�&�KK�dN�׾����x��y��>�h�O~��(�'pСE�Ą�s\��;W��6�$�]Q\F�@���>�	��E?�x�"�F�W@�ý�����]P6m�Tr�C�7ܨv�6��я~�|�ӟu���64(�@��e�=���Q0SQ#A�B�x&��q%��J��+����YgA�$���הo�;����.�[�6+Ae��D��Bb�l,��a�vb�I�X��:ܰ�Ox�C�p���y��(/��x�.pّ����q��j��s��\y�{�+Q�v�t�%��\(cya�+jӹ"��K��(��Yើb.� q>�э���i��_��r�"������|�;˷��-�܇�)ǞR�:묪�R&��t!��Q��p�|��B=1sF�N�ӣ�>��$#�n���}��o�+����=���ɟ�s�{t��W�^>��U���o��\n��k��`^Υ�a>�� �d�8ֆ��¨�������o*�{��̚|�0� ��Y�����5O���@��	�
�D�_\Չ��P�y��׈�c��|�����|��Y.���b}>�����_(^|I�� !�s�4>�@�mĦDz)�>K5��EF�P����ފħk��c��i�ֺp��7I4���Yܵ���E	��*�=�vz>�~F�'�>�OaZ#�W�A)�G ����r=��dL������&�{��w}rC��̪/�ǡ�~�z���OF,���G-d�dy�YXT�25��(�A������Ac?�Y�0��z`��<W��֪��L� ���x�a��%cW��(����;��ۋ��c��M��}�-�Eь��f����ɚf�3�(\ﱳ���>�Ϟ�+�RViW7������{G�¬�N�?t3vi�v��L��Mh��*���q�л`lm���Q��;E��� ���/��\tمe�c�O�'=�g�㽫����)�������J"<9Jg�� h��s���>����?�:�s���} ���W�,檩���b����~����o.��r�2�����>�<�ϔ� �����W�0�E��Sb�N���8�7�Xd�V���y��p�J�N$�E]T���>*���c��6������� P����>��t�D��p�Ŝ
=�ua�IP���h`�4�� N�[�9��L����*���»��.�3�:���MZ.���2:3R��x�����=��h&�mDv!��#`�yp�3�׬��_���9R�q3Sl�c���-oy�ٯo����o,�|�9���//_��r±�;�h�X
'� �]�Y��dGV�ŸD2�2_`��|>V�X�/���z	�/��²{��r�
�����q��%%�
�;�|���%��N�Y���$"8+@��H�2�M�ܴ=���sIʉ�E������|�_q:4i�T��y��}��5��	6#]����o`����:n��W�Ĉ���S�y��̒��:a�fs�D�%~�siwf�(��2��U�N8�2�,�o�Ԧ�U� ��@�d1���Zs�Y�>ǂ���)�Et��E}F���S\.D+�?-���$�3X2���Wh)j��y��|��j`4'Iag���G$Z_)��|�B�ךw��|�h�FW�ő:�^ #�� 0�����X���v!�۵��%$=u>��0Z�����1T�޶m�w��׭+�>�Q��o}���W#ˮ�Ӟ���{/�]-����P�~ja������5Qf����sF-jb!��q챻5���\�4��З���r嵗����m�*�-�)$�?�6�+V��� �4Bڳ�C�V#�n�
T�'��t��>��{��q��»\yQ���/;���3�(_��ʍ��X��������/��8U���W*��܏����-Q�Q��@�evC?�n�4������������Շ���T��'>�	�ÊR�lذa^��C�n���`���p��7ㅻmF9��ah~��'�\F�b�)�p��������90t�Vm*/|������Z�K*��� �3�����A��5L�X�t�)¨2�¯v���tDy�K^b��[�EW|�lZst������聲G./X=
�f�-Ν0�"�_ͣ�  ���o�Cߥ��.�Z��t��@�s��g�ּ9�s������%D����p�&�.GRD��s �֯��Nm��3���'������ek��#��-�� 
n�g�E��O�W&���t����]2㙿�Lύ�r�1q#�U�h��-��pR��w)�{@c�};���)��<�X�?e=m���|=�w^P���O+���i\�����y�Ѧ)8�[�<=l$t�ZFHr� w��+��?N=��s���(1V�>�y�"2��Bñ ��
���F��7"ن\�,�$���h8j���H4~�0�hm��ūߏ>�L)�\}��XY�fU9�Me�Ļ���j�Y?�0s�=�Q����+_i0�[��L��򗿬<뙿&�i\�k3jwIƛ�<`,-���87�KU�k�:dkn&����ҭ�Q�-n�׾���6�ַ��r�uז��#W���!��{v��zY��%�J���+V�Qw��zP���u�+��h�P�
�K�V��w�m9�r���_*/}�KZ~�U׸H)������@,3̈́0<j�����D�!M`�;}��n���a��o������ovx9���J�.���lF�x$ӕzG	��Ꚑ�(�T��yE���fH�� ��s�u@J�G��g�g��g?�.J)�v�Z�9	q:�=?�*�k��e������a�O��3��m��~���屏;_���o��mxO;����W��\�2���n�A0@�`���"{�y#���?la�Sxm�����YC�t�a����'�׽�u������g YƈW���:Q�=Ϡ#�"��8�"�^��툣�>�y�s�� `���������|�|����&[��N���Qr,����!�223b���*#�m����f�����кW'c���x¬c#}���B��2e�?��1��~��Տ�����-��vq��"��](��FVYm�4S�70B-�h����,S&i6�c1X6.Zx�������XA�7X�0;)M
ތ�v�z@CC�����1�����)wL�4��ra�A���P���C��gA�-`aA�!�<�O���'��c�._����������� �T#ڭ�u��]U���ᢘ��Jų�+�����׾�<�)O)��r�v���EB�5`�ڤ���Vi�F�f�$p�!�J�D������O�)�B�۶�Gi7��?z��Q_}�U���?J;�9plV��i�ltL�L�4���թ���e' 2#��L?�+ƵO;ߓN<Q��A����<�)�U�z�uS��}B{Ө���ŬScU]f��b8�_�=�[�7ƕW����;��y�'&���7�����L���N)�5\�>�e���Q����f���
� �t4#�~㪠>bQ#��`��@�r�<��/O����k��N�㖲jժ`��W��2�!�1��Kw%�]�js��H����I�.F�?�ؾ�i���)�́���e���H����<|�1�k�U��������g��J�� �{�_������8��V���W�O��dܸЮ�$5Kk��_�j�]��F���
Q�\���$mUd܀�9�5֮�E��k��*t<v�Ƌ�y���eG� ���Wq��|�@Q�"�D�j��$�ޠT�5����r�r6FN��} �b-��Ԉk���v���K�{Q٪����m$�Zy�z�t���Kz��c��]�'����j���XA���bLv�ս��,-RH�Z "��������@��?�i7��S�4o�ݔ
0`sXib��ѥEN�,�{�;˙g�!�+�\��;�nw.
�N)�N���FgU��]��c���n�ŋP�G?���m��#�X|qP�#�8�l�r�Ԛ�Hݡ�~"�������
����V��b5%��
N�>L��E�P�nz���v�a��u���E1 �}ܞ��%�a<#<�b�V@Ye��wF��C�uP�����c�H�~�`a=�łq�|-aX�X\cA�i��`�^X�4���䈢���>�*���o|î�
��B�:�0��`gޝꢛ��<4ڜ���� ��U�v��ۑ���`<��J(H߂ȗ~�I�1����ZD�NnT��k�(s3�3�,�w}�P�y��n��R�Esf���	�a>r�5�\:r��r�^f!2lz����|����9*��>+ǜ���߇������8�h�F�q��\�Թ�ݵ��b�����}���Y����D�)W���с���h�����W�!� (j&R�-`j�6�ʚԓ��H?��<�7)��ǟ����6ou�V���+��Y��kV�&�U,�˒�J��{D��{�z��?�.ߓ�Ɍ���08��j? K���� %���N~�Q�]����_���1ю>��ث���k7�#֮.�ܹ����nk�.N�hmU$�zp<Z[D7.��=J^� ��ڔ�+��C�Wc��;����+#�E��s���hG�����������;v��Uu��ԏ�J�to��7�w+�GG9��ːč�e�B�^'�d��9Y�O���sb���[&������8�@p��p�R4h������O�t5mc�Hُu#s2e( .��`�G���\SEZD�#��T훝��yPٽcgy���Q���z'r��&����Z�T\J�p�e���˖�{��	��;��py5�2d2B3��
�t����?B������nAeܽ�?.P��U�7�7�M9��f�ʈՙ�������O�!�/��@`|0�����.-��a����~��}U�!��V�5�& C�SW�n9������#<\��8�0@�>a�M�)�F��0C�b7���b��&a����5T��7��+��m���r�n�D��Y@;�̾�� ��9�����x�)������-�@�|���U>�W����;�<�ɟf��>�r�񱰙�lxl ��s���^��Gc��Lf�IkwԞ=J%���E/�}��� ��HGs��7������Lb���6Z+��D�r>e�p�M��Q	�a]���0�$���d�fܡR-Ѕ~��%n엾���Q�>�����.���g�>lg4@�j!���R"g�ϥ����9X{���r�D�9�\��&@�`��q__�L���R6o�Vz$�n����C��X�^v
��:"ti�W["/$���L�����WJ����7�������τȫ/	 [|���":��FX"��=D�h�70�.�0
���߬v~$�?Oc��c��,���F��<�.�C:{Xv���O+�=�Vt/^����N���q�-�v-�hH��ޮ������qS��KY]��/eFm�Q�UsRHD��7e΀[���*��J�`)ιC��n)�ַ�?��?�����w}@: ���N@��?R�"��DEA��\@L�hY�]��N���������WJ�i��3%L��׾�E�.���f�5Y�^%�C\:�H(J�ȅC����WA�{�\1���
 �O �����ay@��G�������Z.a���o�^���~��ڟ��g���R�����t�2*������
1O`G ���W�A]�DY_�#0�j����|�ϕ݃��	G�P~�E/*��0�[F�+_���P�@����b��`���	E�����NJ�k�r��:@����P�åyC�D�Q��8�fI�������S��d���_�z�K^�1�-��w�y������6l�j�v�b���B�|,A�1.O@9�R��Pz�Y�?�hū���T����|�3�g���7����;nuH�Źz�)�k���'��a�=�@��	 ��`��S��C�����o���t���e/~i�9�������hJ\�_�җ�7�PN�p�F���u�^c��Z!��Ө ~�� Ak7�9�ŝ�Åf��n�Hv�M�^0^��V�C�X�}�k�y�=߮�W����VQʀo�������E?�ݙ���P3�5�������])�s[������������������4S�G�K׈��\��q}�8�7�ֲ�@t�۾��p���ʋW���r�� �6��ԓJ<׳0�*
�s��y�a%����A�a���Gs��)�Pw~<�a�Q�;��7]S��
�x��ӭ�,w���N�:dG� �f�%t�(e�%�=u�x�_��'�jG�����;.��k	���NHfbbT�e�s�q��c6���S�i�>�B���(_a���
��� )UҴ>1@�U�pǎ��L�_�������?Ӯ�k��/UD�[�t�)'�e����˺Z�.�S+�+����r��LJ5�U�b`���Nѡ�h$F���?p�~�#~�C�+^���'<�|Y����u�/w��p��?$*����EB��q��&��RV/�h`�X�c(\`�p� ����ժ�m۹�,ʳ��[��������c ���߉���w����o�v���m�������˺�X����<?��0v1�j�ժ�Q��믻���#�ź��g�f�%E��^�Gv;|�;߱��Z%�2a	���Q|�+��`�\��/ ڬ��ss2�v�B�d �Ec1VKpt�ڧ� D����g���e��!	䟾�O�^\rɥ��\v��N���I�� �� �w R�ƜhBv�/Q.& �7$�������a�TDխ���?�1��/{�4Q�ʕW\��I��?x��������m ֗a�()ӯ�~�-��<rn1vu������jT# 
��l������C�:[����D>��϶�mo{��Z�	�spۭ���֊�"8FS�gk7$�`	��L ��{�3�j[�k��S㣠��0D�����E���V��;R��8��.�`<��qJ�Ԃ�0K��$�&7}r睛='tփ4Ǘ��%���`m984(09��P�s�r�qh�hC�9�rg�ah���Iz�� {�uM j��m�����+��Gʵ��Y2�kc7�����9�&)3�>/���� �0�O_�p�F�����̀
�A�N�{�[�M3��3���f排��ˢ�?�E�[o�N=�+��`, �U�:�zV���as$�X�~eq�$z�ݼ�B�)�`#4W0\vQ�����s�G<��7~�Y�x�p�1��/����o}K��eҥ��3ɦ�s�b8�X��.�;Ys�y�h3�E�$��]G�E��uQ2���4�v"��:�(�-g?��J�xC9��W)r��22�wlw$���v�T�G�Kn�X�3��� �G�?F� #���1�ʓ�~�~�������v��;���_��[7��~���ƀ��8��D�s	c���ꀬ�vs�(�:�g�V1WC|+ )��N�K_��W����S� �
:���+^�
�w.tDz!����[�x�� �s����LMQP���2YM\9�gK�B惎�Cٲq�!C����w(_�-�%e�"˙�5� �ח+T��5��mZI:�bOm(�C�
�+�D\7�'�%�C5x�~����׼�5~���9���?��#���W�D�p��)/C� �n��<sV?�D�֕�B�˔�q�>�Q����|�����v�;�=�O*����f��Fy�sQdX��E�ab�5��8pa�0.N�Ȅ�� :�s��ҋMS��ՙ�?��d��="�8�5\�h�.��b��>�_zu�s���p����'�p�7i��q�#��{��u� I-1D�T�]R��|v]�7ma�P��2~��H�:�(9�B�am:�]��֬��CC�p_��MS�O	������X���#-�~�z`�`�'b�	C��@�n,|�Z�겘��=QP��Yh��E}���>���6 zX�� PiZ�C���[�a�tZ��:�,�-�d�v4���%�~��*�b���r+����;/v���p[�m���ؐ#���-�'#�J߽��?A��s��\aoV�X�Mb���V6�2Z�ΪR���QIQ�"l Z�%���%���H$`(���P���<S9_��^֠�UJ������S�?($�O������T�q���J�8\`�aa�"�md�cTH�3�9��c40��-���1�?F"�#�R�s�dzYg�]�E�`�ey�pyE"N���yFL�<�P$^Υ"�ӝ��,O��':̾����w��{���<䡎�!�w�����F��|]���{�O�hv�2 ͻ�������$v��{/p"D��q޼es�V׀�qM��RGMP���q	0+��n�T�	�3
���#a��*Ր�:m �v�΢'s�f��݊��y_�D� .G5
ppm4-� ����i��2z��@��#�=n9W�B�G? P̧��x�y�JuL�����Qp����  05����M5�=fVt��N�1gYWߒ��.^��h�����p�gh�R�}���v�#̝���Ĺ�`�@0��s�B9B�؀*����A>�� �?&�C��\����&�Eg��LXƚ�:��!3��z���J⇵��g�C��(�k��:`z��el�D�r��U�����L�?6>�4>�'i����� �Fz'*�|��cQbMB)���	�7�!��Kc���H$b�db�p�r��+�6��qhfp%i�_ w�>�}����U�<�%�t���}��^q�ŕ��N
V�.,��;L�+Wh'�t�,����a�.M̙!��~z�����B�'����
<Xl�F��� ��)\7z9"E����T��ڽ��?b�M��~� B�ǔ��,��2��L���𰢣��.Eōi�I��ԗ0��O�u�K�=�x�8�
���x-W�V�c�b��	Y�=y�&�5c���w���v8X�{L�Hm�o�!���fW��M
�����HװOb���G�h��"�vi�	��V-'L$�#��#��0��*�4S˄��[���[2��燎�x������cj����fn����Q͉ A0 v"�2/�(�y�Ffm�45� X�է37�J}�X�)����> ߵ�|�	��@0N�MhL��qf��� ���2�	�v%$�2���A�ܙ���I[̇ ̐�B�j�ؿß5&��YȖ1��M���戂��q�����Jt@A�ٝ[��e�Ll�S'�7�&����1?�w��)�������и�g��>f�����ɕ~�p�r0Q�囪�G��cUw d��2eCs��Z�t��&���W��*�1X.��rNٛ6i� �������p٫��e�V�Į�r� �6"�#��g��R��ĸtO[�����5=�C��
pc2-�_6.������":�!����l�{r-���n�����t��9���8ޝ	����6�4&^�����xSx)���:�@�����&J���N�hOSC/2��|�k�co�%�Gdg�5��%�h��h10~�e�r�h�X�K
|�N&PC�@!�����H�����Ȅ�P�\�rx�������Y���)��\@m`��,��GwM��tT�ay�U�v�;֕W�F��y�m "x��6ch�RcJڶrx���.�.��"Z��1rfO��[ ��jL0�y&���+�`9��<�h7�@k�d��p{f��.��%䱯�1!}C�p\;�� pFj�0���,�4m�	W��M �;t
�"��j�	�]վ�G;"l;��z"Tֹ9�c;��*B�)����B_G�� �����\�9�9���!�%�W��F>ª�O<f�N{0���5a��&�y\tU��閲[G���?]{�\w	\q����dv��y\�y�e#�'�lK�=m���pvm@n�mh�iQH�YO�8��8+���K��pң��=�� ���l �k2��� ϊ��EYK�ch��M/0��s:r!��˼�T�*���>�A�%7�W��߇�����	�צyE-<�w�ޝ.��W�<�o:�E�Ş�_ ��ۍ�0w��˖�S��ψ�Գ�v)#�sv��4+y�]G._�~獷s��7�g'gf�Q�l�h�li�5#?Z�F��]��g[5�5�x&[�u��\-ad3u<���g���yr_��p��?T,���C���rO��"
�(jZY�t���{���\<Q�)�Bw{A�h1�7���Xd��#y���"H�� )�$l��`k�Ң�-���(�97)����eK˥��3�h���)�V(.F;��~h��P'���w�͂�b����:x�E�0"T�Fl�:t �6�&�ȶ���܄�g��a�C�̮��t��໬IDw�ؙC�[/T�C�&�7��nt��i�W�/ Z��Um��0�I'��y�[�Cl.��q�c�${=ae�_T-�� ��(q��e %��� ����=�F80,�h�ˋ��)-�h� 9�֌/@��XK��h|�0n62�r)�?�I)���+C�q[9^R��Y}�k�e#����g��^�gou��Y��*(��\JÜ:�t�eC��1��f@�4�W� 
���a���eܒ�3˨�H��kFPp�8��P�;�S!���P�,�+�}�o�4g`)���r���*1^ ����n���> @,х��}B[�,�cP��S�M"X�x�B�,}��>�˽ N�4`��u��^�vݼ����pO�7��iS�u�:�tS�
�x�mr��Nڻw�>��8����.�Z�����((A��I� {�;���_sF�kk׭)�y�RJ����'�)4�w�ջ�v�l���)��H�/^���/�Wm,���������W/Q4ٙ�iG�����jmj3��F3�E!�M�OM+��&Mk�4��0ݦ����M�?�z��kVϵbP\WrN}1-Q��9/�ֽ�+JoLc�8BJ���1)VSt�dOg���s�nk����6���������֎�aٝ���W�����-�ց�0e?�_]Ap�o�7����jL?�a�̏b��.�{��p�4^��:��O��4L��G�I����r�5g�bâ�]����
�;k/�=AB3��D.� 5Me��:ch��G*{�J/��c3���/ᦩ�A(j-fֳ�EHu��s��JhBT�=�:��a�n!i�v@ l�ݺ6:tF<��4�S	��u섄ڴ�s�7���w�n�
�! �k��tR���C�1t�c�}`Z���0 /���ON"�V�MW����`�~Kf$��=Ɉ��2� �4P�G�n�EZ|���?���I�.������� \��С0�Y�
&�����&�g �� �2;�a� ?�f�1���8�9���{�o��H�c����0y�q]��\?���id��9y�K'(���_���wf�n�y�d<�ېJb���$���;��,�#X�(&J�16 �F捿�N�Y�-昣/+S���c?��`J=H����b����s��/#�`WiO�DĄ���ql�~��LJ�"c�gn��"A"�G>�>-���V���WX�GAT������5�K`����u(���O^��*S��=��d(}�CU�1P�ʭ�3�� ��b���P���`� lK+�:��&�,���6yy$���w�q{�����ܵ+�ꤞ���|\�Be7f[�ȸtQZ����M���ilxpE�����VLu4��j�X�1���* �ǈ�l��J�6�Ƥ�sOb4db� ?n��-�ss�L���M�qff5�4��f���J�ߥr8����Q<��QC�y��sV��Y�z�����:����,���_Ѧ5��.��W,����]G�{0 ����=�@�������{ � A�OCC{x/���Z�F:=AP��Hbw�k>Z���i��`Ե��������\��oc3k�0��ᅒ��f��j>FCoe���������j(r���	uȽ�{�u"̹2,�wkDD��M��-j�S�t�^$�� *M��w�y�܇������V�<Dh-����O�c.�c$d�_]������^��9U0�)�M�D�Ic`�*����>��4���ۇ{G(�
ظ>�k��� F-`���HX�­�a�9ҝ���J_3��،��γ~z����Nc�ȅ�����`�5�t�L�}���_D����e��ڬ =@¿����2]p��o�D��*�q�@��xc	��c�}g��=i�pAu/ѹdx�+�����!A!mu~J>�0-h��C�S(�:�<��X��p_�F(�\R�N�`6-wF�q݅CF��<�;O�p���>u-�偙��������ј���`�_R!�Q��J�:L�~�`+��Ql�ꜭZ��T֫�TO4�p�_�V���\�A:K	�8�?ֹG�uH7$׹/�\h����n��Zbb� cb���K��2Q*�GJ||�[�)w*�ę���.��g�Z��:N��	����_9�Z �=��|��,�l�]��}@��srtBd_GG�ܧr����=g&pz�)�<� �ʺ��\ϼ�� ���<f��͐]����:�O,Qn)\O@�ǽ�,�kF���}���Z'��Z��o�c�_|�>��"�O�t�aW�vl��4�@w�%,��2D���7�	�hI.:<�Q��� f���صZ�"�Ц(���ף�Ŝ�p�B|����v���w�e��N������f�� ���&��!��̑��7�*�S�T���]ka�VD�z��n�i}֦v���umNXp�Gϱ�nA2O����Q&]���O��1��NLnTF����9G�ՑY�޸���������̦���ۋ�o[f�&$�����ٴ��R��t(:שF�sY�+0�F�Q@Zۤ��H����(�a�W;Ӎ�@1~2:.k"a8.�0�a�X�C�5���}���Na�r���ѷ}r��W\FP%+n�x�[�c�v�v�[)��[��W�^�q��>%�Fk\�z�]D��wiI�Ř#h���� ��M}�J����eZ�K6,����$Kb�
@��u�<ȿ���>���쇜Şy�F��ĭ��x8"K��ui�#�`	`�`3l�
է}z���y�h� �0�c�Hj(�����|�䠿0��7' ��좋�y��Q2�ߑ. "��6�{!���߸Ϙ��p�X���oJ��=�}�Q��R�8~D�d �1F�J�h���N����$�}�ވX�r��(��M���/[�s)G������۷��ؽ�ܶy�A�I����>�6$���թ ����x����H��%K��?��mV�f�VN����Jsrv�E:������z~,�ieIP�X+d����1��ߛ3MaJ4k]l�&bnvttnrj�����Uϑ���Y=6�*������Kc�{��&�=�[�>:x��\�c˶m+{z���t�MԿ����U�����[?��( ��4��!�9����[�Z�o�O�n�6PD��D[���=� ���%?�<���`��o"%=zv�l���ʲ �PH0�諕;�a>�lP������Z�0���h�csy1�
����P�ι��*��Y��ܷ�'�|�$j�a`6�^uY(�b��ϭ� 䗐n]�s��`�O�.�R��>�5����hR��<����f̽A�� ��,�����i�k���s��n�-s�F�)B�c�4�����ǘ3�{��¬��^F��,������r�l��s}@�@���c�(����}�ͬ<�ݕz�������+0)���x�h>Uu�3!�q?�d:���s�8X<�\�+�M() %��v�c���܋��ȿ -�Bg�*��U���*�_}nh�ѕɪ&0H`k�	]�@��Ww��F�4�ݷ#|46_k���d��?�\g<����#p�����ɰP����F\�&*�|U�7@R �n\���c���"���X�ڗ��.�-���2N0�Y0��ʹ�d���pUF�
��u�h?נ,�Sq�ޘ��^vi9�ӜHQ\ߛ��|X �(������;����w�( ��v��Qe�7��nO�t|G�ɛ4�lǝx�˭t)�]�=|�yڨj~(4��Mt<��r�)RlF�.�ы����][6�ݷ�i��hZϵĵL陚��gRB�I����x�֚&�f�:�U�\i3ۦ��o1Q��L��w�A'W	��ix���M�3y�	��
]��3׻l��1%����t� ���Z�w�0�\Gw����n~럽u����*o߱����bݿ�"��u���9�hT7Չ��4U�?/y����7'JF�З����G�"��qg�A>��ߔUD��9�R�")p��
QY��â�wn���+�b�@�*i����L1n����ؑ�B"�v��O���R��0FDaq�v-�?�3,��6x���&��:��BR�Ӂn� 7�lZ�5�t��2PD'�7ax�c�0l, ,89g`����ݧv���0�ܻ��x����ݬ�.=��#!C��r�z̓=c� �H�<����x��y�.��Y�p|� r���r����l�f�[��O���ܗtvi/wV�����iCAfv��ĥ�{��F���p���	8����ȅ+��0����%'CJ�)ݶG���> �ǐ���{]d͚��א'���s��8�Ϯ���ܰ[T�(�P�J��2v�T ��V+���Q��Ԇb|�tP�`z4�Z�#�"
,���5N .�?� �!�$�B�n��Z�Zc��U]P�q�]����'+U�o�����5����Y���Pb��zZ:/����02�>��0"�sa��͑q�0�r��s^!�1�g8�&�m�Z[z� Q��"SN�A3b�FT��4�t� ���޲��b^��
��OP߂kRm��r�-�O��r�
2���)O|�T��(�ץ�1�N���a�t\�Sd�g3�9��}�� v��Ng��3�Ƌ~#�&%zp��k��HC4���)J�g`�&��ظ�5V�]UZԗ�
�z�����Ǟ���֦z��I^ׂ�k����n4��̤��M�O���7�� 6�Zg`�b�0i�]����"jKԢ9�K�jh�ĵ
�=��U��.�@�9m<��z�dwWOc��=���7~t,���G�z�v)L��b�5�'����_�ii���f5Ɖ���t9���ֽ /��7�n4��j��XDxNà����"AZ��u´�A��Ov�z�j-�wo/k���#N9��ɸw("l�έ�̳�p��	r������/�4��W�B߮��42Ƹ�X�i���%J$*�EtF	;�ZK���bZH��ު�\�����l���)|'��}���]��Z�`�� �'��!1Ȅ���h@�o1��++GB�9��^Չ�G0���`mt���ݸ
���E���M�� ��I�"�}�]$����lۈ�act̰�H���U#ѯ����U�(�}?��psoD-!���*A����0Έa�*
�93�zU���.%~rX��^E��ݍ�S�9r��xh����hK����׸bq��D�@����ɸ��$���#I�(pe������d�k%¬��Т�x��,٘� O�h-��.N{��\/0Uu�^&�A ��{l�yf�"�ML�*�@�R
��d���2�#�>� � N�����'��eH�,1v����>E��H@=��`L6�jd���'���$8`*���f2{6ü����L�r1�)���;�|GlƜ��?���7d����?R#�a#Z�y��P��=�y�#��ی~e��T��'����(��L�Ђv�$�=z6'��0?�>���
�ɺթ�3l�p��z�i�"�]wp�U�+��X���ʯ��T�F'٧m71*�t�y�
�t��;�)�b�5��ɤL%�-�z4���MO̖�#x͊��҆���2.W5��1��R韶�ܫ9��)�}�lKSk�p|��X��yP�C�y��e�k��E� ;�#�]�"3c�f����\@�H��c�RT�q��%
`¡l�}mN.��Np�hK���p	̃�
�,�s3�Y�q'��w�_���r�QG����o�cV��=;({�]��ǚof����R��L�����-	��A0�]�$( �T�I����j�s��|�u�T�/"giFt�=TmJ�S0g��c�(']�#��)��ΞϪ�%Ȍ��ܩZBv� N%��� ��YÂ�'�JF����p!dY���@�����[�0#�����$���ƫ0��~l�z��7>F�U�9c-`kw��.�pO��=�q}*J;��q�n0�	��[��t�����C�Wא��4qs�#�O,g�q��!��Pv�T�W��e�ve��Q��8o���U��\h�>� �����qF"B������,p=3��t���6�Y��2����e�gTs!E��'��GG���-�0_�Լf�ý~d���b� �r.x6�{0��#ڐ��|F��vPi ـT�84@0��>�jm�Keu�l2Y�!b>��m�r�hS`���r��~�;���~�Źs�nϣtq�e�Rϻ�
Q�B�X\�f�6;�R.�f3Y�}��$Z�V>���(����Y*��y�:�@����pX��W���wP:�f��1��?0<�~��9]�X��d	`;�Y��Ir-�'h�"���f�������R	0�c�3$X�C��X�����53>�?�|kGkK�X|�T�����?�r�n2�]�Ъ��{��;�Wa����>]�G4{�y�W��3��id�Y�M���e��/W��������׾�\�;��}ʲ�\��]*�x��%���K���͡�����,����DF�pz�����0���+�/�S���a+� `r�ȖcYd#��Zb~�|.$A��7�g�`h��qI�u������LFHi�
,�%Z�~ff!�<5=nj^R?AGd'k�*��v�~j.��i�ÛkVh���/ʲ�<Q+������V�j�|W�J�3p�ErJ��{`���|�`�8b�m�d�Ȯ����"���T��s�qB���P������ɪ
������gq[�}Vn ����ӧ�#l
cn���v���2GM
j�KΛ��J�LH��'vT�^�i�t	�� ,��� #���滙x0�gy��MWZ���vr��L��85A@��q���\Y�H�8>��l}�w"�s0Hb��.8�8��Rk�nK�� (��yfGs�,�\�䍸�����g�O���<��#�$�1�(C�������)�>=Od��(�&J�gZ�y�;�s��5�D�� 7�A��h*�"w� ��_d\S�P��=�
 &oD%2Z��C�q�Pр$`�sS'�tR`~�V�̵�?�,/��y,��� #�2[�W#P !���i�����6#C��<Gw3O6�h��(8e��kWHV���A"����MG������m�*���W��R�WE�[��lF��\��F6��:44aT�
�
(33Ca���`f�pD9�����`���� ���,�hKԧ�D�F߷ؽ%��D��M�^#�j�4<'j�u"jTjH��rB�q;M@�A@��:v�+C�3�s7������ �C�
֊vf����
p�4�}C����eU��@w^���Z;R�5����C�Z��6�Uw��V(�HF�:gT��UU~_�~�ڲ_E_��nh�����?���I�@ ,єF۠
�%��V��S���:��#���V@�h�} �`��1��J�@p�}�Ѵ�#�^��>� b[�6�r��E��7��r����ՠ�K�=/�`��0[�@�v��H��2B�ӦM���n�%=�Pw>�Η:$Y�W2I�+���;.Y����Mmwm6mn�h�8S�����LS�?�7�s83�f����p�n�\K�9qe�s��o�UN�fm�V{~nSh;l��7�,�nf�߰�Q����{��O昂~"=>����b@�(�(o��$�JY'���"�6��Svj�6�s�g|Vc<���-��9�_?M=���h�4kQRГivW�F	w��ŧ�:U/�Uא;�\��O3�n��O� ^1ų,E�� ��������W} �%b�.T����
�d\ݠ��ZyE1I�R�d{�6��{e�:��>@�i�\�`D��ˊc��-'��r�ͅ��X�����~r�r����7�u0�|�����"M�2��8��HC��(���1�ac�lE�~����cXls��龎��n5Y'W�;\��PF�OV'ٝ*V�Ҷ-��Ic�ƕ��}\/K$0p�Tƭ�pfi�"�q�Xԉ#ÐEdQoB�e���p��}��j1ͽ��ۧ�7���q��������A\j?��-�N��?�2��[����z߂i�	lٺ�!��Q�@_�`�����(����ka@r?B�����L� �t��|�J1oӵs5�4�J����c0��c��W���-�E�'�g���"1��<���H7����T��̈́�-T�qnBpK�EC�<�.��K$�H�|��L��������:{f�A�uE};�,׊�& eu��>�t�9��>�ktЛ���!!3����;��c���UXh/st떭���.��Uש���Dc�U���ci��޸�C��Q��U�Ba�N0��P�ճ=FrC2�K�?>AnJ�Dy!�4�"TW���_� 聏��@s-z�%'q"L��w2A��n�L���댙���J(�P���w�-��(2���@X�b�r��%"[/MQ��\t35���ErP�-�݊���]gr���AJD��XT���Ż�LU�٢��źJ����k��b��pa��
� �%��п�{���O9CH�O��}h9��$�^�H�D���<�h�������y�Qdqo����ܹ�~ K���-����>0(�b�Ƌs`4�DaT�!X	X/"~0�yO�fg�7��)�e&��nk���xF��
;�yU�S�g����01��+U�;�9�C$`l|����w7i'����_���d|�\W�Z�{�XJR>�;'�$y���¥O
I)�:t�sNs&Y�dW�7�u�J�M��Ƞ��'�K�{K�"�`�s'��\++�3W���$�LSf*N<�$�1Os�-�U7�`�1J]X �V�[�6	��!�h����\��$�*�/n(߯�a %�(5<Q��N�66G���\��g n�("LٍА�π�d2�����ϙ�����=߽V�7c�w9c;��]�x��;KE��>�Liؖ�y� ZbiF�<�g��'6!�&�#�w�{G�Q�p8Һ�N�u�8���Ǖ����T�C��Q�Q�G�K��_���m���Y��7~����6/���� ��W�`U���Ñi8e��F$Z[/L!��>��Ǹ��H���k���n9�-���.JbE��*�t�_ީň�M�Mc eo�n��7lX�Z=k��v�̳� k2q����ga^4Q$3v�ro�#EN2�F?o7���#�3Z �ó1��� �����v�E�Gj�>L�;`���!ȕ��r׎1d׊�)w�!�U!L��5cH�<�����qs��w3o
;e\9�M:��4�
F�,�@�T��x�u��GD]���	��{�J�����v����Y� 4C�3 �v�H/U���Ũ��Q���煱A�f#�Y:JO��e0�#�0RT
\�("MȰ��w,��U5>�1�6�
�� �>�7�U��?�c�'@Me��F&4APjz	�wj�K�2�']�K(j[�g�z}V�t���yM�$��|���&��ۄ��|&�0�Q��qA8��H�G��O] ��AK���=��މ��꺌	��D�K3��]�^��p��k���2',�w [��;6(�+J���L7X�9E������/��9������˳����v��իW��N=���S�R����9�xDy�k_S��ǖ�|��J�y�}µ��)�7�v�o�ʘ����v�^m��sOt`Xd'����k�1UDf�@���4���ch���s_<�M,F�=С0�A�Vr��� bծ��6���ڨf�^�|/ڤ�����!�uxxB��Ouun�7�̪��f�0���#��L��8(wҖ���	ǝ�]3�iІ���0a��2�-��)��i��\w�,�)`�d�C�)h-Ad��Y>��z���Øu��Zh�m�x�MS�$����0;>/�����!�����i�K?蜸N u��a>����
�:)�9��)����U��]��R���dE��;l@�ݡ�Q,0r�J���T�B��( ���g��޽��h�Z�	���Β|0�(?X�HD{a0ƕP�	$ɩ#P�ѡ?x٠j�$`%�L�Csn3B�`#�k�N�b�uRj�m�Ů��r�۩�NiX�e�n#�u'�7� �Kԝ���b�rӯ���Ξ�&���|N�0��F��Y!�͈�=�BN��Y�q�y@#�E�����@����D�U���	]k��mkF�Yg�4�h���r-�1�FD��� <�����NX�`r���W�缀j�)-���A���xv���W�˦�2 �am���^�(���oh�"zrґ��@5��ɒ��Z��<���F4\��lh�x�6n�hWn�n��|�K_�Ɖ$�0��+��ԓ�)�>����_Y�<?�ڐ�ls^�,o�\`M�2.�aD��\���U�(���i櫊�����En{��]�4cc-���D�1<?��Yd�����R�����1�.<��|8��<P���6�+��d4X�����N�x��Ϊ�׈�����P���"-�9�2X, �S�}��E~��g����bM��1�����ڐ\��a��®��r�	� ��횯
���'��Yޫ��H��L�:/�G�5*+D!Lt�v�]t�Q�h�p��06`alc[�\ 
'مԠ�&q!���E8�1��['�S�H�ƥ�<��g+Zg�<k���2XQJ���|?vOx��0f҂�	��ڔ��/D���Y�7��q 9�+�_wݵ��~�.[ج�PqJXv� kv�w�q�˯�_���j�	���X@p��W�Ez� ��H�Sۓ�FF6�]?v%����6pOb��7���<s���ΕA�mH`�����xS�Eh<7A�|ޞ�R����4�rY����zX:�(�B42�1ܼ0B�9�XZ����F��7��/ܓ���<�!ժ�E��z̨ P���l��L�Y�s+]�#W����bc��s�C_g:�����W��o�Vey�9ڬK�|���eZs������n.?���GM��/+�����*�Wܴ�͜�樲��k�E��sĜ[�k�5���J��ҥ~�����H
ݦMذ�	�&kڬ�Yڊ��{�������c=��=ЮtR�l�vyAw���6�G��J�BR|���QߋE6���"���>�ì<�9�*'�t\y럽OƎL��%&��uʀ���g�񛔊��r@I�f���F
V�Z�Ij9�P��[O�sL����?�]�8�~Ȣ9.��@̋�h�q\�
�05���6-�U��1eOypt	�>@��!3�̤�-�U� v&5�����S������@��<� WU�L{�ݴ~�:�ÕLF�D1�3�(��_�$	/���Ds0T�ci�[!H3`�.3�- ���Ťy`�̶	a����D��F��BS�4P���{�SN-�|�#�\@�h)k֮.6�P��\|���i0R"Cv��1H���bu�o�=�	a�JR�t(;�<��<=	�2�<�I0$	R��ioj[�ա���Sp���Q{ӥh�۹�3E[�MLA2T��t�W��"�/�QE���Q�|U�ZD|����4Z7Ui����i��3S]�m�o@1m��7ne\n��ʄ�[�d�\�J���9���r٥�5Ks�ǘ��H �oc��Зըˬ�\�ṁ��5*���Q�zT������E1�w�G>���g��8��1�)�M��ct�ח�|�[�K..��Y#fH�Y����ISVe��)��O!܌}$���T����6:�18��P��
)�/���p������w/������{`=�!d����f��0v�0*r	9��u%��]���}���K������H��4;uv�,N���w�W^U�Ĺ2��2� '"@i�¸~�r�-���-g�ur9pp�CT3�cK.�I'~l�=����^�Hw������cw��L9�`N�/��<#խ�;�f�G�p�TF$�H�q踒�Bࠍ�٥����� 9��ΓU�'��å��"�Ti�w^�I�1X.�!��kV�I `>iu�� ��0 �n"�"����1��.�RF*"�B�E�asn��V�2c4^��K�>������$ߦ�D�;�\�h����s~c̸w�'�a���`���qS ���_��cv��c���'��Rf������~��V~)D����r�" 9�1��ZU�`]�%�p��U���`ب�΋�ѷ��i�Y?��Z�ψ���չ�wy/s��2`	���[8c��H2�G� ��Z]ɶf	�d���cT����,����A���"����wfm+��g����)�Y����3Y�!ږ�,*����r�E���<�bA������o��Z:�`�g��.R��b4+�:��>F�=:sA}Ja҃҉�~���ѩz]/|��*2�h��'�ɹ�����a��5EO(/~��#���򊗿����Yt\��0���q�	'8���n��e��4� �c�=o�?Z����VE�]q���_���e��3i��̡	Z@��i�]<�ǹA�=꿨΋VEi�� �h0P�����GQ�f�%O�B=�z��i��Qĉ�,ɸB֯ۨ��l��=2P�BZ�ĨM��g!����.���N-g��`Q�se�����M.��AIڪ{c�n�/��{�Nh�)�@z~���Re�Ɖ�����:K��J�����#�� g��5"Q/�?����i���Pu?���u��jakR1�cd*����ݫG\Xfd�kE�+�2�	�5ە�vF@�M�t���0I`c<�q��4���[Ɓ� �I��[9����]�i��/\���!P�M�Mԗ68Z�'&IN�NI��8AD���#�kF��r*�@9J�2�|Q��4������;��A��%�|2��.��o֣�"�*��W+)�Iy�����?�� �e��O/k�V�[o�Q��l߱]�n��a|\�Yms�
x�U��O_r_f�H� �&�T�)=�6i��>���vQ�!��v�7�C�D������h����~ m/���$�R��Ƀ�3Vh���x�(wrG�,:#�H�j~��[G||n�#t�y� m�ڥ����� �́%r�ڭ�����oص=�}B�ʂ���p�X��%��Pb���Sm"o�����,`�Pץ�v��{W^q���A������S9=���^ JPKK5v6*���ٯ�,p�c�=�J���\~�����C4�L�{�ψm:��%��I��lV��K4�>��O����-�~��+_��K��?��ҖY����z �{�E�:�@O��LMj�#uv�> �r������J��).~�]��-�+M��Ӫ;���J���맨A�l�Su�f�iղ#YT��`��Q ��t~������0^	x�w��7N��<�ܡ̬��EZ5��e�\&ZԦH��«�ӊVg��,�nW���ejh����r��.[���TX����fCX�����
����~�9;�Q��� ��ݞ^�?�Od�KA�0u2�T���&��	m�� �&�0yp��>MV`g��Q�WB/�vЂ��S�	���D�������I*3袴��w*�$��Mclw'�E�!-�T>GЬw$�kՂ�ZJ]�)�c*Q1�h���D� ����IQS�\�]��Q�t��b:'F�Q�P��eBQ ���մ�$l L�j�\c��/4#�+3C2��G�&�d�. |���
�?&����9Y��0W\�}e��ڎ�����(�E�D�U��#�в�#����^:U�Nî(E��!ͷ�졿i>G��I��0 �Ax�ߙA�5�Y�$=KRO�{��i�8�L}U�̙�a�@�%���!�+�v^�
�8��Ts��f�/��artg\3�c�N�9DS@�1\���� �#'�$\��+!0/g�gKĬp�{�l�W�4m�UD3���1.��
�d��X~(�
��o�"!�� -�N��ϪU�a��y�� C�U/�~]g�F	@Bl&\��`������V�u��w��{\��[�o�<`t睛ݎ��:��x^�6�c�:ʐua�@��?��_�%�ξ�q�3��H��D��K�lN� ����բx�;4��XݹT�\�����ƕ��6�̦��z�c�l�^���fT�Q3.H���OI,
��@������w�>�GP0?�.5� �w��,L�>����Av�i������;�;et,��ı�-c}��WK�x��]i4��0�.|*�3���2g_���D�j-غVc�EDQ�a�=#�['�0Q�
��@��9g�&��ĝZHDYc��
��e�\*�Č�/:���hV�'��r	s׵<������;P�;v�>�G��4_����@���!�M11��1���8z�� ����H.\�m�jf{��]@��Z%����3���,����T$6���r�KƂ�8?Y��sλʜk%�2��c9GQ}�Q�>�kP�_�t��#�BP�BE1�ލk)KJ�^��-yf1j�u����B/��0��#�ÑV���uּ����c���֧H���)��ӟ���ֈ�Uø9Ÿҧ��f���cT�'�&=��;����I�����m����,]�����q _N����:o��,���d�2.A����3�Z�y��:�s�2Wx���#w"k�W����}���p3F��F��mN̯��r91/�C�ںu���o���.fͱe�Mv����۲e��'�VX��FV�S`o�����������g?�ܥc�D��6	���ֈq�Iަ�����P�%��Lu�Z���cr*�h�ԥ�e����srE�j����63+�t�Ĵv�����Xd��Pk���qF2g/TwO�SC�z��a>47P,���`���$٠F@�2��⸅���f��"F�G��Vj'�e�4�ٶm���ڡ�#.~H�v�֓ஒ�b��S]�����K .���.���0z�J���]��������3�3�?����"�pUw��@������am��`42�p�p�D�.#���A*ꅾ!:y�|�fP�=`90��YD���MF`���,_ ���x��j�0��Y��d|:Čp��)��l^��"�a��\fc�Lک1�R?��Ȱ�����j �=�po'���!HrC��EL�v�s �0~0Im*J��o"�\@-M�$h��y�\ߠ�j���*�9��"��<I�b9�H���e�{�(,��'C��鋨���&���1�莸��?���K.�:7ʙ���k�Pi�s�ŭ�*�
`g6*�;�!����X����ߝ���'�4�eɌy<�S�@Jn\|ߺg\�fq4�̗t�s,�9˼�vtY��6�,Eep$��eɜ�Ṡ=K�*���&�&����q�b���B�\���.���D��>�;���������*aϾ�
|X�qnes�g�6�5-)�;UFc >l������[����|�(�77�8.����Y�i��:�1�S��	m�ȵu��t� ��sIY�98t`�R��-�sJ}�[qh�hW��T_�r�,�~jz`=����W�uGIT�o�ㅕ�H��@t"Qk#�� h!,=@ͽi�o0B7s�8ɞ��~�4���Xt��#]8�Ek%�UT�2�(P�΅h��e���d�V�X%�a�,��]���������0%m������o��~�ca��,��Ļ��棖��.=v�D��sgq�dօ�8F"C � aq���F�v���E!�
� �����L���V8"H0��6���C|����rX���xA_3���v�Ez��q{Tm]�� 3�]w��Ԕ4F�9t]F��s��.��,ӌ���-]nvg���b�*�J[S���8���D��D~ M�j�j��0��Li��VsF}�+��_��U��	)q�ے%��A���=�f�-��7�W� �d�B,��X$�\����P�����\c��%7-&�̃G�P�y�7,���ǚ��ZX�
�/� �|�_Ѿ�}@ ��|�&�L&7C~�v��jɒ}���.�#}��hf��v�7��{�$��h�O��	�U��ʹi+`&#iS�"><��}�KPdrF洳,70���r"D6#0�r+:y�ژu����f���y-�gnV��}���v��G>�b%ʖ�p1�g��
1@��=�v��~�ʿ���?�g����I'���c�W*�ǈ
�H��G���H��m��)�i#�Z��%��̜D�곎)"k��U˺��[�p{"/�~*z`=�a�a�;w�O
��:W�.����?�dq���o']f�+�Ʈ�gk�L�^ AZ�"���uk��O��ʄ��@Yrک��*`P�V�ͬ5�@� ��5b�"2�ňE���v�PqF#*��*�E��L���!���K��'��8\��QM���P`���U������M����){vc\U�[tt9��m�C����'�BAi�9Q5( >G���bQo��2#��WWS�aq��ާU��i&fO��ŵ���^p3�c�!hi�+2��t�"C��������$�CB�>�Qu5���6u����\ �&Z�r��n� Av� ���X�W�(0K�c�8���x0hcƵ���K]-���<��
�e��g�;~�x�"1�p=5�E9�p���-C�~��1g%�ձ�K{`ҍD{x�0��6#z���t�.i}"�LI��p\5�\��}�^�>�3�<�,P0\胂ť�N��3����&��\��E]�X t� �rʬ6�" ��Ͽ���|R����Y���Zh�̮DT!��T�	
��ؽ�`�\D�؆ul��?��C��zV5�hF���.�3Z��Ҩ	���[�~��y���Ψ;�*A��q&(� '��Ji��cܿK�{��n�x�*`c�\_�֬пr (��-�3~QI��կ*�\v��SS�L>T�<����(�LrD�'`ը�kX�B�ވ�c��ٵp�z^Ft?K%֢�ڰ"@�5-]�jtfr�@����w/���]r�T��-�� ���Y���Uy�֟Y�Y�o��̂7�)�д��S��	M>�xI�Zf4W�[�~ǏW{r*���g�A�m�ņ����{`=���|f�MYT��
� �=
o�O^�3�MJsɻ����:�)�F*5!k0��l���qtJ]�x�Hd��"�B�e�G�ƈM�NǢщ���
k�c1����e���!�"�R�#�d��Ι�cM�0<ZP� [N���L0F�2���K<����c9p��`���h�!�(�����5������W�#�\�M�a��y�Aمq����E�+Y�S�@ꬹ��;\����r� ��:�uY�#��53b��D1J ���7 �SQ-�p�&��<�Ŭ����G7l�·Qw�o'�����,tAD�	`�с��l�}�ƍ��E��WJ֗�aE���5R�X8	_��/hς��� A�7�[�Ȃ�5u+Nv��K�]'=�#��~�̒e��E�ʍ*� ��#,�s9�:�b�0'-b�U���rS7M |D����]�k8a�A��2�[l[�P  @ɐ�	WN�����(�f0��i�8�L��ܣ�վ���Z΂6p_��h.td�^|�"���Uq�D�#}�����4��k .r�1��Y��E�zn"�G�Gb�I'�l�\g^u�����a����)�5\W:�BԪ���%�;�Ĉ��RM� ��͹e��}������.')/��&��(���W�^���
�ԫ����R���Ǘ�T/��w��aH��λ�,�����#������	�SoUj�j�q;v�(�(���_#�NmV�}[�P/`ܳ������:[O��;{������˛;�:��`�Eji�v�1��kij�$�eNsxNk���V 3�-s��Tb�	����M�ݏ�� G@�� D���lJSlR�������>����뿲�[��њ8��Eӟ����4)@E������9=�S�ө�����kVi�劌Ea�u�z`ݯ�Z8ؘ�A��b��
�*|��+�`��{,A�}��	p�zj
x/ĮQ�'�����&q�K3���hؕ��c��"����6�v��τ ω'�\��DVZ��֒c2=��H|hL{ئ��&�+�a��Y����p�NWN��|�u̊@�u�rp�(���*�����W�8er!��*��P軴j��pu@��dKs�����t�R�� �Ѹ�����������.2g�óuo� }m��E�w��K�F9���7��_��dwϹ�_x����z��ﳋ���<~�?jv�}��U٠C�j$�f�K���` �B0r��qfgC��#�q��+5jo�r�,�����?�?� P�+5W�b�v ����C��>ùNu� I���+��R~F�p��0&�vSٲm���׳��dy� �N�{��;�� �s��="�l�u��Q㣎9��*�s�]���`�)^:�9�8�}�&
4lA������quz|��LYX����I��F`7mdY6�ӼD��C�����a�m�n�-��M
�1��,��A�=Ǽl�$E�C�2���F*ܖ��(M]�$�ݻ� �����s��\�\Z�a�>p�D\�z~��h�M�s�"�G�[ν]��˵�{$���䖅ɚ׎i3	c����i�֮Y[�R4٫^��r���f�X �$U%���6Z�s��ru�ީ������4���=��G*�gl�4�.��Gu�+�c�Ԏ��]G6�]���ܺjzjNI�ۚU"
tV��g(;J]6�����'F�gD�"S��bd���5+g��h����>�Q������8���ig�qїf�"+��m��r('�{����n�K6��o���s|���`��%7����g���B<�����=���kO��q��)��h�M����G�S���Xf�m��I�f���E&�;�h��Yw�)H]����@Mf�#J
@4ƸG�ݨ/4"��~-<�c����8��^u�D�BtV�_֭]gC�%ѻ]7����8���*�}(�����8�M�\\��X�p�5r�`�dW)�ߗ���J�xFy����ъ0s���.��)��!���M7�����-Ĺ��Eb�H�!�Ɋ��.F{kxԖ��dD��|����+�(�y���6���0,�c�A����Q��N���kVd���\�R&�����w0�>�>I��(w�~���]cD����� �r�-
-W�]p�bV�6co�	��xp~���Gm�a��Z~t�U��`.���$� ��AEf1�  ����_>��f�֯� ���2.v��[�Ns3^��}���s��E^��;�ӌ���:r��&���:ѫ������7�I��G��n��@hㆍ�B���g�
��B"����]C9��ǎ�:d���L|�3��&���3�E�c�s�?�Q�C�P��[��Y~㙿^���'��3�U���ed/�L\���)C��.C�î`��toW\~Iy���]����w���������̜ݠD���3i"Ӏ�O ���)J}�7�"��[�m+���t�m�(��ǟ�T�0�Y�9�!��k���7�5C�l�sK'm����:���.���O�Je>�����.){� ���s(Z`��z�H�m!c�s��bZEkOw�55-iokY��35;95�f���1���l��� �\񘅚_Զ@
?�f�=�����Y.�E ;	�}Nt�z�p�U0������fm�i��V�Gk��ά$	�W�v�ԉg�~��yȐ��_�<p�j���� �0�&��Nv��%2�f��?�u5Z�����P%J����y�����묑�p�X젆{���W䀉�:<�&O�X�4ȏ��,p#2��+���'���$��|��f��ŭ��hHFmH�׺#�Z���P,���hwyAy�;����LYٹ�>~7��S�d�H�oq��� ���4�R��o~�k��^-���T�[���jg]~�[�Z^��ז�?�g�nw<�mP�A�V�C�!D������ �F<JZ��8��  E2EΕ@sx�L���o�zWWw�������,��?+W_s�2%/�B�Ї>ԟ��Iב!�0��1A�=A�Z�'��re<��,�N�`���'�]r%�������s��\�<q��g�"xe}
���c�D�fs�@���x0������p���Y%�H����}�/^��姝rFy�+^Y�h��S@l ��LCM�`.�����z� ��/|W9�|Ԁܒ�����O˿~���ŗ]\���^^�җ���)e��@\��2"��������1F[��`&����Fr7�����gRWn�����<��ǔ��;O�㧛����/?����)�_o��g?����d D�.���[�顇�NųPۑ�B7�3G�VdK�VN8�1�|nڷ��m����"`����/7(�0�[���T���2 G�FBH�k�)�9Aw����t$$�6�80���	7#�0md����;��FH�<���,�|��5kVK�����z��t�4k�7.�q1T-]*'�k�T}P��1ԦO�1����隉���o޶�����O,l���.=�$�?K��sP]jQ+�ӡ�쇤�U�_�!���Z$�-H@���uJhJ)f%�G�꿦q�,�\[�d�@��s�%-�[յ��Uʋ��&1�Mڔ*�������EΌ7ͭP���N�ؠ6�A!�\|ݧXA����� ���Q�U�����L[�����l��W��n6j^EG��W�0�6�����ʿai�\�"�(��:���)�(Hbh�5��x�1�S�u��Ț�Bn����b���t�A�b�]b|?��ϗ�k��S!�'{\yƯ�jy�c��0Y��S2ر	ևQ&)�}�-�_s
��b�Fj�Ҁ(BI�w��]峟�����[F�Mox���*��c�w��Ю��~��_�N1
J���-\��w1,�M���﨤�9�h��\JΆ��~G׃��U��O}�S��`����7O~��o��o����P�0�s��7;Tw�����6n��1�l�w�(ѝ�9I:v��7,��_�:�A�Q����z�<G�v��U�o2`��><��$k����9�*���R3�p}�D���[���1jGy�J9\Z�+��s_��tZ��R~vy�+^%��,3�DQѧ��l�A{QǨW!���! HˬD�	Q7	%J�& �(��/{�����|�|�k_4�x�@ �����	m�/�5�3�� L(�}�.a"@�ƅK<\���nUN�}j�E߇�OpG��QɈ��/��Mo����/}ы�o<��]�d�^%��;�f�V;�ě���E��\	�����v_��.�j<b�._�W�����{�k�����g=�\p�N�@0ޛ����c7��tEE�f���EFޭ���&��Q�ct��ro�_��<C��==�����(�'��D5u�n5kss��ʎ�[�B��|:��qf�z���v�Ye��#$|.eUg9z`E�_�Z˞ܾSh#*�y���F�ygg�Ԟ��wL)#8���ۥY�Җ��`�R����t��^m��8�J����R��n���C��
�*`Ӯu���Z6ϵw�L�(�F��S,LO/���X��4ף��hS_��ζ7u��gm�T���x�C2'�v��_�� ���Et��,����0�Χ9R0FD���}���>�A	|r���?F�J��Q1P��F��2t@�����@`!���U'O�������ߺ��{�x�i�'�F�ta���X���u���r��w8iަ#�*��v[y�{�S�p��	�7�?����'?�I�]Kz�Bʑf앺�8�Ǹ�u~Ƀb,뽭�?ijD���0�P�W��6�����˵W_S���w�?|��G�5������け�#v��=�U��]>v�q��f���1��Q}a��44��	eF�WYk��|����r�i'�����=�}��l�S�����W��`�|5)(޹c���:w�I�9�`�i`�'��:U46D�-����s�9�%/y����֝[�>���O�����	,�r�-e@,X6�����Q�,U@��o${c��@���@қQXV�����ٟ�o~�>�)ǟR^���_{��wV�����}2�u��l�"MX���H��T@@^��WEA�
�Q`���.�{6�d�'�$�������s��$d���/����i�߷�{��<�9�9G �Գn��qt4REc�����5ϛ�= x�!�B�㔜VҏyHB �6lfֵT�<��ԭ��qLz�m۷��o�)��o6v�+_��i�V*,v��a{�8���"�����X?=;Vh�6 nm��B�T|�WB������U�
��mo+�v��!@���b:^���/|���"U��ߝg�Y�d�&m#3�� ����(�}�`.ќ8�e�|�	������2=���?��Ŀ�1_��/��������o��y�p��sŚ5/�{�C��uk���M�'!ǂ����=�ۤB���'��L��ic���T� ��ฺ��:�4=���h�l`S߯\��2SYkv���j�$�j��~��B�BQE���6�Y�\��='��:Ӷڊ3��^�׽���?���Kw'~r|pH&'L:M�s�������$C�$��=�mzJ��(-oa��2}t)�&'���bB����_����$N�Z�ʻL��C�@A�\o6�a�>��Ԉ1���DS�E����m,4��B�U_�ܩ.��-|�9��8�E'�-��N@A����F�~�����[K�����p��X���b"x2+)0(G_��2����1�P�#6}a�:�WT��ب Ԅ�}�R�C�"��{X�������Z�<�L�?>��Ϛ�MZ�y�?����#4]��j��эZ��6�.��b���$����6{-jHN	'ѯ��ze������W_}U���ß�����Oz�Q]��o�-�},�
4�Yt�^�M�@���߭��uFX0��# ��m�7-�����Y����uo|����p��x
Z���������X}�.U��RJ��ߔ�����`l��s{�̨�2mN�<s�����Έl>k١Ř6�~C�z�W�c���\?��O�O�&�(,��~8'�ɣ16�i�TNF*����pČEt��"pxpƷVh�jE������r��,:BcmSذnCx�ަ0���~�Q0 ':��ލ,�����bȰ;�
=o���x�C��ט�P1F�b�,��L�5"p�q�i����~�{����߳=�u�]� ������Q^ &Ԁ����%v5��6��AIF��}P�=����q]O�2�w	;w�1AK���������
�u�c*Z��
�eL]�[1P����9������jD"^�;c0D�X	̭����S2��K=�% �Y���!!���X�
���[��Ă�
'Z�p��&�@<'<���lN?�q	���zV�Q�k����;�����I��WBimhkX�5�84V
�L�h�e(�7X]+18���W麫�D���2�: [a3�p4��ֶ�0Cp�}Eo,��T�i����*`t����z��Aj���P�Dˋ���]����o�@AK4+,�V���� �8�s��|�e!&#��������Ђ�c��]�)�����`�0��!nR�k��#̻��7iW�6;'�`��h1��M'o��b"&���J1�q�&�x�#��C�S��v��	Q�0!����m��N �}Y{x���������`�d�j��{�S��r-�	�
  �	���W�N:�|$�J*�Grue(���7�Q��!�mwtt�w��]���H^��b
eX�'����}�� �<����`���!ާ8C�e���_'�Gv��Z/�y�o�NǴg�>�5����6���֮�HBeez��F��Lw1��i؊�H~:�cO�0^*'K]��}�c�G��V�-��@�bZX  �.�kC�l��Wҧ��O�V�g�LN���Aea-׸<S8�%V$o����#�/0����N�@<��0�ˏ<<F�^�%Y&@-��v?�v�.�[�����/��𪗿2�џ��i�(`��tl?;�����>>I�d@�h�b5c��,-YL���Mp�ҵP�c�ٻ'<�9�o~�,͛�%�M	5��d���_y��^RB����VX`����w6O��x�R��:> ᳔�H��^U4_)��@Mzc�v�1`�9�i	5��!Ȥ�[�f15=����+|�_�_wC��j�|���Zc�E��E��*YA���*��Yi	 �F�QY�:�)���7[� PT-cW���lLo�Cb�j[B��u�is9W�s+<W"�H�om���h��?Z�nU�)����_bd����ҕE��C"��e"h7��l���`���i�����pH5���*6z], !2d���lڸ��/��:�֨h:�CG����[mݟiat��RQT��|Ϳ�vX��nl¹N?�t9�W�g=�Y>�/T+ �c���D�q�
�%=���lI�G��l_��2��Z�'�2G�S�3\pAx�v����`�V%���h�x�'!p��*ɀ*kc���F��[ ��X������&�>7H�0%�8x(���_����H�3 ��.1Գ����m>TҎ���Ђ�:͉����t���b���s��}�mZg�r�SGȣV m�Hzk�i���4��ԥ,5?�	`(^kb��Lꁅ։9F6�O��իW��un����G�-�D��/!�;�}8m2�$
H�n�Rs�J0�,O���/W��6�����p��m��yn\S%�!��5 K�cU�� >���%���3F���@�zC���3��Ʊ9MB�+��2�1�>�g4W�p��`AGSa���(�a�j��Jsg1��J)뎎�d~����ג� g�<�+������{FG%*���8�T:֦M%����IB(�QB�Hy��X�]{wk*S=�6+����lEE�;�}
��ޥU �M#��oL�h(#!���]k
U
5��.�0��o^����[T	�^��AkN\*S2V�����s/8o���XɯG�2������l8ĹI����L�n".R1j��|����<5���.+��E����)ۮQuA,�]E��Vm���[�p�ֱ.�)�4V*d�*ۻC�:��H,����СA�Y�D�<o����G�'����
��;��賐�t�*�-x����S�ozH��zr�i1�hbV���Si��՚0ӣ�
�+�_s�:�U�}Ƶ'�v���R�9Ҙq5��u�pL�� Q����Ub��:OȋN��"6���E$4AX���l��y]PtTI�=,�!��7^] $�&���D�_���ݫ������>��O�hLH3M�li
�[�K����5�Ѧ��	0�S�U��R�;Y�vӦMV����
���1����z�i~��x3�4!�:\�,%���Yx�LӞE���d�5Klj�J�0Ga�`o�3��{D�b��r%�+���c6&M��`0�� +U��_������"2,��*]먞�q=�&��0��ZƖp��C}`�y���Y�(�_�m��Y�К�q��B�eec� J���^d�?�>�yr}��(9n=̖K���O�ح�>�ɮ�Қ12��}��c
�֯2 ��G�,��Y��Vh�8��5���5fn�b霚�V����*%ot:���^r���M��>=۴������T���>[u��������(�7�RY ��%��p�A;I��G��5+$�өoO]O/g��<�I�O��-�,D�O�s�Y����y�G	-U\aHn��v�ko���]�SB�i�
mU�����޿׼
u��x��(��RG^�J�T��bMEi25�����-#�^�ۤ����ᡧ���-��h�?B�I^Y�&��k���0YnҸ$�n�Y����h[�畧aU���<E��}��Ʈ�ƄU+�'m4�����Ru�.��Y��?Q����W��z���z�,;\��hH���w���jO�H�� ��A`�,!s�bw 0ǩ6�!�EV�L�T9٘�9����cQ��"dyHZ���~Y���9}cì։��ԛv_��	��|((�a>�a%�u>���"t34aiuq�m��?�����m�5.������f�ׅ���*L���\�bO����,%g�q0Ry���
YS-QT�ؾ�LiLW�\m�0��{��c-��I�o��ڻ��U��a�{�=& �X��&NN1ǙF����}�{���\e6oTfԘ�s꿥���X�V?S
��m�f�[���٪�D���4�3b\�0.󝂅J+����ˎ�⾱�G�i��c8 �ՎP����5���q��Th���?xP�̈́tB\��[���re��g��e
�K�#��a��笥F������w*kmO�Q�|,%��A�Bb�=*e��Nw^���+Wo
���_+E^i�ej�ºl�R�bq�QezOR�3�a� h����>�|a1ǁC�۲l�Iw�i��;��8����,&���N�N�qn��%p�U�b{NvJ==]��ݠ0ح��jq�*ղs�W=!�Â�%+6OftA ��γ�H�/vH[����VNSG9�u��*v0�B�h�_PL�ea��D����R7�(��O�L�ڸ�T��0F�¸��`_�#$��� �B��b�ttJk�"���:�<�.��!N�D�E���p�������_ �N�<a�s C�jF1V�W�Z��hhRE�n	7�|�;2i|2y8�48��B�{���.H��&��T�>a?>��[����!,�2T���q�F�K�V��< �t
g���`Ȓ�e1�g��f[ݨ�7%˘��\�>i�p�8�z�Z��6U�����LQr@Λ�P�B-���B�dʄ��6������i���_ ,�6,iNY֘��f*�c�b/�f�o��H�ta�3�}b S� ����jx��0��@����;��c�L`��ޝ�k���ya�`�x��t,k>��x[:�g��{��)��8��y�'1��LZsd1�y��z���5UO��m��:�e����Z���	t*�ӔW�3��?��OOz��4��"��)ՠKH� ��2G�,E{8j ��p׸a�ꉍJ'h����.U����p��+�?}�?Þ�]�6�Q��C�5W�j��5�r;��S�m���w�Non���������8�Z`%�DT�ܯ�8}7eU8�yr%W�9�'�\O�N��y�����b�"�E(��'����R{�RT�����k�AZx�G������ک�8(dF��
��g�Lm)�5^PB�8���Ǳ��>&-���>,ɀ�&�8Y,��$87����� 3�]6�Z�j��Tpl`l��Ο�EJ7UU�J[�y���} =
�����k(.��|}�̈� �����&���E�y��X�턔��g		�������cP�� ���غ � �� ����.վq Xb�e�B��\EP�j礔~�����g,�*�Q��|�X��㥦�	�azd% �~��= �ZckU��1�vP�$
��O���`bj~�����yy���,���Ǆy6),g� �̠��6�H�B؀9zqYX���5�盐S�o<'�HxU�����Z��b�3)��@QbL�`"=�b�\�a�#�7@�_�M��[z��S���̰1�P����kO�a/�Y���`����ÊN+�y�� 9p^��J��3mU|��=�浘�5@,F��Zix�u��>��G��j�ڶt�B����	m߼6��٠$�Xd}��
����A7TR�Uޫ����{D)���f�K��![?j`x�KW_n��P��2�!f��ZC���x/�o�u���[�w�7u�[�_�E�XAK5-�4ĳ�,�{*vI��.,f�.��c���X���.�3�"� �`q"L�:�yȪ��:�حӡDb�d-�4,$d�R�Q��Ѥ��)�sBd�>ȓHQ�Gk>�zP �h��筁'���X�V�A3#m4|�
�����u\�.Bl�Z� Mr���!4�^����hw��Km_D��0s���pOW�
-�T�P�L
���xS��	-�� r��p��R��Pd�w��F&��6'�k�Щ�c���9y�S� �rz"qO�z��K��"�lb����.^5�����{������h;�r*�w�
X�H��I��6�\a�O  ��3e��t[�@�݋�e���-��9ՔM��;�s>~oLU �p�Ř*H]� w�"-��6��0cccAz�q�Tp��޳h_�<$�	���XQ�BČ�%�b�*L�����q��92 !��5^��⁉����U�6�y���N��r��A���4R���Щ
	�A�q���=S�A���ФƊ2�nL�kгCr�=�4��o�xX=��q|���Y�M#Ú�B�C�'�R� ^����Eǂ6vT`fh���Oh�j��w�yW8�ÛCI��i+����1S����5>!F����eZ�bX96��*�h��-��@!Xt�m�+Ú�N��W
��BlϘ����R��B���H�@AKm�^-&���a%��1?�1&<�u�t�'��5���O�cL��CN�Ķ��7�&|�+��~;GC� ғU�+�	PЩ��P��@+U1�Qqz�"�+,��\��m��?v�83����. �-b29�D���5�S�K�Q�;:v�d���4=���w�Q�Q���^�	Ǐ;Z�g7�d�=����8Zf�y,���a+@f��^,R�χ&qq�mщ���I7�[�B���>vߑ���5�oK��}��y��7��&6g1h�'c✝��yR[cȘ��Q"(�eH�2�vW[��A��:6 �r��2 �u�0WN���|���SQ���Ƌqdl�����s<����W�M�#� ޏ#U+Uc3��L������yoe)�����9Q�P����
4�ƨ�FU.�_׏��@��n��t\� �\���ay`���J`&�͚��g�y��-3&y8��f�������y�`i�Vx��@��B���)�����;��+�d��٘iz1���e���#���{������.��xm���N�ْhχ����C��F1�e
��Z�\��NZG�drX�yM(4x5g2*}\׌�[O�1s��t��LϠ�V4"�Yh�s���
�I������MX�XNGs�M4�Uv���T��Kf�û8���Z ��%�;}��E�w�I�����T�O� ?���T3��K,P>����ź�k$\v���U,5RFBa�X'�e\)��zD5.Cǭ�-x��j8K�rQ������g�x�p
�p}Ik��O�<R��6��V�>��	���4Lp)�&�[��Sh���5\�!zv�쒓	���u���H�[�5���!��!�P�a�����rᑵ欂e8 N�b61�M@E�0���Y�L�da �*���ļD��Z1,:�o�����&\j�Fکs8���;�.@�l�(�5]�捥�+�Ac�T�29O�lM`�+�;;e9�̱Gc3��D��PQiF%������-��!�gc���³�����C��9�I�	�kd�6Sk�ڹ�Lԗ�����ۋ��Ľ|��Xڈ�f�)~>/>�l��d<\b��f����>~H���y����k�L����C�'�6y�D��J�O!s�.�-I��8v�Ҕچ�4N������͕3�e`�4wKsڠP�Q�w� �|���r�����tK���y����Ѫv=1E��XN�h�fB�F�+��!<%���
ڦ!S��ie���PѬH�R����@AKn ���&d�]��F����+�K���N
(�;��'��6��zBP���m�:wo۶#�t�-V�xÆM�[h�@�e�x��T�bU�%��ߧ�"���]~�(Mr�����ڽzuaB�r��{�Nӄ�Z�y!�MKB��>_c<��zM�`��T�����Cv��A�bIx29m���les���@�ĺz�����!���[@�Wh��"����DƒQL/�e�3^<͏U'ܥ����؝];��p�~���(H�i6��k"�@Hc�ӵh�l=� �Ξ�w�{c����8�t��u��a�)����l�����K9b;��Trމ�I��H�J!90�E �Sf��ya��c�%��J�i� �F���.$9 �Gۦp�}VV@����c���?kH )|EƝe2j�꘣�-��u�35����v���{[���J,��.n{�%��n��ɧ�b�=���O�Y�� ��o� �Tr ۧ��Tj<C���N�iKڌT��P��^��.��k�ǅg��9�߳D�>}��bk27�U}zLZ�	�?Kݻ�p�Ԇ�V�U��:���
1.WH��i*t�f�<cZVu���aeRm��䩭�Ą���gp:�-��V�BU�y�A�9�T�m.��&_���"����D�o'ydX ��%�3�0sr�(i�"SJ��h`�K��/�?�����yO�yh�Ʉ�d1ѫ�����b���J�S�y��y^�M7x4�q���?���Xh�Cc�����@O#a"Տ��ۢAB8pZm�
Uid����mtM�Ky;�6D��Fw�i��8��Y�q ���R��Ս���SB���i4�3�1�U�C=��֠����r�E��:䎒�^��
����Y��2G
��9ǥ��t<��7����|�SB��?���l��{aƔ���U-��ǜ`���ԯʝ���[o.9۽���:Yh3�^�c��6��J)�t&'T�!9H}�F��k���R��f��7�l"�DN���k�9s�~��R`�z5s0��;�j)��MX+���+��9%�ם��� E�DH��D�`i#]��f�lS��������XR0�j���f��ZS[a-W(�ȵ{�x��b �����b�A����� ��Y�����0^�@�?faY�LbMB�]>�;Qǅ�l�s�9�?؁2z��8}�TLP6�c[\I] 
ࢗB�Y��b�[aOke��Q�;�6!��w�czʘ��>)��
��ԉ��6v %B�����)g#d�727gTyZE �1ZZ~c���C�e��<T��t=e}c�̳6+��(p���S������tZ)O_��~o�K2�C���?�[�,2�}\��*5kEG
}����fa{hk�O,���p� h�C&'Y��s��&IG�2���py�X��?�c=�����C| ����Z*���&Y_��[�O-p,v��Y�Z�Ȩ����^��%'�T	���
�J�3V�����Z-6jv*@DL~B�V�̜�ZX�ݠj�̠܍��:1�!����B�.1Z�}��#��4EֿK��t��� �(�6��}^u�uUB���]�s���(�������vE<d�[��<����,��)p,�c��6�)��a�Ү��;��4�d����-�1%�
���s��5@(�Ȇs��S�I(��� ����y��X�ބ�f�,6�e�X�j}�\���Ӛ::L�'C�@��V)]��v�R���!�n\-�-��A0�{���=��3�9�8I��R�?m)|.��plv�8G�[��F�Bx0܋l�9ψL�S lm��,�rR&�EG4A�"�� ~NO8��@6���w�c�%h���Ɣ��զ�N�Wm(�Z��~̇�d�
���3}����SĀ�X��LKgE%��q�Ԑ��z~�<�0�����&"1�)��Н5�as��F!!��R#x1{q�z�3�2�1y0h�>��\��q��L'��8
�y�?B`*�<�k	k׫@�>�bE{�l���kDUC��3��k�)���.��y�Jk��h>w?����z.F���Z:���I���(����
vڦ�;s��Y�m�Ȑ��S����d���'���-��VN��"KZ1��(�Wf��,�S����O��H���Y	SYgi���VT�����"b���G�EbpD��Ic�(k-�c�:蹤�#��7�	�y8�_Rc'a��XM�+^|3��_���'�����ݩe9�˴� �\���:�&��v��<%6�
�y� �D���P;O�P"$��x,����{[ T�gO�Ŵ$�w�'���!N�6�9�h�>�ut|�\x�Ha�8�E;�a7��v��e�%ǏӤT�iY(��R���qL@P�;+G&Z�nL��Ff<���bEa��ϑÇÀD�h˘#n�/��X����Y�]#u^��\��T���#����
S�{r��1��)���4.q,>���_�yĴ`�ʅP�]����=ލ������ d�bj2�(���"*O�!z�U� B ���R��'�Y<�@���S�,L��}��!x���yd��+|m�Zx`�`I9�d�{��Ajݢ�M���p���;��9�9atH�7�*Nb�z/6#TxN��-��9_�b�{�5��bC]/�ؾ\}��<���������t?Sb+��T��C��{(�X���e8��>qn[i6p����2U��V1�C\�l������"΍E��w>���_��Y �����e�ͪ����t,���9�yp�p����?���|2�JZ �����(��z[����Κ�a�������Da�� L�zB�Sa7ճa12��T�l]���q�,z���ݸ�C�[���	�n���K�Z0
�>p2�p8�"CםD��>������)��Hz���iD�]��T��}�_�������*�j�;�_Q��Z
1[ۍ�f6'��i
�Y���r�پ: �2�gi�l��h+�ꌢ��k '��A2U���ݪ��9C�VJ���Z�ZJ���h��+��a���L���c�����k��O���ggb8_bK�%�����&�/6��v)���g؆Q�?�<dU�܉�_<�bsjߛ��q�������!�2�4�&��K�^�#�<��t��	���"|�O�\�c�F�O-I\�7al��&t�:�*zz@E	�l��jz>����f�����,4g� �7��2��'}� ��=&`��R[�poF�s�{���7g� ����'�����w�*��fݪp�m*�I�#5MUx�Fb4]ua�ºzfi��6�_�?[IP?->d� &��7�gA���X`U�ft�I�K����8�悼N�f3Ǳ�=��O^�|�o.�A���=���%�V�Wu_��\ȴb#jYC8#���ÁTjW9<�k,QK�4�v�刔Y���7�q��N3�H�a-��	Q=�s\��N�+����׀ӈp�bW��s�-��M��xT����ض��S8��xB8^�e��x��B_b}��ME��oN =���H��'2L��ς.�ݴ�zD���xD�� �!mwЄ��5���U�uE|ĳ���bz?mF
Ѧ�Ҭ%FG?�g��ɝB�bk @���#��l��N1���38!�����ҽ���1��0��Rkn ������%A��	���iZ���
4 ʱZ��jDI��_Pۇ0���a찏�nG[F����r��=����Ү��j��+  ��?����~M��wc�q��b}R)��A���C��h]�<HvЖj�-����}���4������v���w�zF���+\j� ��F^�M�҂D�R�x�S�����a�$8Osݴ�Uř�+��s��	k�Ú��P�K�]*�A�U����"���B�#�/���V�숊����t~/l��^,��i��z�.�xZ!�.�����}ž����g �x*>"�� h��쏸�f��փ��nYˈ2�	p���,���{�� #�#(YX�ٱAp/�/�({�V��k���1-bc�Y��aR��D8�l�E'!U�E�Ђ�i��Y�'��y���!��qH��4 >@����c�wM�9&�ʹ�Q���bт;��@r2��)�s���S�������<�I{�:4�F[�cw�w�鞽 �����l9�@hA�4q�<? �&�Lwoc����G d 1
dM�p���b>�����U>N��(
Gdl��1�ϓ�!�ᤍH/X;�~1#$a-I;X͝ �����AC��Xd�(Ð�#.w���<~�S�u�-�yikBh� W_����D���c,noS�y���X�L؋�Q�����#a: ��#�Q26����BPr�tN�>~�]�96��i��E&A8@�����]��ەЊdp�K�|MNP���<  �QIDAT����S���;q=p`�l�ݷ��g�{S��Z��D��k�������5Aw٠67�����;���]�����D1��#BK�T���]>L��k��~����>��F�H����L��[NSe�U{�-��RbbyJL��d�M�n��o�_#C�1��z�̍R��� �`�m��-��siZy�>�ZZ�3�_Y�d���փX���z�z�ƞ*�x�-����h~��':�%��?fv��b���0��/���Xf[�%b�#r��ZڲP�*��UW�����a\�[��|��J�E	��
\�;�K�W{r�؉DPV�OM�����(�?�c!�M��0�ʛZ����٥�:)�"F�M��D� -��`��V
��n�r�B��n�������Y&�93�#f��qn�8�Z�=$��އ檌��8@��,~��B�Aڴ��C�EC6O���N.�pR�y�j����J�휓(ݮ����{I"�W�8���W�;D)�ź��rCדBmV����<����#c�J%$@�8de�/4^�NfG��@+D(օ���!��P�s3�/��� ��^�VSd�&�a�8������.��v#��R;3_���� ��B�X	;�դ/r��6H�"5C����z��qc��c@��Y�l�,ܨ�_&\�qM�l���Т���	��;��Xh\��I�gDL)Lt�
`�l��� 6!�K�.�����NaD��k�BJ'�Q��C�:�[6�s�;GÂmUEZ�J�[U�i�1E����Jr*�JK2����6@+�c��e��蔛V*f��Y �]�-�ތJA �5��4�-�;��f�/��� h�cl���ؖ��3u�rl�I�CB�N>��N{L�Ĭw����X�ww <���*��u6�=��MW�֮�V4��?��Jv}�BN���V����$6(�M��$����7c�"��!˚��ݼ3ש5lE��5Pod�p;x?WI����/ӭ\��t�R��yZͯ��Ѝ�Y5^�C�E����4�>�g����2V �{eo��,U^Z+��؀��D`����~F%@V�l�-�8�$�A�P!��Wc@t����������bl�s�{1A��D�I���8l e��H׏�S�Ϝ�ۡ���#��<ܳe��H���V���&��>ll8?����p���3�ź�� �o����Mi�;�is�怋�S�yҌ%͜u����h@���vʘm���.������3N����UșK0cn�q锬J7 V���W�e\ʜ�t���ݴ� @Ș�]��O���"�SK�nѩ��أ^	��r�~�硒򤮕����32Kc�`�V)[��n�:+_���'M��Y(��Bm��A3���=�]ʨ۰~�B�{C��1��Y����è2� ^T��Lu�l��Cp��m�0�f˞��������0tlR�~��e���2l&��kQ��1} ��e��~�ᶅ5:�X\h�3�"Uka[쌀������E��eZ~O�<��֌�k�]��ND��[��Z4O',�S�`��\�pӍ7�Zo��Z��M��,��_�bͭ��k �u�צo��#�a!�F�*Nƅ�/��9�G�<s&i��-ю�z,�ӟo�I�����,�bm�ba,�)h!��n�@��PV���G�G��)��}.�R����M"tc`��|a�iV7{x+�:\��>Q(��A?����9�� d���� |��g��r Y8����7�U��75�8�g��,�ëÜ�@pN�H�9��q�~���C6�sG0c�$�&��YB˄#5]=���H/)��q(��ҢX�F���s�R�;ƒ
�V����@�i���:D��6z��� ���(�%������K`J�o���B�rʤ�{c�q���2��`>U*%�����j�9_	[� ��'d��u���l��`�	����]����`�O�8����Ш�6�� ���`%�� [�P4��0J�4�A���*e�L{)+L(v0���?�;ƛ�^�p�\�R��!c�Rsc�����:�z��G:�5�K�B`K�U���U��9�Ը��ޙ.�D����g�a�,/�j���@v#�xذJ�����ki�`���[������!��z�o�9�@A?���`w�Gm�׌�&�|Bl�A��c�"7�'�;5E����g���g�,{V^��lQ����� �>%Z�U��ږ)�L����H� �3y�������+�x�q����F�H:~w�v��K��S}cq�6�c%P�D�8+q�nF�nD�1u! j�P��"���Uh�?K�2O�aG*��6��NL���VցM�����<�ԑu��������0P�R�q��4 �3�]��1M�<���p{-F��gX ���?s�B!�"�gS+��3���sT��Cu_�����@(}�,��NZ*����*�04��΍��׌5�t�g_"p��&dc�gؗ�U�#4
�R�NF�A�K��ZN��,]��~,�^<�tE�Km³V|1�u�����`�(������З���n�#4N ��W����٫�;K�}�<4�s��K!2�?U}��5�S�i��e�}�LG�G�B��%7�j,;K��2�����Q*�#t�Z)�Y����1��[&1r�Bu�	�Dpl�?E��--9�doH���--�{�l!כZy����h�5�9j���1�k��U�m��P��ιj�
�@kvK�y
�������CG=*��Fj|f�C����S��0�?o�\��]Z+R����y��
�p!��ò�Y�2g<��FW���ߵ8��X�n,�A��<8��J;p���?�i�ҹ�G,lw~,��������p8S��:iE��Agה�6J�N�@͡^�T�U��De��QN�8m	��cD���ءm��"��_zo��S�ARdX,d�\#�!w���P�;i������:�F�XY`�Z��t]Մ��0�U��J�<۝ǝ8H(�ZسYv��:,��$�S"��\o���Y@)
G��l�I��������� �D����v�r4VO�ГbP��;+��D �k`^�%��.�N���c̈́]J+�ؔ[��|<���Z]�U)�ɔ��F�W��zp���o)�1۪l¢.Pij�3l�g��qK���1�H`dʰ7:�d=lF�kf�k�8G����	6�V���F ��Q�)�c�(�1F1�.�0aI��0��s����H
�p��I#Ľ�,�M=�`S���k�{�\����V�-ia|m�fJ�e�����?�{hnn���g�a�V��k�w�
�mٲ%<�1���
�}��{A<�F��8�J��0T�
�ͭ(���¥ R�"g�[�3�3k����������=�ݡIM�a�����+�g�s�`X�fe���������<��P}c+RT�K	 ��C:�dr����0�"V؞)�w���Dz�h�b!V[�";m����-4~�H=��6����-q�y�� �
�}�~i��X=�P�=� ia��8��pG*&�&~�%\_���l'Td�;����v�����;)}k�D�֎҄��Fr$���[Q4�ݺ%����i����ޝ���'T���8|֜���K±,�B�J0s��#�h܀��䜽f!�&��L����.��S,��-A�'��ZX��F"�gfḭ&.�����J�~P���ǰ*��3/�6����.&:&_|u}�Dৌ�����c�#n.���85�4�J���-rL,J��W輴,��/��v�&t��0��s�J�� ��؂6
���>+2*\D��CC���U����������R�Ī>sM�i9dKڜ <Q�,/�Z�;�I�XB��^��u`0:^jN�E�jĪ�q�Cr�5zOE���?�F�b��Π�%�a#��u �E�c�ߺ�j�'���:vT��1;"aJ���(<5*��3A��	�E�?%�P�F	@�XL[�����\���s�0$1m���ha;�/�1X`�*�lP�cY4 9�� 4O���<?z\L���[���v���Թ٠4��5ջ$+�B;��q����y�*K3N�q����@�F�{(�Ƚ�*nj�^c�uo��L��7�>ۣ�����p�S���/�;���#�C�ګ4�4Z�����o�!�ض-\r�B'M�0�~M�w����9�uJ�02@�n�Nئf�"xZ.Y*R�Q��_��������p�:�i� h�#N�<m��P��;M'-�=N�
}��z��G�q�WSN)�\�9P��dd?�l����J�^�0�#M��bѮ��l�L'��%�0�^Rx�=B� ����W-5���s_X��M�������خV��"x,�r���1%��z9&���%���~k/��݂37h����k����d�2�%����;����Y ��G@�'ڒ��� o��uv�ޡ�-4�ԫ�Ƞq�@0�.&鴨�bE�\x�IE%Y1r� کN�����`'l�KYU,�w�_�(ҽ�����] �(�F�0rh���&jt);2'uOh �c�����g+ ���u��gt��'����
�zd�M��5U
}(;�>b3��k|Z����po�um
�H'ҧ��5�Q�l `RN����2hl�u�d�x���0L-�=ٳFA�R��s@)�g�q4��pưڜ��a^��d#8�!U6�5�]�au�t_�H�̙)��
]-�la$�O����y[-䞻��c��a��Uw��������z���'?��p�c��B����K���a�f47p��nR�e�YE�3����fUP�P�xxX̡�dL)��_��	`�p��0^�I�X��z�YB��[:.�@ē���e`�֐�����s",H8p\:�	�|�BJ��:�������駟�ݾ-��8da�;�C_�Æ�kB�f�����2}X}]��w��>@e1V��\�o�>�o�����ϵW��|�������U
L�]'4�6l^jUe�J��<s�
#n7l�g�]��L��, M��z�)�����E�jZ� �G*Х{�>f	c�Tܑ��e�=��j��2�$��J�z��<ОD���e�(��HѴ6X	-�'��~,���a�L�jU��r���^dMw�N��r�H���lh�ĭ�|�C�!�_�1�t��@��P	9K�Q<�
,a�/�8yI������J��{m��P�:>kqoZ��:�[�sm_�,��/�b�-�'2l"�B���Ǚ#J��0�4��=t�D���√����c`����N�3@�}�����ўj�W�^	,��P-c�X&-��9������u�Q�m!L�BY7�;t0Nz�tbӡ�{Ld��ޮ~[a�5�œq�����-Cԁ��gt(?2VSad&u|��͍��;&�0(`�N�YΎ�B��%��d'shC �����tu��n�����2�-��Am�9�k��E�10�D�=��k� a\�8xĘ����N�j��#ǻ����尽�znM���ռ���	mI����nhQ}����}�u⮬�]��(U	��֕X�6����I1���i��ח1W*�  ��hp	ȢAę�/�����1�
�ls�J�h���>r���iYx�s�kl�{�Y�8�֛o
7n�{Nأ��O;=��e/�\~E��G�Z��;wZ�Z���0��")�� v�8���	BM� �E� �ROw��%�_̫V������d@`��z�C�Τ�����ݪ(s���L��S���V{
�J`I�ؖ�����U�t�2��n�N?����jB��{��.{ԣB���Ĭ��5�h|�ll�<�5�]ڗ��v��J,йp�!��{�N�b�"�Ê���5�Ņ
��[o4�����������7�M�P�PW�mf���>)�60x4,�0�Jv"����A�P��C;c�ד��ň�'S�s�����A؄S�S�l��zی������zkk��]��3x������ h�#��S*M*� ��Y����iu&���%�%йq��v ���D��ɗy22��_�����YD�c�"�Z�{^Xl��	Q $���^��A�`ט��p��k��^/}��ڥ���=+,kn	�ݷS�d��;C�~����D�sSr�bW�\k�IV.G���L��Z�r9�Z�1X�~���r�e �����b��W�P��9��|.�Y�z9�>s�k֮7��Z��ش;n�=4�n��8d��7`#X ��=a�}������!sj�C�@ȧ_�cY�L9@�p�T�"�͐�9q� ��a��p��]a@��g�6�_Z�c�n�~[0G�3:��̇��V	l��1��\�#v�c`��/�y 8��Ͽ��O��['��P�0�{F�J���V�����z�5�87�@�m�i2����k`�L:���
g�yv8���6	��۷?|�[�2f�� \z�e� ����ڷo��{��u��E�u�)ï��˃�8&43 ��Ί�0�&h�B*| AXj�j�lܸ�X�Σ��[�V���+��~�/9a͏�;�5�Ҏ]{Cs������B<G�3(=v�[��*5��wBk���燹Ch!��̢�Ȱ@��1Y�ZU�Hk�*�J��V�Bs��H!5l��{��\tX��6Tg^�y�Q"�29��^����� (���=��_ ����>�|�֍ھ��a��ճ��uKT4��(�2@�� ɨ
�b�P&@�F6���G[v`� 3����y�7��C�l/�-���Kuyz�Q���Aa���֬g��9�!�8�£��nиU��3�5b}&�u� �1(;"����0�τ�Q+Ć�͖e�R���bk3�g6���:),��h�� ��#u@�p
�-�-�O��Y ��������0[LC��V2c�g�2�,���F��!4�Xp����%Zt���qR���Hdp���5��)|V1���rv,���\9J���b�ίX"E��#���ж����E���aSxֳ�θo��0��a��[E�2�c�9Ugm�v�0
}N���ؘ�Qe�Q����U|NU����5��iѐ���Ң8A�Ah ��:��a���叺/�^�JZ�M��ۥ]�!���0���8���[o�3hT����u��I�=(m;��?�R�W�[V����^cU�3��u�&BY�6����5�''�3^�c����ȹM[��ik-�����hԅlݺU�`Y��λM\�y�^�,�m�7�:�?��#1���u�Ղ�:.���a�!99&��`��:��
�ӡ����30���E�9.��/�R�FM��2]���r�b
zĜ��|=��~�٦aa�V�6���q\��o�յ6��쐍���}y����cp�IK�ҥ9#�)���½;w�~̯<�Ҿ|�J�>j�A���jc.N:���K�3"�@И5k�.�䒰R��w�����ͷ�e�C؊�9}��v�Ç��l8"�퐀?��"�7����4i�	� 8�ň�ٻ���u�C �F�|Ps��$��n�!��U�����8?JB�5���2�����k�9#pq��C^�\���f.��� �s&02�k���{47~`s�Ea��v�Rg{��}����ٽ�F�ݶ����ф6#e:*w���ԆP�*PI&Yq��p�4Kuu56���L������������G�.t��A���^��&ˤ�?z�Ϙ*6FS#�@/�(����FZ�1���'���8E<K��@��e��$Y��?�5��@��2 �s�̀���\[!TA:A%-�/�O��Y ���O�$���x�2 īA$��,�Ǟ+�L�{ �A�ty@�����SՄ��(��<�k$�C�����������a�������#̕�%D���
����s�Ia]�3�
���6�[�m�j��B�h��Ύ��a	/�8�|���w�1��i��V	����TG�A���F
���D�����g�BA�%²F��19�m�w	���t��"�g�c�(
�>��n��l\���{��9�s�1��o�a,Y5Mqo8�;�u�0A����z��N1D�4�4Ї �H��3�OG1i�t�>���ڑ�����L����ζ�σC dCV=Ԁ�"dw����+׆}���b_Tf��MM]b[z
&íw�c �]��C���B��u�&�(��<hE�(m`)̀ ����lظ>��b��ᬷ)�r�C"��&}8�s����[íw�m��y�i{�ۨ�� �ǝw�i"�U�V���k�B�\cY��Y�ؐ�U�4xͯ��~	x<��QX�0��m>�.�ǥ�u�B�A@�5n�޺�l2�*4� �U�/0dwI�1+pU*���ez�jX ��
����O�~Ŋ�V��@P���a��<x$А��@IG:�E9,V�R�ϙ�n������@bߪ�h��YGŚm�h����%��t��F�%CxL�=(�TS�dL��X���ν��L;�߫����_~�1W��֖Ч�61[Gu�!�X�
���	�ػ���l����(�٭���"��Ex>>�g� �s�گ9ߠ�₋.6�pT��:t��z�}Nj������w&
��1a��ZK�W�Lcݦk]�r�i���s�%��O{��E��r=V���t=�ދ�d�9(�/�S�ke���qڛ�C���bz>�����g[F� ]��{����m-}4��a�Ma'�*-V�-����I.Y<^%�S� E^����bZ�H;���̨��x������V��m}��@�_,�߆��Ц��C,���n��a[\"#�W
�!���_��S�v�=֭�S�PU8��_��R�C9��fD�:3kW]� ]AAuP��̕I��'��,��_-�1��#=á��6l�zn�+�6kml3&e��_��QNF�Q��
?�Z��gF����k�n��.���yv�?��bg�sA�f�s-[*rƥ{�����5�KWQ�p�2|�����D�še��PT�kv9�X�r��1E�3���x�s�㘚B���93eSv�(�s�5�u�ݲ{}x�3�v���OX�v�-�b0��/7�A9��.=˜���L���=���G�K��&��.4}Ǩ�.�,�|Ӎ�5(F�Q�	��u�~݆aL�q�ڵ�
�QШV��Z�P+�F*:E��G=�W��;w)ԣB�
��
v�(<'`�qD r� L��@�L��a�ˠ��bպ�apX��耴-8Sl�?�6 �]����Q1OL��v�ut� �c�f\�k����<e�Be����n^�ѓ	5��� �BF�&P�60��uP�I����U �` �O]͍5������^�98[��Q�z� �v���-l�X�0c����I%psXO�4a\FuM+��5�$� �y*�{׬Xv�Mk�Wi��),x���|-����L��W k����;u�}�b�N]�]�kÖ�N���
3�ܹ�jք\6vR����#�[���\��ZM}u8��L=_�K���!o�!+o�vO,a?ƈ�@2��4��7������y�gP�X����!@���<�ﴍ��F�}��Ko$پ�n��J�-�b��D
�`�K��kB=�� ,JI/�h%#��I^V��e���K�r +����d���8�)��}�c���'�,�`I�_�;�o���]�����+yew�p�V���QQ:' �Bg�X��m@y�@-h� ���p��,a�JEY%VA�= ��uon�!Auv5��e�c1wv��١�ѭ �4*ؘ(�Q��!R�zՑ+q���`h���dVYE	�s�Y���{vW�*iք��7�>�{��fEi�?Zl�J&�܎�k��A�g۽���:���g>M���QN���hPԊM�v��Yao��>���8�so�P��mA�
��
�ᘆ到(�>�����l���"�`��g(y�e�͢l.�A�Y��u�a9�uo��4 �bd*��i�V�S�ʕX��jh��0l,Y|5�0d�Q�yR�Z�Oc��VI܋��n�<B�)[jla��b����@��4�,��u떛&�۶��]�1
�+�k8�a�3c����'A�M�V[+��D�u
gM�v�"m���3o�%�\	a�a4  ��M
Z#X�*� ����PK]�rik�J������_�����-��F �MN��
����55օF����RGH��&���1=�d����)�W�{���y����~�u\@��B�C6?4����Z�	�<����_�П��q@SE��!"̝6�l-�O�.:$ا�Ė�j�o�5�"�Ս��X��p��T]��TM�~M8����ߨ�넴V�z� ����
w���֊+�aE6mۨgz��=��	1˹Wjİ5�铮��4Rht�+��Ƭ�9��iY�|�m�����1��`�i���׹�z��x�6=�6�d�pֱZ��B$�� � +0�l�֋%f^�����j��+�k��vG ��}�����a͖���B禬'^��.׭�Q9MI/DԴ��4W5��U�]�	��L��I����V7K`��Y� �~�F���P6^9��/~�K���U�]���#����	Z�`d�"F�=[�Q6[U���Y�e}��%�r�d�L(�_B�&z,Q�M��Y�I�R�7��Ϙ!��S�b��ۙ���К/|8R�Z�9�q])�U�V!?-^V�_ ����'P�0EA�W;Qj� �����/~�j���(^s���a��i��5�R�N���Z�6¨2���T6,�*�/P�����Ĺ���A�\X?��	�
��M�eF��E�[A����'Mx@@�ki�&��7��bB���ł���Y�&IN}hd�v�V�F�#�u�N!��=��� Ŧ���9Sf��i��ک�>��m,��N�����ڲ����fA׆���9���M�Ӱs�{B��ې B�B;��\v����Dͯ��\d�a�&|���R�� ��WJ��ܱs���+6OʹZ�\�p�"��ׯ�)��p�㺗f�j�n��|V3V�����j��3Ч�V������8&V�g�^����9G�i���Ҁ/��>���{����Wz�54	 H�D���z�ă�֛^}Ku�J���Y<�y�@U]���E5�v��T� SY�`��E�i��J����A��Z� �B���̍m��;�B4M��U��e�j$.�}�����Z�V��~���O���kW��O���x8c�&�Ȇ4Lϵa�ڰR�M�"I��l�� @v\u���Vi,���*�u��5�F����ᱣ�h���=LE���	�h�M� �oVL�%)��Р�?�x����ՑB�s�������=�b�
��y��5�X� Ԛ�����5qwu�t]u5��S���TRA󦦱Ul�6{:�u��T�\�ta��k\�Ț!8Z�^�[�ƒ6(6{����36����\G���v��g��b]�q��Ϣ�%z�_܏e�Ա�s:��z���m�JՔs�|;;�Y>zo��^�a�2MU��r�*��#bK j.(�`x`�i�tw'�g��m�i��%�yq0������L ��e�-
ͱ�.���'TPS�@��Ӡ&�,6u���� �2�B�iRvI��r����!k�X����T�`�hn�U�jG� �Q�'ۤ�M�9Mٝwt�#�#��������'Ѥ��*�!�`P\P�*��8�0 @C�1.`ĊWi�g��,�3T��i��eUZ�u]�1$hDN����V)[H�#2C�D�k;V�� 'ÂM�L�0c�uV��6��s�y٭j�//w@�n�ś���Ε�5Nm%��+�}�{��#�Y���}��^��A?Á����� ����j�j^��ҁu�|P���ѪR"$�g �؄�<$���!2�f4wתHz�={�+�"p'�F��Uh���>���Z<���Zjl���,�0���u$LN�0!��i�FK�E�����H1�U���mPsKU�Ѯ()�Z�!~	XA/�m��C(���
0�ku���0q�	�Jr֑�P܏������|�:�w#b�
z�*cm�.	�3�P�!�^�{wޫ�bT���ׯh����_x�����������}��� 힎I�v��J6ќB�~@�a�&��ö<3#��+Վ���k{��(i�������W���N�  ��DZx � ��!�J�����2�؅�/�jk�Ko��󁭻��t���ʧ<%􉄜��l��xJ�~�JH�V\Y/�'�10�}�2Ϭ_���}������l]@��y5���.�&Ⱦ��q���{^R������]K�=Q{�T��?�c���8T����p��r{ ��?n�o��HhG�+�G�F�w����e�e�=S�\��xI����u��U�
�&XXܭ"6��SoV\[dy��'��%- �0'�����E��Iٶɏ_)�P:ESE����QΛz �R�Z#4J�s"7V,UV�uV�Nj����p��<Te��tl+D'�A�oJ����w�)���r����"�%*�{Wv���� ��XT�kgQ$���d��O���f�P"5�k�{9?NG�Z?���a���#�(ݚ��L$��O�]2�`%��AR��G��<f�J��q@׀�H�`�
 lX�I�B'oB�f���tK3����%���~Z�f��)O�n鼰H�^� p`��(���I�nh�-�u�����wT�r8 �L;�J��?������Ph��<){&+�d��#�
�ɆU�,Ҽ�s���b�	˫T�y38.G���b��R>��%��'���4�G�*��3�e�c��T#�����C�!�N��R�	�CS����z(1D���h4j�_�'=S��l�0��4�$n�@�+�5m�='�5���jn� 1o�^����qB��i\'Z<&��I1����m>' W�y �̧?-�ᖻC�j����u�ݖ��K]�k���c�N��j���� �ֽ���?�� ��j�6#T'W�����zF��}�z�/��n��blm��m��
mP�H���p��������~�-��}��![�ɥ�O1G>;55jʣ�r_W���bw4����Ш�$���!��K�XW�֮ߪ5CϦ�%
��>Q��8�M<�܄	%�LJ;	#&��ǵ����JI�C4�lMæ��Xu��R��V�	�]��֎n�.!��-u�@���	;�
�J�"��bI���^�OG��90>2�qΦU?ش��v���%R`rQI��R�0Y�{���M_��ܾYq�6Ux.�]����/��ɟ�"�e��"b�����Y8��[t��P�E%ڝs�T1�!ЊH����P�X+I���Cr�X\��lrH�q��!���ӄ�X�tl2�X��#��1�yL�"��U�J���Y��W�mi�qܞE�NSM� Nfwk��C�2/�F2��- h����G�HX
�E�Q�d;J9D�t�~��$���B�7YNUrB47-*��,�b��NDǮQ=�)�!�v��$~ެ̰�sq�>MM����N r�.�$A�Ϝ*@�XE�ESQ����K��
�9��z�{�w�)�:W��
z��.���µ���v`�I�19	 ֐�8��u�J9E�T��"�;TPAGR���<+��������0����7���z1d��l�սh�Z�B$��'��1):�J�Ep��
͐�gnIcf�`�d�i
jR�ܗ��F�P=lR2�q.�~C����8�3ij�=�����E�悾����� ,�����o0�:���<��݉,l ˓��ނ��M`�*Y뺭O��kա*d�
9�����n���w@�Ds	�Zk�}˄�g�_��5��CK��0��G�cD gR�B�#z_sKUhY�Y��B��W��ZB&�F�&��V��a/���J�̭cS��J	��xm� u<o,+hgh�f�|�ќAW�f�N�ذ^�v�6DX�&��q*��MU�*��-4��ڍ�	(���g,uz(�)FsF��t1����=�7�7�Ċ��k�l{h����2�jb�YI7��_�K���f�M~�탘�T�׼� h�>��s-q��H-1��Es�,�z��mV@�j�XW(U��ÃS?loj���s�n���>��o\�姉�������ǿ���m;�ٴ|͕e5Z��L �E�(y��iaqA�@t.�RMML���"@Z���vr�_�>;s-,4�{f�0Y���J-rr���ɍ[�i-A���-H�2����)�c�v��+~�K�y�`q�9�ݡ�l�53���f��U�f��Dt^Bl�׊8j�c���9���*cD�$�K�[(H�RݏhM�A=kH��^��҉t��#twxի^^������S��E����ƵXO�!6����ƨScV�=:�.:��g�u��0+S�0�����{��������D�K���Kd�XA(�p���Ӻ� b����e`K��Å���t�ւ6
hr�o�ճ��U��9�Њ�6+,R-�S �Ze�ؘV�8%�K'R�g��)Cԫ��ӷl
�}�U��k�PTqL!۱���w��бgWh_}��-6T�G�ޥ�K�X*����@۴'_�,\��a佧ަ���85i@h�`U��(Qv��h�&���7�ڛ������;?�jOBr���E�;����M�F�C{�RQ_el�lEI�j~r݄�d<J
4J�Bo��PDhXl�ب��lP���$��K�Q�����5�=�Lْ#W*oO����y�y�H��F���	�qғ�8���u��H�
0ʔ#���S�1���NN�R��Q!WD�*�sT	
Uu*� ����I�I�C������3I ��}C��������F'�͖
C*D��m8�|�R؂��f3�Q��PU�jE�oC�u�ze�q٫B���m%�U�1)�6miVv���e S=�T����"K��	�I$nl����MIC{4'������HF�%�V	 �ia��Ȅ���c ��S��:i�3�"mh}��#�-q���U�(���`B=�fT�g�E��x`����sc�u�c/��Ӯ|��_=����>�s=岭���c������W��cfr��u-�[��F�@� � vs �a����@��M��M�^DΆ;;����yfi�����C�����)ձ�-�d�@����xUW��3����(�L���0��݇�!4��ò\�?v�4�� ��1���$f�EP�2\�8�Tk��(t�29*~��w�$�	NNN^[?�`���X(��P�A�����B�����w�����Rײ��*Ԗi���n��J��,0l�n�*o�H�M��p�%熿����xs<�����W�/}ɳ�{�����w�9F�/z��Z]�j�()U8B砇�Ha�RR���5�]��%͇X�:	b�vT��������+X���H���K� �H���{��<�R�ݴ����r�aHN��da`% Δ셃�ƦgT��3������g^&��nQ�ot*�/_��+��e��-���b�z��;L�������e�H�=@�FNw��`-�A��8�R�$(�ac��$�U+���k�B�:=+�1+A�c�?=<����L+ž��o�j��� a@���q��Yh6:кh��&�JJE*��{ի҆�zN�Ū���U��V�a�Rl9��%b�F��Ј�B�z1A%
oRJ ���M�YԼ������.����A��x�l%�����%�O}��#�_�R4z�~i��`6��o��+M���i�
�XSY' 0��-S ߦ����-�P.�1�9�f�@O�0jU��,�8e{�T��\- 3(���Bx�����J������|���ZD=bY9����!�]�9��ӞeD�s
��
4�c�
E[�ѓO��4�c�=U3S���JU̚J���3�:F���pkQESc���PD�?=�\���l&YGK�U�R6�I�4�+Y~=r,�A���+�*�BHG����;�ƪ
�3e#�{�?���=�?~�O����<�����/�����>���V��u����qcqiy�АsJ�@(�"�>�yr�qk]�&���܃|P�v(eCXj�I̯'�y�#�9�BVR���N�[�$��ΒF	0d9f,���̑�?޵�K�������[~�Μv'���C v����5c�p,�
�}���6\G�"E�S�e��]��ء��w�#���O�ݥ�|�$_��ځOJ�FOW��� �i�(t�0��s�>K������3���
&�ʲ�	}��xCx��n��a�V}�j��U��M4l �Ke�v�
5��t�eM�+�k|M���u�BG3�N��&��rD
��\5u-v�8hvχ:K�T���ׇo]��p�_�u��n�fk�4%�4G(��x!Ҧn�2�LY�d �}��_�w�T ת�������7�ax�K^������v�Cb����e��)ۨI���Q#6�D�nlb0tv�W�N8C�)1#ԁjV`���!����0�K�/XIfϘ޻R)��׭Rqʃ�����^���W?W"p�ilJ��T�`ɍf��w��$"G�"�3�kc�
շY	b�W0!��ݡ]"�J��L���1?}mh����J��B �q�́tib����Ⱶ7�Vb{䔩��Nh�[!e���J6+誘�0qbfaa���my8,�${�H�^��/���H�ޞ"1.</��-�T�[��9���`=�R�S�Y��=b?�:P,ۗY�:K���ժk׈)�D,=��,�^� ��3�%J�� <�P�-7�d�A����V�}g�*�K@��U��:ZH[�3�?������#���^1�%#��h�l}���!���`�Mճ"F{��۵W{;�n�����<}Ǻ�+ƚ�jg
�`j�thd��Б�u��x륷o������Zժk��Îl�h����tI%V���W���_dd���#��A�&�G�@���Ukg��Xul�o�+�� @K=<�{�+~�����'�����ӷ�{A�J��i>�ř�rP�-�ژU�<���@�B��5[}g��8@��~9SC/�Ң�o�Zp�ny�ߊ�R|ֲ�&��6��9�nN������S<�Bv[��On� =���뷮�1��Q��l,�� �5&@h�� ��rml�7���S{���p��������K_������:>p4��e/��_���Kj���#ݾM��cd���n}T�I�X�(�N�bAtlٻC�f�s���tw�{�zo���}��t"�{�S���,5�����M�W�P�ޘ�12�{�(�?�q�j��L��.9�^9��pM���k���5��}t��{0|���+ܽ�#,_����;���y�+�o>�2}>�׮T�Φ����-pTר�r�%���O�BS�:wk�,�I@c�t�e��F�~�����o}�{��/YX�^[����s^x�ܧ����`'%����d���#*�)=�e�����Fɡ�Aŉ�.k7�v�U���K�^�r�j�	� ,i\���õ?�>l<�B�v�?��Ԧ���<�4�yv��*2��wy[m�����z1����{Ͻ�н��j[�\�Ju�UȞK1��6�}�c�)H�ݩv���K$EQ��|\�d�K-�FFƄ\��&�� Lw�ҟ������ĳ�۰ hD�ٳC+p3��	�W� e�)L*�/@SZ�vb&���bCS�1%oH�!BD��Ӂ�#A�-.�(��Q���E[�9�?�i@��2z�}?��@{C��6���Ѓ�6ǀ���y(a!HA�bk��ƈs�����Ԩi�*�R���\��ª�ƙ�#���ɡk���K>w��gw\v�9��j��W�x����7�������O߹wە�U�6����3M"IK6��^���hc���=�Uy�A������*rTZB`RMcU��*�`��o<�O8��%{��^�����������γ���G&��I��CFTK�ɢ9Xd-ƄOLc�e���2?L0��ϩ����=h �H��j-�P�T�M7�EU��E d`v�H����r�A�[=��x��p �� ���4u�jت�b�l
�pa�қ����
+�|��v�j�g�Q��y������^�!�\�.�;��r寊��	��?K�'o�hz�D�[Z7BNBK��������S.]�/�5M�>��)�Q���}�#����=?<�I��=đ�E1�hj��o5rd�x���o<���;W�(�q��_�!\����Z�p��ݱ-\pچ��J�^�7��p��#�S�F+��څ��g5G�f�^���A���w�X[x�h)LDd��l��غ�#���Ĝ�fmKh^��å}��d	a�F�O�{��Úֲ��n	o矉u��9�{�bx���+��u_h���)W�⎳r�����Ӟ���<Ӵ&�r2���uN�K�s��yW(]%݇2�i!����רΕ����CaŦ5�}o}ChR�>�@���p������a�u�	�^���7�!�s������GՒcm�R] �^�ꗨ��y�O��Ca�ڻ��٤4n�kjL� 9!_!@sF�����`�I �}h�56�,%c,)��K0�*(��ΨH`��ܻ�Sn��s5�T�.��W�iVɊ�4}b+��dJ�A2���Ђ�����ssT*�E�-�+A��K�ä���d�lލ ͮ���vRT���2�f2���:JC�ź⏰}��<�������t^��h=�ةJBj���P�6�?�v|a������v~�U/~�?�����`���u�����#���S�zǵ7������W��h�|�-@+�r�K�Jg���DN�>����B[ ���qs��b��)Lq�*��F���wΖ=�[�p��PNy�i�&?���^�����_Zװ^���5�N�e�K�-H,Ld���n9�](,p�U��C��ve�ŀ�;`�'<B�2(~���"�P�|�˜��`9v��G>��9��O1c�5���O�\�:͋,�.[4�BH�L:1i��'禦�hg��R8��&��Ii3�شY᫆�Û�rL�r�ii�� "�ٰ�4���fhZ;��=�B���%DĈ�gX�R9���_?��bk�@�-�0+A���m��a�G�Z�,�v������?+���M��кБ^a�����ó�����B��~��jG��w^>���T�G�f��?��й�@����
e5�z4��*�������+_	{o�!|���~���7��]a�ڍ��mM�PhQ zv��E�VC$_, �c,�V��B�����g�|�\}G����n�>��+_��/ޯ��2��,���3����?{G�O��^���
{��1`R&�̊u��WVK]cآjҽ݃�O�����fU��6/��������uo�sc�fH>��&��pX�U03T�T���H��W���rI���g�^�����w�W���I�t(��Ya8��"]oB]2:���V6oj�X�j��@����Ⱦ�&Ҥ�Y�M���#q��-�䖨@v�\�	���l��704h�J4?a��q	ݩ9T$FnRmHJ�a7;�J�G�
<jnQ��Q�7��A����S�1m�B�ZS��u�QE�z�}U)HE	��u��!�R�B���e �A�?�@#��A5%��U��R�r+H�͖aR�Չ�!����r�K� ��ځ�/��/��<���m������877!�^}���s��}۾��?�����W��P�M�{��+��u���_�F��z�LmE啥��zq>�\�j��@�h�z�:)�Y0��e���8��R1�.�׈�i�3G7l�r륗�G���z�c/���?��������u��P�ش:�4�r��Ce�^���T�5jk�CK��(؊d�%"4����x�hPh�rJ�؉l��C��y�9L��(������8�]������d1��Rp�5�MƋ�[�U)@��QW'7�jv(ح�e҆)������r2�^���4_xv���1|�s_
��5-mZ����~�V���C�Eg����Ec@�Hv�@�R�9��d;��ü�j�N��fF���i�bYښ�;��D@��h/.U��ȑ��O^��v5�<+\{��f�"��Ғ�>��S�WJ[���I�&&��k��?5%��]�+��T)YBmX�a�|V06�H��ck��a+|é5*xX"',�	�'����c.`����]�#1C�}��-E!�߽K镵���RS�4O��ϐ�'V�t�Y/�K��"8��S���@'�R���v�]�t15n����v����F8c��p� ]�J�ֈ��߹��T���������7���sT�5�?��7Æ5��%/}Q8����WL���px�!��t?ý�]W�.���S4@pB C�X) 6Ť�+�f��5]��U �u���,$jb�N��`d{�����������������	-��հB-?��j_x�c��s~��7��$گ��y�L?��o�Z�4�:������e�O��X����Wÿ}�;��M��J��:�ڀ8Q���ރ0�<Idt����:) co+H����R���=�&�R���x|�a���!CO�C�V�-ٚa��jp;7>|d�}7��ן�/K@i)Y�Z7u�w������~���i�RQg���峉cSS\4��ʰ����z�X ��%�Xq1ץ�5�%T_�ҎQm��W�Yu`Yk��{ʏ�7U�}�_���o���TQV(�)�<��11���G1�^��91��a�J/4z���!=X?ö�H{u^���([�f���\�cD7�H_����lV��W���#s��}�b��!}OE��(ѝ�BI ��_֗�����FJ-� �5,��Mq���}�I�AS�d@!���u�y�I��Y�Il����%�zZq��n�M� ��S�� ��E��0�.�Nm8��aSb�p*M �V��febV�D�pX;2��VP�D_��T��	���� �`Ũ�\����e:����B���H�oQ-�Q�
��+h+ֲ��M�X9s��,lC�i;�h��; �c��E�d"L��I2�>_5a�}/1.x29D��*�?e�����~�]n��Z���?��M1�%��mo���4f��*�z�����Z�P�դ��
�'i�z�=���}���&�J�2��N�uP��uj�Ю�k�u�Pxޯ>9����V�RƔ�A��3�S��x��qr:vk��m�d��jt=:K�M��@�D�d�Uڒ@���(��H�6�g"+B˦����)�<)��WTo����/{�uJKT�l����ܾM�������Nx��_�'K�Q��^��g��3GGC������hoy�o�']~a8���孍�O�������*,[���Ԍi�'toT����jn[Ɯ�uϱ��^�\�MKD;���<E�����+UpN�:�ȴ�_�Y����P��H-;�$P��Ա}����e�7^��������	�4��l;�w���|}wg�	�וh@�z\戴iM��ދ��tCsC��ʯG�2Z�PKkR�Ƿ0�o&� M��TZ<�m~Nu��5#���t�LU5.� <Q��=�-:D|��ҮN�4&����,	��D�������UY��.O
9���M5"��Z[$��ϧ�M)�FF������a�i�3�@|Y��ź�������:/���*1?v��~c��-&�,���c��Bנ�'�)�R�n\Up�
�Y��@yJ��
iy�%P%��J�E�[Wj2ߨ�LM�&�AT�nN��*9��/�<������β�.P���~�$�8{U���������:E��:z�'\t�i��xr���?�.���]7�RCQe")ck@,@��#껥�Sa��}aBmZOo
=�#�y��VZsuX�j�	iv(<�b�����!�0ƢT�kt����͊�������0pxO�~O�j��+p�c�3�x}��KU"�����sW]$2�&n���oSH�����o�|�+_����1��*e�U��BgBJ�D�N��
��ѥ��-ר�K��\�
~LvV=�9k�Fh�E��9፯xv(��K_�O�lԉ��5�ۤ{W����zj���=�r ���<)��T%cx9��N`uN�ŀ�u�91�cbR���y���۸Vۙ 0�*�N�P��(ܥ��9)���~�������d�}��Xs�"<�O�G;��V�ii g��p-/RE,U��e����j�Eg�_��p�~'���.�������/}~��u�B�X��7u���a��A�c�&�ia��,���,]�&���5��� ^܊��w�	qK�}Z�i�&�زT�Hr��@0h5U�Q�9~��_���Z��33~��Yk�>��������ǏN��Ըk�@aXm&um�V.?��+.:��Z�i��e���8�J#(U�E�]ԸjXXk	=�!��]��c�V�]�lY���љr�j��C���8$j
Y�eb���0:z�0�ؙ��E���%�U#g�y�f��v�Ľ�j�PbV
u��3�@
k��=�x��2Y6��f��˳P]�t�����ؖi���b}RA'_�-��E��m^��b *-OKS2��p\N����XTH�J���P�Be�P`pF5Z&�f�Ճ���s�*9�������.����W�vز�p��'�[�.\q�����P+��yn��I�R-�9��Ë^��p�Ĺ4�,x��g>��Y!���J��]L�\/����u�>d!��=����+����S�|�z2u�.v�j�9L���fi�:�W������<=��տ�ᣟEu�T�*�}9��B�2sEL��g��۴L�������F�Gì�R[����/�M��� �&����Z��OSGt�G�~�O�nTO29ezDU�v�W׹=��c��5k��K?�9O�T}��U��oڨ"��l:<�O]~I��ݲߐ�q�T� Z"�u֨��a�lQ;	F���U���O����7�Is}<��^����	�x�3��V�Ԥu��c�X;'�w�Yᆛn4�UӠZ:�}TF�Buu���I�D��i���U#���c�i��<&;6r8[�,��hH8���j��>$�3�;���/c������"����(|�k���P֊����@�\
�JCF����>��de:mE�Q���d��^ce�V-%�@f>Br�� ����db		��7�m��&�|N��"��֍91S0@V�ܞcv;�A�n]dU�았c��2sMdYJI֖�p���G/:s�w�ҋ=���c.;��w~���޽��%�EEm4��� ��fKssg}]Aij��H�@AKq��:�׆ʦ�*k�gkj�TA��/�^__=��ֺ�P�a:V9|���+�zm��� ��r_��:�	J��I;i����fd^Y�j��H��qzIb�x2��-zY8 ���\L�1L��"ĂZX/�q��9i,���߳xG�X� ��¥6L��3Rd��RS�0D�e�z�����/�~�^1
5U�{���a���hWh@�jU�E���\EMK�~������-��ȩ�y�
��1_�}�=�{w�{�_�W�.�<<�����G���uk%�}ax���rd�O������?�����������i��i���֨�29���%�	�� �t�}��36�7���w�o�0!�J�ݏ)3��r��ן�k�z�w�R��kTQ m�M�cs���������~�	Լ��oox�)%ۦz���o}�����Mi��¯��s����*�o\6m����o}o���[�*�*}���5/��ҹ%hWqD�ղ�5����#��'�#v+�uŪ��'>�I9e��+<R#v�4R��G�7���p�B<o{���.:;4()�C���}%|�_ ��(��������+@��p�c.�"��fX�b�U�P=�Ç�����û�����������f��w�&Ӕ£z����JV�#Z}�F����ׁC���j�F�11B	�������R��Gm�:�K�\����|�����ד��87\#���g_iMc�}����];Á��l�B�z�+��c����k�K+�*��z���$Q���дl��Fa1<�^�o�.zؘ�獴���@&(��F�'W�¨ .�iJ���H&��f���6��6��
���%�?�v�*��ѳ�I�qb|lv���г��巜���a%������?{Ƕ=�zj
�mi�g~b|�\eH�ͯG�2Z���ӍfbJ[.�?* 6Ewg�?�/d-ZY��4='�ش�m��T��vw�ۍq�А�aZh�u�R��X @I� Z�s�vr���s����i�`vX�-x�ύY%�>�=\P��q��t<�Sd��n�ɝ6?�5�=c%~o���YϺ�B�rk�x���FAԺ�d��@CtM��M�x��_��K8[���(�Bw��51���v�h�CGyRn�!T������{{�����B*^XQg���9	W5�^r�.�,|��__���TO�'�/[.�"��z�5��f�@�ֳΑ�����7��@E�ո����O�2��/��Cuk���g�-|���}�ƥFm�����װҬ��()����f��C�?a��K���/;��� �؃��1�
+��j��榛n�ÁЮ����ub+����w�{��^ۤ�}(|�[����&ց�-b�zU�X B�c۶{�U�4�z�/�N[;������תN�5WY��J�`j��À����WT{K��	��v�����ưf��[K�^�a��Χ;l�z���(V���e�[n�5����^��ɑ�*��ad�/���1<U֟y^��W��z��ޫ_.{Dz9Mx�<����QG�X��	w�)�TL�OM�A��A[�A�Rޟ�7�ĳ+?�,,�9�~����\�r;�3��_$|�o	�y�;�Y�~t���[��Q6؜�	��7����>�#ij���G�}����\����*��y_�k������� �Z�*����Z*�@;ڕ��xf�g}�.R���H� �����Ș/��� �_�|��A�H��^�O�o���Os�z�����g�����i텖����usϷ����#`�($������=(�7�i� h�#^_Y6�P]=֧�j�4����?;6��C4�B��K`�|dx����a�����j�5��,K �̞��)���Śth-T�}�Α�d8�q�\�`� cb`}e�(�u<��[w�R�?�;��$/ X�^��7�C�p�m�*��Oz��X?C�nBl�?�]-�ֳ��S�J�+`��&g	E�-��fw��h�-�L�/-9*��D�U��$Ǒ�_���:
v�����W8�P۴v���[׋��Bp#�1O��TEW�;]Yd�]3����&�+U��5�\�i�P��ມu���u��LZ�~U��g>Y����W]���:.��:��]�*�)LԤ�mZ��� ���kC��c�����H h(	4 �%�2��q�{��Δ���c��l��F���.�ތ���OA6Y�v��:��ڿ?��O>��9�P�@�r����YL�@�!������8�f;e�0-ب�Ya��Ȝ�T��C�����}Bb�~b���J�g+ugH@\������9��Q�#TӤ��B{:�*��CJ��;��3'�9!���	4�gk�ig���������m�jR�����������ܘ�}��5�	���i.��>�*Ǥ��0��I��'�M����\`K��z�)�b"h�2.�U�bm����b�fҥ�{���~�b{���5�ݰ�ĭ�Y��|�[
�Մ���{�%gn�����}�>e�	$��	�o:csht�
�\mz
'��5F3��ఴ@�J��Hi�8BN�a�_�!a_�"��6ր��=v|��+�'B�V�Й^��jc3�(V�.Ku�`KƫѵL�ό�jm�XV���"Pnjh����?:��hlvV�
���R"�o��U�w���89�#�j��/�2Z��{�����]�����OL��JX"fw��>�ǎuu������*�7B��19��ʡ��f%r��j��,
���*U�&������B��y����|�Co���K���Vq���L�$�0k�
�-�u݇W��wa2�����r��?^�� �|wy@�tG4t�b�u\�����3�SU��2`9:w�����Mz9��)P����b9�֊P�{FbVB��Q��ڵk����b��u�	��Q����я	�VA�M�k�-�	��7�7ܭ�����7�R�z5-j�9-�M�&^���_�e�!Ԫ���Aiu����0�~i?2)@7��u�)lԶA�a��l=���2S��{z-�R�h���S�mB�U�]��B= ���IP�]&��q���A�]��E��� p�a�:����B741%ӬG"�Ze�+���5b��S�eU�VH7T+�U�̪�e�Y�������F]v�槴�5T�h�
�]r�a��X�\v��Om����@Wݭ���-��ebT�x 
�~d(��e�~�A�"x0?��Ig���-m��B�5�},��W����!�z���[nW�_}x�^~빏����^��pݏo��f�AuuJ�Ƶ�ĭ��Wx�߿6|�K熧]����k���G��_c����pDU�ר��<������0����0���b�0C44�`:�ɂ���d���'2�_f�4�b���9�$���ª�MP�G���*+����Rgmъb�j-��*��..���d�b=Uך�����q���;���?_� h��1�4������̩u3�h��f�;g�O�`�4��%����������-k�X�)pg�yZ_�p��5|R�Ҥ���#���"���3I��=�~��,�'���v1�J:��?�Z#'��������I/�O6�e�&�FJ;M��=��`�F0�X"w�)��	 �杄	[_D�����|X��!��<�rR���c�G ��bu(�V.&�pwo���l}��tPՋ��qf觞���5ᴆ�IZ�T���%�ՙ���������Ђq,�c?,��m��L���c
����*^8"�  @��ƃ"��_,!D�Ǜʌ�9�^����ɏ�����r��-�s��A��cM�����l�J/�I�\Lsa���9$D:&@j"~9�r�O?�YӤ���@)IP&��/a���u���7�.���ŧ�'���4/�J� [��L���8�#��dr�r0 ��T�����b�?�"�m���T'�m���Z���+Tʡ)|熛��2�KNZ���*���r����½;�)��U�\�	��R��w���6�����m�����Vv�&1�0Q ��U��s��	6&����#,)��n�$�oP~�!�O��7��jZW�=�m�NC�R=�|�aD�Ҳ͔V��A����!�z:�yŒ=�*BMq
5%��in(����B���,�A�M=>;W������kZ�������C��8;3�y��ܾ�ˊz�x�>��xO���O�v�UujJ���!&����`!'[,^Ls&hx������S�=M�T��ɿ[����N�����µ�x�RRi�V'I�9+�e�͌=�E��3��F
���Gl1�p' ��8������c�135M�LYO�	�=hƨ�;*q0L�+�[[�=9Us&if�>�H4TXq����F)�sb>*q,mT�8%�M㚀��Z��ċ"r�`�y'�{aX�JoCe컶�-�3�j�
� tt߈��F+��a_B�T}!�����k&gJ���՘7ԥ����Ұ�`}�K_R��!�[e��{���+V�2�5OX�"L��]*�^��XE]~J΍끅�0�gO�J���{kT'��#��^�����C���7@�N�k��Z�cǔq'mz)��FCECU���Y�~���4mj���e�m��}Ki�-a�g ��;Ø�$���y����6��������-�F����Z���wu��I[5��,7
r��o�jV۫4���	���H�5�����Zs��\�7_��,n�E��L��m�aЫ�F@�Q��x��lC����y�٠c=}�Uu%��UE���T�@��U�$�O?��p,����� h��FNB��Ւ)��sF���]yþ�g_�o����羽�TJʟ�u�ۗ����D�Ji��/�~�ŗ�g��O����S/8E���I;���D�H{عO���N~�I���JN�����{9ձy�-�ѩP��0z}c�B�\�'����Y5�S\{Z��w�Ƨ��O,-�M�9�� Jhd(#�D� �D�-䆎I�!����U6�K�ȸu�:oڪ�̣c�ڦT�FO��Ƌ]:@�m �z-�e)����z���CZ��/��ԣf
p�3�c�G�"����f/@�gU��
/�*n�h7�K��JúH��c�Qա�\Sbp VU
CK�V�l2����8��a�� 3�E�sF�� ��S�j��_St��(5���EF�!��Zi�Д���j�s\�ڦ~��견�e�9�"��T�Iu��yƔv^By�$BX��c���kv�p�A��O'3�ㄝե~�y��b�1�_�6T�,7 ��$z��n�i���l�O�~e�U�5�Q�a�ƇB�ŲM����^���	��1/��Q��^,��� o����7|s�QN_O~��F����c�R�Ê&�����ޡ1��{y���utb��S_�޲���ͭ�i
�������U��|����t�0?X$�������+2��j�Wh1�~Ȅ�9���xު��g�d���_qW����v���y��5]���+˦�"쾽����%�"��؍��8EQ������ ����-��z��!�Ŕ�)��@wF�A��94�{KXQ�;�d��|�4���D��X�v�iG뇏 r��Oz2[�:��5.�����c�|o�MD-��-���� �S�@A��I~�u+.@Ct:%%ʞ�f\�WZhKT�b��nl����6�6��BK�r2���8�H8B>˸9rD=�v�:1M�UDGp�b�h��`�UPś{�5,d�����(�g�ki.�P��:T��>[� F*���%P�U�RU����(@���g(�c���|�ۤ�V1���C�C-,X���je��@H{%��q����' կ^Z��ej)�>�ܰY��2���J�6*D�^�T�A���r+�i�<[��T��
f$@m!��ܙ�J�����d�J(iA����տO_G����&��2�(���B5�J5��B��b���T��A��zp���ҿHMdQeD�ٰʘhr���fƟ֕A�+�ܘS�������σE���_Z7��
@�,��3YI )�*�ٹ�ؿ-��F����i�w��G�O�+������+!N�-�A�k���#�-q��r��xV��5<�����X�W�����?�_}��A�AK~]s��o�뾗�T�n*��.�⏓4-�8��R[N6�"Rж�Y2�RKo���=��uq+�T15>\̈$�b��Fqg7��pqX+��	h��%��x�@N;2��]C{X��E�� ����ig`�b�0�\�#7*��J�5?.,̮�Y|��}\/� �[rZ�C>�צ�p�t�^���ߌC*^�
F�B����� X!�kTA�2�H��:pM�ƪ9[m}�R�@�tw2�`pRaJ�pd���Q1t�g�3Tn����tn/iOĖ�M|�Z�H��s<�u�b�J�6��� ��8~��p<g�$p����i��븴1@�C1D�
� )�<o��V�a6�}E��;��V���YZ�G��5.Qp��r�J��r0zV�*+�3)��E�_'���
A���F5���J��lJ����?��Q+e�����r���!��l1^�emK��2��:�J-0��>�k�R6yo�C��R�q��&�gzt����W�a����xhs6!�rZ�gT�V$}��q��B�\.�Jy3����\HC�:�3mVb�.=���� �������E������JuU�3ݧ��$�[(�*��M����+����S��Cݶm��C=��O��t+9�X� uX���Ɇ�ꮆB�Úв�?���$��⟓�������DeY�$�4��b5�bv��-a��3��9�������7���]�e�ڻ�\s�ͯ8�?�����eԤAӀob���!ʴ�܂C?yN;�ű�����Ď?��ݹz���!Z6�}�69�t]���y����
5,_�w�:pց�V�-�
]��\Ӕ �|Hm�v]j��;֟�}���Y�'Υ���]k��|8H�
��~v0�},�g��y��hg���iG@9���M�wB�pjF��ӵ���~;yמ �b����n�B�;��tTa�RlK-�*�8�EH�ȗ�V,@B��¿x�Ƅ�V�/�e�8;'GSQ�����2�o�H:�)\F�M�=��<�7����n-,�{F[�Yo0�:!Qv���>I�!0X�z��dz5��U�M�I�Ka.�Dr�֞B܁k͘��;���a,QdM�AHs|�\3���X,,�Wu�|-�.S;�+f2Y�7����;e�%�MFk�ߌ��|�ar=_��B�+��T�̘=Ӎ�c,��`���){�o���F�0h鹧����ʶ�zN۹������=������{�145�Ue�L�%@�Ҩ�ǌ���������r��zY k��8حu���E3ݣE��M3څV�V��בɀJ��[ղa�����򚳮��ES]�����_���_��\�����K��x��׮PCL�+��gFxh~��>1y�b��>'�P'�5�o���'̲(�~���Y[f����CA'����̼��y^W��b���{4��k�`,�1U�D� �	 �uk��t��g!�>]�O��"0IvJ��9���^i�.FE�LG���X̒�p*骑Up~�0��'�K�!ZoDw�?�N��M/�e�gEd ��S[l�yh׶p��lҌY�Z��b�B�@��V#��j�n[;増�� :���.lLX}'}���(7�V�3���^�Z3{1�gi���EGz�v�@� ô�ƗIS5)V�O�g���x!'��<��&�h�QUSzLN�z�Emw��	�`��h�Q��a�k�u�����J����y�9�����|�,}:eFZF �$��6�`1���,;^6>���2��g(6�5���1d-<sșw\[�>��X՟��q��8�L��æ�ã�&�/.)k��~��;���3�n�rP~�ׁљ��~��'޳�೫�V��S�ƼBe�T@�ácG�7/�o�M�3\z����2Z������X��G���ytY��9��,�J�],]�K�J�^|���g�5U���������M��SG�u�����54�M55��ssǏw�t�l���笽{�?������w�l@vgM���H���h/,;)��Ӓ{�4go��W�����ŋvJ�~(L�bg��XŬ���s<�hXp�񓛵�t��Y��9�3ӑD���ȼ������o�-Td�X����T,E�8N��� �A�t�'j~ _�1�/c�����7{*�Y��Tw�.���5���޿�� Qr�&D��*�}�0^z�J��UV���5c�5�k�� �]+���X'�������?k M�VvarıכP��Ҳ����R�{
eΉ���9����P ���P��k?Q~�F���ʂ�E��ήcV!��vu�`y�4:z��A/Ay0N{�c���I{����%���Wl� �;$�n�FJ��r�%���TBB�SXbY�X��DB:�$����}~ߞO�aΙ3sf�+E�D.����^U���b�h0j�E�K}�H�dW~��Dz)� V��&�W�i�%W���D	X�����8�j'����n5Or���W��em=�l��#HD�����`��Z§�)cs����L4Ϳ�>�33zݝ�F�z�?z��^q��'��YX9��~�<�+���g��+����g-�7�?n5�յj���ZV�z���&4n	(e�.�/f46�P���;������:Z+�`�O��}���5j�a��͍���8��c�,)����=����yj��2Z�6�٫��	�S,�I��N#�`���?�Cc�k޷���c
��%5�?�)#Qy6�y%��1��ʼ��+�]�|hE���s��07r̀�v:��v�Z��Y�~M�{c�X����Q%�}��T��o�$rrs�L#"�<B�49Y[Sa�[a�J{�̾��tܖ?j�B�����v��w�4WLb���-B�ؠ��Z���8[B��7�+�W)y�O♇vE�?=x��u�SQ���wLS�����ڥ|��kK��C25���1��V�x�}$�>>��&�Y��� ���>%�t�䩪�����Bz���W?/�.U7c5�y�ꁶ����^*�Ӱ ��'�R��8%�ت`D�A4�c���jQ W)�l6V���O�=|J3mbH��J������n��}U<>����y�W��)����6�2ʃ'���K�d�'��y��y�iH��-�J�e�^K���DK���[��v����m�mAJ�jb�\����Wb�_*z�8/�/:#�C��J�>f����e��"Ҿ��4LKy��?��i���I���l�9!�q��u/�g�}����x�7�I&����w�KKjƟɴ�A��_�Ǒd?-B��BT�W�0�b�s���\=S���2dh��"�?c�ޓ���w�Ŋ�u�7k��1>�+�=�0�w�x)�g~`��Ӊ^3h@ ��#�­C(ͭN����E����p@�V�҂/�����d%�|x���Qՠ;�M��V���ff���1Nǆϐ	��L��mEѮ�}�#����s2�񿞲���X8����h�"*l��UcݽN�T~���ZwدS�柤H+���4<�4ܶ%xG�V�ݙ�9k���>�0ҙ�\���B�pS8?��3Vh��*�G&,iL���C��!��Ɉªҙ�|H���K���t�74���*�b�{2��$�&��e����[ǳ�1G�8ô9�� ϔ0F���]9��q"l��ʍ�mZ��ԥ�ta��C��3��1r����*T�Ÿ�T��3��ۮW�q�Ue��J*@�L��u@a���?�?�/�rj���y����i{>�/ڮ���q~_۠�'b칀|�-��:��v��-&��ۂ�-�'��R�4U�u�U�Y�݈�SАbI2m.��)~B3~��̰v��f~���0}��in3l��C8^�Ig����j ��
���`���7x�d��&NHdR9p��C}J'<U��4�_�O�ŴO�)����"���y�4j�P���3B="�;^�����Z}��-�г���t9�j*�@6P5$�lkrx ��e0ԡe�v0���.ݶ.��8}�&�>�k(�~u�03�=��h����e>w�����_�������L�>�8�q������k�F�G�]je/w�u���W��:����]�S�>�:�;��՝L�^\�m��'�"��E��c��Ɋ�D����UH�h���k��FGKw����$8w0޷� K��n�f���wR�*����!���M�\��o��Y�+y�=C���}����l<g�F�p2"�k )s(���ɠ'��?G����I6��O�7��*֠�3�bo����rJm����@kr ��M�-���9����jW�`��āT����.�d��UD ���Ф*�_�uW���9�3����ΒP����4�%���/7Љ���Zܤ.��C�Wk�[����TC|˥���:�6�њc�͍]����u#\c�$,��ت_�ϸ��r�����;���*������ ���cs�U�[Y1%oO1�4�� U�5n�6΄A ���Q�^�f����;U4)�y݁�\@#c�B�8�z$�H���:F6BX����#3]�/�m�A����Z{�M~j¥�|g7�߼�qqfC`[N6��}]�f_��}�$��g�\Q��n�T�d	9����&�����6z�b�V�_l���fJ���E	��ӑ9d����l���M�s�;�|���9���MY;4�-]Uo|��t���@���<��ĭr�op-�_4���1����-�ű1P
�5 ��(�\�j�W�n�>��������ۅ�eJ���2�����[cg�_��
�L^n?<�xY���� ���{�ۍb�k .�>MZ�����\:]��z:�X�%�B~fwX�
:\6���M~���m��H�������suC2j!�����`������vf�6��+��b�ū�=%J�ˑ�2DDR�����|5�㸐^Y|x��VܟL���~�&/�ˋi�����@� گ�{����K�
Vh��bDG��Ƥ�<�H��%G<*:i�Ax�0L�K��̊��_����x59�������N�?1�Z��1�$��M���{�P�x���E����RGJ��;����*{�M��lh,�ᙅA����`��)����c���1lD9q�'�+1F)�Lou$|Ø�	(s�N.�_���,�v������oh�MPT_�W
C� �oUǭ�k�Jڤ翵�ɾ�ƫ!���F��G���Dsهsc��J��Ĭ�F�!֫�L��?��Xvw�z��d�$2J�s�#4�Mc�˸g���H1�����=U��|���Ϩ�g��g��]f��=����5�!�f�FD��"M��&��_�������)�E��%��G�RO^���7p}ǽ���*���w�A���\ķr��G�Z�u�<kz3@�TjS�<�K��}�Zj��v��^�2H�Y�"٪hg��n�|�&I��^�OF������$dd���,S(q�W�f0�f����Ӗ���U����9�6Iw4vW>`�c*J�f_�g��{&��t_���]z��q���|����/��Fv�٘�r�v��9�ڄ��S8��-����y�*VV�+��f�6ᕮ��M�l��	JB�t,|Et,��Lu���$�&�}-�r��M��6 P=�G�ԏ��X]��^U��	��c�+�C!P�r��Zs�ċ!��̫ -�9�}��-�m�[�PT:cM�z��UnV%��Vs�j\$06��V�M��}��Ķ%��!�5������<
��K	�c7t������������̤�ͫ(����''�T� _P����\Ca��Y�,N�*jU�L4{��Du�Yw�'����|y�o;�`�?�,,��_ʌ�RHWb�',���֢g��=����2������34���p��'�s����F��²�'>y�ա��f�7���,.��B�����0�]�zM@��It�w�iM�u�l2ι۹����WM{H�S��Ÿɹ"��[0-׊7;}�9*|q
��y����	�|����ͤ,41��P~��z���il_�њ?u�Q���ף�9��5׼' �%p1�\��`t�����%�W���D����H���Vs#���2����dJ]���޸j{6�Y֟�ӱ�38�N�J�,�$���٩5���q5�������5 9d�I�Z~A}�m�<7v^=&���F�f-���(kMuS�O��>�yW�Eb�i��ix��W��kL�*�$`�x�ko����V��㴑����l�J�"
�X�����9B�����{o��;���b�m0��s16���+5[K��r��]�0�Y�/h,����I�q�H��-[5l_iQ;C5�����2��o/�_	`>�'o;e���|k KX����[KiB%�/���V^qX>O@.W���A~"�x� �k�4"]����N�$\������Y���<;f���^)�vh?�OΙ�0�((�O����&���*�H�=��Nw�}F�_��%���İJ�,��шw۬|3���g.�/g`9(��&&���sB��OK�q��G�k�U$A�-����ь��X�Ix�V=�cNq!���� /���gt���E0���]Ll�k���AO �R&'MyvG�Y��������ӅnR:97�o:�\�+7J�d����.���������%ϩ���sf�ԗ/��Ņ]����>I%N5z;�p��g�^#�"����dl4�C�2���[]6?Ȑ�/M"��;���!����ǉ�']hK-&@��d�V�Zt��x_K\��lΊ�%��'��m���o���8�K%��<���]���O΃��O�ϯa:�Dr����О�� ��3.�u��R��}j���	t
��^�gSD���||����c�Pi ��-E������MDF������)#Щ��'��e�ֻ3E�K�o{~� 敜TU��]�?����&<��1��g����NW%<g5��.4J��rx eX��pB̮�cl,{2j�}�6��q�b�'��n�a��� �Hc��� ��"y��>I�(�=4,i����>�>��;�&^��B�I�]����IKt �:B-�b�Q�F�@�\�Nm^�3�2�v�\��ⲵ�r�bY��L���"Ĉbc��1���a�0�J�iP��[��Y52q��
"	~��F�1fNk��v~lI�)Vc���^�~G�����3�*ԝ���&B��3���O��}��-�����"W���Ե��Sxc�d�X��X?J�my[������L���@,�_�V����QZ�Ca�n<�EM�A���1�p�k�f��� {�h*/uٲ-���v�����Y�㷫�	���ʟ������J)�s(�v1��1�8��}G�7�cs<ǎW���u4����9CC��ᓷFji��$�i	D^T�o�mx�}��٦7�-���99#�ΤN��z5�Y�D����4�E~�F�獓S������۩�#F
��.��;v�:ԓW=H7��Yç�Z���|�l���4�l�a;2���m3��tcɗ 5��I��HHE(S���eγY���Z����ji��RV�m�ZezY\��k$� �];�#z-����!!%���_���<��g4=U���<���E����;�D+F-~[��t4��u�b�0\��amַ̀���tS�2TJ�U�uehٵ�(�Kj�J'g�vlQ�}]��U�#��x��N��d,��G>�y̡(��㰞p ��4���!�2��AA������(kp2��	���ک�е�
�X��F�6Ū�_"M�
�91!�h�)�Q�hb��ph��6 !!~�Go�i��p�/�@����>�A�n�=�u:�8��pK�0W�4�n�K����q`e	wW�;��?ET�c���q���6��a,d�.CZq�/tX� ��ϼ�%J������O�Kͷ��/�Wx] j��,�MUjB���ZtV� �SLo o��11�P����fO�D6���h�i�3�b��I'	f'f���ct���������R�������N��6/O\\<nI<q����&�Xh%G�グ��z7ҁYyS<���hbcE�jû�[)i�ގ�+tusc��4	

j�+�GP��@x��a��|��eֆ)Х[oS�k~��;0j?�T�c��iy�u����xe;{��j?Z���B�-='�ɟ�!󷓯�\��ke�
er�������:յ�ňm���p� �0���i�#ڱ6��6qO�����(�X�5���C{	�n��)V���A+�Wɛ6��!D�)�u)��Y�E��/�	҉)�������a2������V�Id���5zvV:�c�.��ݵ���@��27����XK�&$m���_��/�Z�����?����[����,sN�ti�J%�OSUO�^���� PK   #aX1ӈ~�� 7� /   images/ee71944e-6ad0-4091-985d-ee04a3ffb0a4.png<�eTM�5<���$���%@��ep� ����www2�&_������Uݧ�^�T��{wU���<&  �TT�� ���T���F�����@�$�	 @P����1����̸������yu����^0:��&O�N!&�^����1�I�7�dH�1�
�O�X8��r|��{ZV��a2E
%�op�.�N.݅O/�����[�c���X�|O8q����.�y�y�GS����,rP�s	0�8��������� ���0�B@�� ��Q �!��s�������mx��of\^��9��'@���@	��g�F~�{@�����v��-��A���v�/ ��߀W!����E���AY���.�-�,TN}M���Kw[��>B� (���׷ S�o��|-,蕒�m�d��"��H0"�J�P�:M�O�-��*8I-��_���1"��v��w�#K��۝�?>�`������	���W�E�=���)�Z�*1C�����{Ax�n ��$!��@D e��ی�
�j��ݝ=�ЂZ��ښ6R_ي�n��F��ƽec�G�ƹ*Rn�R���S��M�;	Rb���2���`�IZ(���IR�IS��ס=̨@��Z-1VB�A�9>E�W.ս�n�+�e���\;fŹ �ٚK�jwV{M_���ʢ�ы�����yKG�b~��w�j��އGG�yG�o��9;f��fk��ot���9?F_b�Z�4��G��\�s�̅�Q���҅��9���0���[Om�`%��!����I��ZL�VL]���4�yJ�~����>���t%��Gj{�h��6@��������=��@j�\ �#��F1)���o�5��{�w;fչ�#ߵ�#'���l?kGK�z㚚������8y��\��՚%�OS�v��t�?�⤅���__����*�8o��	d���7uvNԟwn���@	&�_�N�ZD3�NdH��S�Kv}MU��rJ��廈��U�ȓ��-��|FsI���� n�*uX DP��p��@� õ5'4~#�1��B�k#�rFmFT v\�m�򻥳;���L��*�v�^�B�:]V��P��f��j%�U
jj;�{�
��~�i���W{пj�y�5�#���i��;���$p�0�N�6��"WX�u��Y|X�\�X����U�X�v]�܂ x���QL�bp9>Yf�!�ߗ�p�Y��s 4@�~��F�Y&8�R�l�4'E�#w�u�Q���^����Rج��,���)���S���zƮUIP�J`�X{A��RS�a�Y��n9��b��agR۟Q�f�:%��ET�8�?lx���P �:�06�"�zaR�[Z�|=�X�N�-�45-�u��o��t�TO�ډ��Xs`���f�geMs����S�:*%O0��k���V�f�����"�}6�;���N㊼K]K���/I�����l���N_P���X��l}��Y�Q��'o�Z��	bGj�����#/�ӕKf�;%~�^8ό9���"2���i���� ;w����W�?��N�''O���&`A�n�-+Э���0��L
�&������<�`����e�<��D��p�������7������Ǟv%��]p���)�����@�0C-(ze�TbŹD��2ݿj�ASَ����9�ǗM����n�v F����Ф�Y��ܨ)�=�,����k�1�~r�w�kX�U���D�{�[�b�X�d[�Z৐�`��dp�]?�:ͅN4�D���F�"`�\���= ;;}H��?{̛���;���Y�s��I-!�Ж#��8+����i��B��(��`D���"*Xޖ�\���S���u�a�i��{J=���<{�F���_�����c9Ha[_ �!�+��4<<����4��E�xFc~�{�l��V��%�&�|��_�a#�#�К���\�g��G�fZ�T�s��g�z��w����R���OqO斳������͘�����/�������ѱ��vN]0��{�p�wz���	��$�K�__[s3ssϒm���5��y�O"���-~Osw���]k��_S�;rϏ��`o���9G�	�2X�^�Yܧ��[��ԩj=頡� ���`U8N�A�-�����o�E\ɜ��u'�j�]! NJ���E�=d�EKq��h\�-�#��^a���`��9���>`yoF�᎐�2���0�c��o��;�C0H��*�&[�K�\��7h���K��IIY����c���a�'��#|c���GM4���s��p��AIi.�_�%���%�����n��p�l��eI�7zP�U�'A�1���)��Լ�[k�=���$H�9�_�^����}�<ë���>�k�nx�\p�~�gcG%�!�sj���lFiԍ�YQ3�_��Q?����E3� jV�Ӑ�'e�W��CP���8��P��z��TPi�`Kg�ppeW&�i��d�~�t����(�j:8F�#7
"�k�߲�(�:b��C��O������N��x	7bȃa�������ˌ|���ǡ
�uE����2|qqvS ��l�sv������ln�Z{�:�ݵc,�>ۍ	��-�AQ�Ds��B�V��ͮ���o�m$V��L�v��	q8
�	���m�����B�ʳ�"�(�T@�J���8�[ނ��#8'o�"��ˢ�(q5"F~�dMXE*c�X��nu���]��Cq{zR���L�rz7HALh��@mV�o�&�uy%$���y����0�
,6�g��g��\��=�l�c]wd/nff�rb�"�z��:e�U?��������#��[��62�?:�"�����C��������db�����Ő��S�a�@:/�,\C>Z��׏5'���E��<R�<;�Uk���Y���>�]3��@x���u�^��L8N�ob�C���S�n9Z�)�����m�ۤ��C�  Ғt+"T��x:�#2�4��w��A2�Vn$.R W�&�e����) �����b4aA�WYrrW.2 ;{���3]�v%����;��	/A J(4��I5���#gs��K��ӯ��!.1X���&_ۧ��v����n ��q���x���d����n�Ζ��-k�?uP���gH�n�CiH�'�*�qZl���B�	��7��㋇5+�N�����=a$8`di��P �$��i"͔\�U .��b�<>>���W�~�K�D�g��^���eڛ�8�T�He�e���K�����ЋbR{��C�*6v!|�v�����TK*M�\�;Pz �.�Y���ď�l�r�tO���;5;M9 !�B�*�#�LћYYAvf;�#����/Ek�����������#�]/���L�ϛN�Z\ƫ\�ŧ������z�y5:ls].L����Ĥu�D^�&�,�6\������s���F�{/��3����k�큼�����'Q�ܑGo ��C冦�'��4K�t(�C�ic�	� %�$���w��0�"!�}HGA�h'+�7�̽M�@���#r��Їn�xq.J �����wE�}����4D�
@4�u��G�x��� ��@v��%2l�5���xbd$�e���t��Ѧ���9�!��R��x�uѻ���H��^�t6��t̣�MbK�.JUr�D	E�����4�ڴ�ۃl
?ݻ�&�nma!F����Ȋł�JY��1�[�
�U���tz|��3�D=���}�	/A�A~��RT#\bC|J��P`ӽD�����b��9nʮ�����K��S����)��hʏ�C0����ו�F�S�S 6P�b&�k�ty�TU ����Q��|�Kζ6)]�u��p.��NLJ纜���a��t���-���!����Uo3�M��Q�_�]�N���]�M�l�|<|VWW�3�/e;x����<a���Љ'��e�t�������$ �'7�SI�X��5Pu>\%+R�ݑF�Y��Gj[�x@K�)��1=���� �0t(�VF��m)��Z�����:4`݇�_j��d_Y�P�xfU&�f<�E.�f��[�C���n�;�OA�(Y��e1��L.fCS��~j��x��f��׳���
���Hh|d���Wl������$���Q:��_Ǒ)&Ք��S�G�#��7��n7a{������[�G�K�t<�V6�X/	�L^^8�-v�(eO���)�~Źe@��v'U��9�F[����ӧ) r�4�Zc	�*�g"�r9�ڮ��_��S�+Ϝ�m М�|\�"@��4@��[g��U��Ʒ�!\�kq���mOQ��"�4Jc0tUc��R�{���@9�(�Y�0	*{�y*	�)}�&-�������g��r��C9�ז�{�+Q��P2I �8�HŰYFV �jS(����Y������!211+�IU��۪�[0������]gE5�V�t�Ť������>�)O�߫��6�p��?���tP;��Y�����M�KU�4|G�+}�IJ�P61�'(O�gF���bٮRR���Qgx�N�#�adq�6��ã"PZ�o��������!BF��2)�{�܋F-�h�>�:X�A�")�B�����N���	��c�1S$C0��9����N�I��>�����1?�n�\c٢���#�B�;����� �sM��[&0ʑ�Jd�4`�d�0!y��X4�]�$9���ҩ$���$�B� j�j��>���vuw'��4\F���L��N�K�����ӣ6�P��O�L|��^�8:�:�[�,�z��c)���*�
�ι��Pd���O�IQm��[[YM8:;�4�8�G ��Kd���  ����y(R��u��L��c~��h�&�i�<�?�?�<�^��R�?��jo�ć����=_�n��[G����m�Jc@���_�4^#��:��;|�N��n�4�5E#r��ێc>�P�,;��k@�'^�s�O{����NZZ�'�A�V��+�U+߫�pU�4
GX���(䬧�T�]����QxW.�f�-�:L�U;�
�N�K��/@�(��D��9GAǓd=7�.ϖj����~�N��;<x�u�a�J:I���aS��o������L�Q665:�N�]��(t�"Md�Ϫ�Ġ�Z �G�m�Fw|r�i�H^粟
�mT���ܮ,2}ٺx4q��)ߴ�J�����u���UGa��^h|��h"���l��Lf��D{�u��^�ɸ*elvUU�'��~��V,PTo0웹R_^�Fq1V��r�����V �z�Ǒ�G��EuKp�d�D�\	�.��Y����˜W�aK�S��i�;�x\��CF�SM�B{�gEo+�_��ì�g�n\S���π�m��vޛ:�vD�h*���'�!���/x��%�\TO�]�^..��M���J]�5"s�|��s����^c?�(�:-�d�B8s� �G̃&��*�ʯw�H�LE܀m���A�+JPD�I6�4,�Cn���Z[ �Y�d+�3񬚢��$߽�٧�ϧF̅ӣ�O@���u��j�(f�w��ڧ�*`[��K�z�NS��;D��`��:���=�������|�fSD��Gj&��~�Mj���ɔ�-��Y����n�"<�M�{#5��SP/S+R*���kZ'H������L����|;"|=2�~�~	�����z��?} :��$������̆��% ����(/���,�Q]��_�=�����.��a9qNs�|碕Z��&�Jۦz��.�e���G�l7��_��g,�E�����j��d�.�r��>)����˅�+��O��.��
 ���v�*�I��R��6��M%1�z����.?�]�t�����7��[������72��!	9�/�h[��0o�����O�˜��������u�oT�'�䰡���$�Tv|%X���ΰli8c}s�d7bӤ{�(aﱳ���������M���A�0ub�-n�&" P�낽���ޠh���b^B�����?~�"�l���^�74~]��ll�$�e��L.Ɨ��z͐�5ZL�ULö�����Y��X_���d;�>�[�uZ'3l�`5ܶQa�.=p̟������;�	�Ԙ��e�!�e�0�.��e�W>���]5�lqCGZ��m�r���SN��Ð�GI�C��i�3RKN��B�H�+��F��*������hxj��.��<[�d�51-��&��3VVHN�1G�����b��ζ��Y��3ZJ�K�}o��[����%���o5��Ku�򿯻_.�爹6���7�c�T%/K��Y���,Ñȯm���rh�7WW�;T*m$6)�.�i�I�QĂ��1pP���To3*�*�L�O>�LZ��*�T��C	�l؁���,ms�6��	1�h>�i[��W��n|�[{���.rb�3nKG<ׂ�eW����{&5}�{�#�/�Ѫ�&�@�&�W�]C��ta�(X�9]_u� ����~"FU��ke��I�� ���4���p@�^^����N-�ԟ��DC�)��Bo���*ݱ&��������n��)�\!7�3��a��9�������K�~�hK���	6><<�a�(Ӹ"�Z��n\����K�����݄�=�۳�/}���u��{�^�b�8���\&g��FG½�YR#�uSS���'[�Ӑ�̿�Oл��
o�ޒ��:�n��AEA�R�53�8`;[$yHd_tw	���3�|d!Aк	��g�J�v�=�?Z�����	��`mJ���0����v�0�O�j��؆%�CSs�	��O���g�''333���c��w���v�����	"]�ٛj%�-��7R��Oj����IK �U�0Yw�M��|���g��9���B�N����ii�X�MH.�H־�+U�N�u ��fUk�[�o�E,�;U_�8���ܑ�ӽ��+���!>���_�0Ӂx���(�cn�i���7���5���S�@��7�GW�X�"���`�P<�^��M��]�d�	���ďj�MAsQ�!:��Z1H�py`�H�ɜ�gĿ�5=`B�6��'d�*+��,�ZXt��/I���X1�2���WE�0��J!�\�3.UV�Z;0��-�?rMM��V2K�n���$=JY`7;���]�E��!�0)J|�w15����s����F�O�)�t�V�`x���h����jT:n�z�2�d����0ĹD�D%ʘI�r���0�,��u�e�����$������b��`IzU��F8���H�?���T�b��/V���Z�m|�R�d�%뾶�����}b5��v�5\C��gKH�0%����s��E��dt)z3�8ǜh'�fC��"�Yi��C	B�;�d=��e��-��7�Ͼo����G����{nR������6]�p��.��k	w�[����z���SW�(%��c�>l�J{U��;�O��"_��N��9� .�o�<��Bq$�����]VD��2�u?8/�=|AP��q�����xH�.�2�tҊ���[
����]���;�{�u\�ȫ���RV\v��Bn��@7f ��9J[9�hB4����TdIyT�Ϲ�v�n��2����	��������v�u��)�"���W"�&S��w��1�䦈�ZԘ���X<{D0>�}�;"�D)r�U�5H6S"��i咈�|r�XEg�m��.��?<���
�{&�K���Oٓ����7�0�����W�do�����.~���l�bۆ���8�������v���!H버<��rYCH�>��t�ǥ}������2wk�O�TǊ	Ybq���@�i�w�	^��rl8�@��D
[nd�"Fg�YqhÜM�ߟ�^�beѶz|%A9�i:�a��C>H#e����A��{�G3��F+r��'dY��.d�'+GmMd���y}c%������A�Cqp<�Qgf휄�Z��Xw>�kc�^ ����������c��.Ę��R��93:����)��[o���������(�KG����S\�zB�KO݊KZ����=�Q��V���.����|d�D2�uyK�︍��Ԙu��7�=�:�������/����?�q��p?��#�Bz����Q�.��2SSuaAӋ?�쫩��9��qq�V�� F+�e}$ظqhP�%��G�쉆��!0��(*���h^_�*q4-�A���x�H��@��T�e�ɔ��ѱ�|-��w�NqM[vԽAb�%���e ( �6���壷*b,��^B�uA�r��6�M��>�|"�V�����'3�����OA�{ �7u@�`�*�N��#�;e���\HaEP!�)�}KxL���y�=�x{�|8�H��da�'0��9m�����O��w6})ٺ~���W;��° �ŕ���>���j�r]�L\�����[�&�Z%�'��D����}���{p 
�h;��+��a+�[��|u��4Xi�\?�*����C ,t�͊�������e��O�@��<��O�A��ivѾ����d����v�=���Z��^]c��쎀�!�{���"���L'Lce���/.X:�-%mͶ)�r�'� ġ�bҕB��I=Sl�\�T��_M��r��v*^�_�A��*���"4�j��N�*��͆��ZEJ����+aC��s�[��?�\��AD&�z�$���YOO���r���p�T��������f��UN��O��y>��y���c��A钻Q�Wh��_������m������׼��\�-����&��ͤ�eZSgmt4V�{�,fOջ  6�����O1���k�`��k������c�<����c�ޮ��#_G�F��S�qS+_jv���̀�n�����g-������R����9�عc5�sC��?�]� �F��Ǝ2�
��y���y��>����I�|\��n���67.?�񇂟�zd�{*OM:���oߋ�]��up(]cS��.3�'z�n��xA���]��A���{��~@�Y*c�1e��u� ����{C	�+m�NI�r�n%{�9��_��������[�]n��[A�C5�W=���� Ob�tb�ENcѮ?^����C��N������zvv�.
U�޷�_Z�
��6���9�k؁��V��h��g�f������%��7a��>�������륱�m6j����~Bš�xj�B�jE�R\3p�doa�>=D���,�J���5�;ɩ	�"�f1;���s$��f��55烅��������[�"�g�C��f!�����)��g���q��
��Ѓ��v�11i�����ȱD\���r���|}:�&��|�M	d�eV���wvH4"C+�´ѥ�Ow��$^��$$l577[ ]�kk���=�ҡ�ʿoǵd�SDR�a[��s��S��ZδL����'J��}�:]8�N�6�ϻ��n��r��Z'3�1p��;�l��?��U�[�3L���(�0��K�!�\��/n�
��$�s�-7;���arQ�@i�`n��(V&ҋxk�f�&d����7��s˄�W�h���&���K�1_1+� �%!�yy\GPI�L�P���t�7�M��U�}��U/�j�N�$�+$"[b������{U��!���g(宅������"9;��黢7�N*���M5=�&�gJ��#I^��/���B��"h�E��oVq쬄|�|�d���65�M
��o䩑��}���O�kk�vAA���/�\�=��+�W�˰K���k�Eس���q�=��ȣ1I�Ã�=KE��	6Z� f��5�w�q5vͺ�4�|�U��ǹo�A���d������r�1:��*����N*�I�+�L�e��)n$Q-ah���+�!@��eDKA^����*4C��S��]*i _c/�n�U��Nk/ ���� I�4|�՜����""p�&����8_YJ��a�Pnb���B��ɩ؃ⵉ�V�\�V0�<f����t�:��Q܂>>�$���P5r���A�:q�5Ȗ
�8v�MJ����}� �?���J�'͛>�T��.U˨#�N.�ϖ��i��%��[�0[N(��\q4A��V��;͔|�/��/R0����oQ�~iu?�k��l��ʽ[�<����\�c�{�������9��]���]b]g����N�+qFXm�G�!G^g+惆몭��� s��x&̵����j�1 �v2��k�ۖ��%���rP�ٰ���-�����-���l�ڰ����:�7�`Z#�+>F[M(۽�H�U��@`Y8{�Y3 Y
 ��q?8�F2,���C��	{�k�1�%��P.�?�\p�U�����O%�!�9tS(�w�Da���#+g�~����
b;jN�|���R��)6�1�3�RɠQ���P�֮ԟ��G��G�'s��s��~�e�[{x�W68�9���'׊]��݅M}���/�%����xpg�p��'lu��eg�'����yz~��b ?���J�a���w8-�/�J����n-~ڃ�N�-U�v�D=$>��/�}��� ��*�CT7u蓵D�:p��32�
#E��qtR�dVH�iey�g,�u%i��� T1P����pB�8��w!�C��ֲ�f�K2�֦J_�	�A��q�E���k;T�E���e T�H��h�8��uϱ����l%�[��.�Y��I��V�B��E����!P���q�d��P{R����u�1��T���`Ej��W�J���G��E�}9���h��1#<��9��?�3��T+�AZ�q�KO��ک��Im��׉(���Qd[ �[:��20��]��g���i-X�rp���o��$��Ib�'ƮI��"p���1렄��9$��e�<�O��D��S�@�GO��C�$�����'�ò��oԊ�l���k5d���Z���e���2唜ʩ�-p4xmw,
�V��v�q^3l�z�"������4�*�{���MN�$f��Zz� ���'�sPq�gMD*��9z�*�t��m��\��ُ��2�����O�ͯ���g�p
��N=ۨ�.��������Z�l=�����;@��` ���.��)\����7Sf�gu 
>'�ڥ
�R]*�I�������=;�Ś�T�$��k"i���͂��3�ε���YG$�/��$��~��TRCh9 �CbvY~����3gK\��mMO_���\{ޒ�\}�����3+�����g)5Kl͜|��X�P�ח��dp��~P3g�'ɒ[�]۪*;E�������#��v7�Th)�/���:F��iUGm����8��P�~c;���y��� �WF�ծ�-�W٣i{�ŃA�q-Ki��Xq[��"�;k{���8<�qw]����Ay����t�&"N������JS�I!�����Ic��)�>�f���-�V�A�Q����w�bwH��e���]�]ADF�$����hйp��C;�bq�n�f���OZD������r=�a������J3%�j� Y\n��k�I��Sv�K��Q^���xf.u���m�?�=����
z_s��X[#�ԯ\�F�	��y�)�K���d�a��C5�����"�� wc���
j���L)��x:x���u����,��zy��������}��q,��C�:6��������&�.�y��������n�1r�2�����<�r�XN�`={�ӽ?H-a/�r3�d����(;2�z =Ï�H��~-��n6	��Ȳ�S��N�f�Ͼ8�Y�a�@����#��?��A��X�DS����O� U;�H
�g5���R_A`?Lܘj� ���?�
<�4���O�t�	}2�ӟl�G�n�8���I�Uss�)I߂�+
�ZZU�o�s��z�n̪��L̥�n��a��>GC�x�`���l ]��}��S_\jן��o�z��hA�ڪ��>�~?=�7֍��ؽ�5��1~i�e�����q	3?���E��5zE���(T��j����Z��u(��H����P��{w1?z�	��*s~��7HUi)��;AY-�Ѱ�64+��#I�H����C�d I9O���2*ָۨ���O ���6�k�Y��t��4+����;�}�]��ӻ�,�$E�V.�/,�������_:p�-Yu���b�
TpĴ�׷CkBu�@�;(��>j���P&�±!�Qu�|�w�=n��Wt�QJ��?x��R�e� Fx������>J���O��SD���c'e���Ŗ���c.,fD���i��v�M[[a评^"�����R���yK�DcW��X�ϣ
����Q\ֻz8@~�n���ݑ&Y�u�`��'�;D�4�c/
Yd%0����8�Y}wPOQ)Ѩ��@�����8y�f'Z5�W�N<�WG±�7E����`�l����%����*�h�.�r�p�Q�	,���D�%�^80��������M�;�pyD]^ ��sZ*���.�{[��h������ y�{HZ^iN��!���A�u�i�A�!Z+�7�������Ou�{��Y�q�p�XK�ϥ�Y���:��I�Ow����������>t��aUT�xN>v���*]>W�"@�q�2�,_���}��E�c�?YZ3>9)�q��qY�R��������r���=-�5q���Ҵx%]ܪг���u��[��mЩ��]:	�S�Ê*߆b�3k�W���6����1��ø��Ft!������E�o1�'�?u}�L�R��v_ኧ���q�8��@�'=�ye����M'��9�(���(�Aj��#�qUIq�Fv���cQ�z=�!H�p2�!!���Ճ�	`@V<T9d��}����)��:�O�r�w�w@�p	�0F݊w����Q��p�ĝ��	�����+�b*��X���v/@5���z�?!V��~�w&O��0�=�/N���*�	_L��C2(|]�Qcn9A������O>DDD�Q��fs��=ыO"�S���:�����R��I=\*H��Q��6�4v��	:�\"w~Hl��ic����Ȁ�.è/��/�OP����
��@1�X�xv�~�YgC6���]N�f�C�A�������*v\p%
���Z/�ʗ��@�\�V���Q �h�}*"��H~�� ������d*As]^��B(>J���� hO1H2���_+96�8���3����: �b<ׄ��e��_�*AF��X`&��#$��7>ʼRlY@�&V��m��`H=\� ��fP������,4R5��a�T!�."Hvf� �������a�5���!W#V�a�gK�ž����1�A��5/���az�ٲ��ںt|�����K�E�Q�-A3W-?���s51�||�4�}�wb2�s��$��G�t����lS�R��݋��(t��C˚����؁�¼���,a؀ј���GG�G�F�aZ���Q��#
ƈ�EZ���=}E�5���+ɹOn��q��Ei�5��s_X�yM��!:��JY�"����Κe�l&�I۱{�gr��<^Ϛ�{��h�H�4���Д��JQ�"�[
���'0��V����t��8�S�@gBa�|�|SQ�z!4�~."�qf~"��9��Gi�A�$$���A2I${xѪ�\��c��S}����aM�HB����k3}y�5P����@�`J5Ak�q�;�ޗ�N�@�c������Χ!���LbG�q/��<��&�zj��5P-� 6����?�8vOf]!ɲ�:g
�B�f�G�2*����8'3/���=Jt����#y��Q�V۫K��Q��U�U�,{0���,�3����uv�}���롿�|)h�aV�e�\;���g��C� 2H�ř�na��ӟ�f��Q�M�yu�����OA�߷
���z�#�\�E��Ȼ�{)��ms�vI�	�a:姗j3$���z����ef��I��8sѶ^l�`��^?��^N��������(��8�-�����H��4/�����/��`6�R�״�D�
�#�q�r�ĩy�������Y�z�a������#��d dś�Ä@���M	bGx���)�����npQ��6%�%��>��Z�+�ɹf�鈍��Xʂ����
�t�d�'���k�D�y�C��@�@B����ѥEt%�ct�[����\�vk���C��AG7z|?E�=;73MF/����-�\W���E�PK>_?x���N�ܷԽѮ%�5��A���_6}���/^;������Rh~�(�j?\^���|N�ز�7�5v�Q6����MM�T���p��k��~0"T�r���ͦ��r�q	�g�zJ�_�ڡ� �m�y�Wi��M��@��˕�G�0���A��xlK<�k�,��嵪�[�k�aN���4�R�I��;��!�CD�	��)���#�J�ĄTm;�r�L�2�b�9��}B�~���6*��D/>5��V�؎�n��ב�̡��4�m���8��C�[{E�Ca������[l�5�yW,{������u�_�	����N�S+.�V��ߎ&oE(�c1�/�~Q�}�e#&Is���;(����B� w;b
;�R���7����jk����b��A�sgwi���C��g�����J�4��	���O��o&��n&��ۻ� Q�Havp`(���s%; ����be�):�KC��n�|>s�=90F����{|B6����X_��/? Zn��=�಩`����T��V��A�#S�7�PPw�J,yԈ-��>`a9�cA�S�Sq���ܠ�A������Nj�u`�p�MLŸ_��Lo�Qyi�/����U��攬��y>P1g j�z�a��8C�0SmC��<��� _U˕��:K��5[q���Mp�r� �e��:�Z�4|&
���R�`�Hw]��僚0t����m87ԏꑝM��PuR��ӕM�`j֜~�V(�Kί�%��ryN?����QU/�Աfm��5�R->���AU�J�W�":?�)��$�x]�t�q�=�Iq:A ��n}��eA�GSLZ������N�0k����+� �60��4��p���[`��EF�������b�����4�:]KwsU��$� L7g!��1�����n��\��F�d���W~���]|sy8��i��bi�3��	y���ý��=J����K�c�u��<��z<X >��+�b�9��߰����}%H{4�jhȩm0oA� ��Q�r��GkfE �����e��T�����/�N�Y��Ɖ�i��Ѽ��X�j�h�1qZw�S�J[>��wp#�-q�H�'�E�q���?s�X�V�S���Q��d�N���,:`��)�O�+]�:�'#w�G���x���x�^��ߡJyam�I�w��]thr�M=��{�������L�� ����4d4n���t	~��4��ֻ�{~~��o��'������i.�&�̫8��l���~�U���}ڔϾ��/�U��P�E!*ď�礜�)X����[RE�fM�+(���6���xBQY�}��d��0�d����Y���d>�(Dp���'��`R�f;�a]���P�c~����nu�9�yr7�/z�c�:�v(W����k�SpՄ�c0b�$�/'�d!�D*f�^�:�����o�+���M �W�8E�u\*�4A��K�q{(;���O�̢��%����џp&5��\B��dM']�Ȳ2i�6n�)iVccb*d��<O�w�P�-�T'��±Ʈ� ��6�~�{*���˛�lA�vO���.��K���!#-�v.m����S�����üEF.j�i��PW���üw~E��m����r�^=���`:�+�n�J!Gt�@�k���n�2����Q-�� .EuGg&"
��Wݖ:I� H� �(܏96'��F��@�4�^b�w[�ɇ*�� ٢� �Y�+>!���UU;.�aV��G2���P�}�����=P��G+FH�D�K�ʡo�]�2�,�GǴƸ��/�K��:�4?�έ�M��G�_0��8󊗊1R�~��Ts��m#��&�n�����-�gF~h���6�]a�Ic9J��K@����W���^/Vɦw�2MJ�*F +��[����@����\6�} �T.b7������yΖ��Ho2nB�����5?@����2K�7�cb\'�����e�z���Յ*H�~�����BWUu:QҸ�L�l�$ynl�����ر�fl�.�R܁�vu�R�n�a�������������hF�j � � j�--]z�����۝���4=�$I�$�O*ѭ����fn\_�xh7�z�H�%��h���J)�{��Tn��=L�����rI(��{ʛ����U#� ��%
+Q�Cf�q��������z	���p�j6���ٱx�Ƈ����ziZ2E�?[bǝ}s[�FFFF��k��I�{/�9�;w��T�*ڰ�N8V�d�Z%������4Wl��)% �.=��}�� �R5V�-ս��&�I������o[[[�e��E`̑#G�#/�x�(T�X���e0nK��� -��m��s��slaA����_�n�ܹ#�.xe��64��w�%���?�F���bU\���\  �5�@�@�w��Ҏ5�n��'uT%ʪ�>o\e�z,j�e�,���Kd�W��&A��4f0�K��'����)3wdN�Ve��]P�}���k�~��O?����|��`J�* �-o�ϝ[o?���wm8<?N�q 
(Kf�{n�Ke�{�7��
��M���[�5����b���K`P�7x�ݿa|��p����0 g��g5K?W:�rˌ��
�`�2�d�W���Z�ZN��Rq��㫖5?'�r|D55�������W�(�Ԍ�c�a�����2�3�nv0��������7o�Q�Ǭ��c��'N�Q�w�m� ����u��聐��-Pg�j8z{.� �e�U]d�a���4�����>/8�oܸ!�0==-�ω��L�R2%[�u�0i���L�ۑ�*��5�.���G���9}�����g|�|�������v[�Uj�Y�+HDp4�_����XO�����
n�@��uB`��GP�㈄dƁxm#��.�D�č��D(ӡʲ1�*
���O_�
���Ic���c�'t���r��'FDq'�#����{�je��|��_�=�Э��99� �����v��_��w���(
?�l�N��GWiQ_!Vqg�{�U����1!�d���2�<�oF�*��ထ�?z'�j���)jrĩ�Z�]
n쯃Zg���W��V���i�)��dOZ�2�ǋ��j�&4��`�I���0 M*�����Q��=����3�W��0����x� ;����0���9rd��#m[C�񙚚��dl ��ᦁ�vd|me �zwJq)�30;;;:��n��&�`$f��<0 ��mSD��(���w�c�]�&�G�r-0�z�L�O��QT������9y���wfmc����	��7lkgk��H��*~�0���fuu�<�У�%4����Ѻ�ҥK����$�$֥|���'G &��y�6�Æx�6��e)����&�z@�n��.�N^=_�8'5L�����&�D`�� R 5Q���z�� "�w��JP@�^w�[�6�sW��#�fn~J�;��Oj Z��-�������������?���O߷��0)�~��������J���^~���~��o?��uN����G2�j��RN���Y[ݔʉ�w�h�T8�ZUg�0*�S�Va����(0��V&�8y���y}2�jJ�jcO��8����E?������㱉q1`x��,�df���-+eh�
bt<���W��S�!��&�A�lll�k7n�7�|�\�tU�� �VWi@����{��
��q��S�����M ��f�8����pv�����j���[ �|-_p�0�K��r����ڊ�|��o~S����Em�UJf�V S�Nh*Ĉ���*e362j��3�N�2�V�TG����9
Eg�'�x�R�����>�essӼw�y��۳"�\nO n��r��.Ɖ���|�Z��a�=��V��RqA@\�Ȭ}����������T��2�H	�w��[�&C�4�Z�H�H�X���RߴEx��'=n[�Tr�Ry>��f��3��±yS�E��!�{r_��Vm'sitt�?�����s�-��ʡ_� ���-���6�Λ/=r�����K��1iD&I%���+೼|�,.�1{{��R)���TG��Xԑ�^F��^������LIp� �:��N�am�F��;g�0�x�H����C�e`�([�b�>�S��J��n�R�.SJF�Je5���:���do��f%m��۠� R0�G�-�X�={V��9;;�/���s��A���zR�L��K`K�hP�ޒ��Y`��@L]���3r��Io������mn޼i�ݶ�$��j�퉷���b� �jT1�s���h�=IK�����fs����C��# X��^xA@�5հ>i-�p X7n^��!(�03�~VsMi_��*���	K�U3p%�}�DaYc�~�T�X��{R�[�!뱻�^A���V$��w�U;$t��Z& �jN'
T�!��d;�
!n�} %ƆB<6�z���ψt���	��GF�1��=z�w��?|�g�������{>�Ӥ�Ow�����=5�V�ܸu�ܺuKb;;ɞךRZi�
1��T+bD�ۃ~-%V�����`0���zG@hT&��8�g�e	�8U�E�,_O3{���H��!�I7�D�����q��#8[��3h�rI��20���Jy`y>�*t��^ZB^�m���,�Q�m��7�bAǏ�4?�������A�c���	i������,^�9BJ�0oG ���!�Ù��5# e+
��OP���q^�cS6ƃ��k��
EE������Ў����i���-�61����=���i%�*Z�^!�a�~�ٟ�����W�c��$%:r/�w (9b�����k
�c��-�l6�`w�]�z�AEq�8�qz�P0��6�'��&'RnJ�պ�f�R;��B�0Y�&V� �Jl.��^B!�t�@�<k��%y�Ҙ�j��5
��Z.���������"T@<�Ƴ�l6��{gfz��_x���ս�>��7���z����˟���~��o��r�ʯ�����1B<�0�P�ݼq�ܸ�u�4��R�q��x)�in�fE�+5��;iRm̡�g��s���D%-�/1�;B.^bB��=�L�Ħn��cl�&�5:jx"yPa�����Cʬ�|��U����ܺ�[&��o~��<� ��ׯ���zˬ��ݶt綌	�Gϱ,����{��{�3S��<&�|8��zl�֠���c}��q�LB�� ��@c,����ᚡ��<�'��B9b�4��0��R�`.R�1a��~s�٘AWK�A5��]���8
P%��k0���`@�-ʽ��n�a���r��O~���3��Ɍ��Z� ��~M����r x/^j���P�G�eAI,�ׁW�I���0�~�*/�9&�i�@(E���Bj�֗��-kk�LX."X��'B���8v��rnH鸖 �}�8�{���v�U�D�$V;;7iN�>e�.����J۔����tz�R�t�׏��7���YQI������=�s������>��;���H}�776���av��3���n�kW��ֶ<�Pci	 � �M�4�G�F�g q= 7�CC���~�30��<��'�CUm�/���ܹ~��6�D3��h*pi�<t��
�_+��}�c���+���
u��8�����b(�Qs��Κ�ꈹu���ko����m��0 QjE��;rT�gN�#4	�d||RO�c����0V&�
�2z=18^��!E��<Ɖ^�K��㼰�,��Ŀ(;f܄�ڠK�͂4�'z8f,�8	��8� ��I!�D����TPRʼ$�,����pn؎�C���z�l�n�L����~�<���r0�y[��eRd�n"�@�x�y�� �ã�)�u������u�t{M�t�����m�����V�s�$�꽥	Þ�J��K:������Fc�:R�X�3FI���"_��?�����e5�U�ޡ��5!Y�	��YaO�7�rd���j������3�^K�K��6ٸ'��`8�������������
 z���v��w�_�z�7�t��F�����p�e���k�n���n�;�[r�R�I��=,���:�T` ����! �PP�-���৉�TZ%���e�۠:g�H�n���@:��ă�����h#L�f~�Ν3cf0�%��s}uM��ˋ�WL���oe��y��7����V�Ê*P�������b?ڪbI�	��a&�&�%��o�m�e���bTNk�`H0�%�I@��I����4L;lo�Հ6��ꈌ�Ynt���9���Q�ò��1C��&m�h��d"xV��{����5ǎ.�N�kF�G$si� ��?.�%���c?�� �k��5�x�����H���
XR�� ��p: ��o�v�)���$�����RhB/��2Cm�^��~h���u�Z|.��1 ����q�|��q-Dp��@r�,������<8��`�X�@�gT�&u�φN���
��<~∙��4�����x`�#�STB�շf��~�s���?(�U��
 :0.��z񵇯\���{��EQt7"fl��v�u�x��MQ��:0�S�J�X��a<��je_\�)�,�-�w��RRf
0Z(����!]�D�C�Y�*�Hk�o�k��ó�B���k�����՘�B]a�9��:���>���J��7W�\1�{��'l�m
���f������L�`l���>��r�*%�c��a�r�FHea&H,��c�s�74mL��$��i+h �yA3�p�l[��H_��h�ׄ�n�Q )"[���' Ƙ�HY�	1%����5Q�G<l23� ��ph�''�^�i*5퀋x�c�=&� ��� ��rD~���8����Aj�� �h?Q?�;�,��ŵ��F$�3&�`A�,xH��6�e�I��; ��yi � 2 T�u�z�
�vdۍ�1 ��D� }�4w��<%=)~�w*��z�|�p���
F�4mӷ�>Ą�{���B�Um���Cɞ��g��Ԙ\#���es�v��{��=g��y�K/�U��
 r�$M/�_~��o���o�z�����S4`�{-s�梹uR�u��l�a�e�5L�A�t@����h��{ @��S��$�g�2㴅7���
Ǌ�i���!�B:BfЖj���l�	�C�އ&�b�؟���| �P��s�=rܠ+dևfq�X$ʩ\|����W�b�y�]��4����wN�;l1���u�h���Ĩl_x��J��};�Q�-��v�DUj�������RC�gs��w�!�#��0�@jH(J$��v����v21�5����F/ ��xh����C��s�[y�L �X���
h�+�ΚqXc�������������ѿ���PtI�� c�A'�ہܛ�|/�c�T�Թ-%l��E�t,m���V~�X'�Ii�2hl����Lz|���~F���� ��7�[�S�A���Ѱ��g�:t,U��Dݞ7�A`;H�bE�q��Zɜ8>/�Pe}��l�q%a*�و��+���/�������������M@ε啿��{�{�7=������3� `�L/]�,	~���+K�O@ES �:4w�f"�����&(�V�Gk4
.��<�x�'�x�C�G[����}`aL5���C�rˬ��c�8�"�3@|�C�c� �߉QHu��02�f�P��L͚7������3����Pm=���x0�Ķ���5�fyeY��g���S��YA�=���ehЛ�=Mʵ1�=$��+7R9Ճ,}ʨ��"Mq_�8��r�Z�ב��oB,��Wƙ @8'P[X_d�����<oEbv�f'4RM;�ez�x�x���5�`� ��dG��ZQZ��aH�o4��بRL�\�97���w�9�6m�1���K�l%\s'[b*Ԧ�' <��B9�U�l�"��7�r'V '
z�t�DO� N���o��a7�ng(tb��7� �X��ϩLp����5�����"цh��������K��{�x����ȑ�����<�[��:�G���8��/��윋����ntt\nH�m�����j"��$Idqk��1<D0�"�X�MA��nJ#h�9i5��\���^����wJ�yb��%�l����E�-/��A��"�(�¸�U2�}�a�H%��`�����-��%�-����*�]�������7���	��D�����4���y�h|B!	@փ��z]*[Ǻ"8��v�\�"��X��[���@H���cc��u��,��
7�[t�����r�1^k�bP'�hl�x����u�a[���Lp�bYP�:	�� ���n�����,��ڈ�'�&����J�B��p� K|Ǚ��_ځ��D�?�!�Z��ZE`y�ذ� � ���0� �7Kb����[���AFs�_���r����ym(.�5��N�b���֡��ɞV���!�	����G��Vf?vlA����Q㪙�?IV:�����ԧ��'����,:���1W��u�k_��?�t���h4��Gp���%r|n�Xn
-�S�"����k$W�z6x�iQ�Xg���:bm�R���%��h\Ѧ����<Y�6"c��>ד`/<��$��ZE�Tp�8�J�����!� �%r$�bc?X����(Ӄ�El��)#� q�n���e'<L�`@��ذ,n���w|�}��Z�ȉ��r��x�s�c�z��S�=KejT#WYol���q�6�MO�����9A���������  ��8�����ȳ�>1I`l��7ܛ/,��nMh8��A�5���I��3�&�魛rc|�	�G�4�zDC��D%S�*E
�Jr6������
�R��*b�rg L�����D�T��q�gy��^@>/�]g�oHr�m�^>K]V�k)��nŘ8�y�qR)�ۑ{TYNī��z=@`���y~ L����j5�J���{�����/��w=�ӛ��= �X�跾�����������yc�
<-}S67o,�7n�� ��̶���4Kp��y<�nP&_��m�-�F ʨ��*�ܶ*JQ�}X�\�؊��Ȗ2�x�8�aQ�Hc� K9��x$�uzrB��y�[s����}l����]��f��=�IU`[��b� "�I��}�7�8P!�����}]���v<ź�x�'�g��'*SP �u�����z�y<H�y�F��񘎍6ԙ���b,H�mg��z�aY.G��Bv6E/D������d3kk�(l��D��8��q�<_�R[- �=�33#X���)s����L���R*EJ��v��b�!��Y6��0q!Y��W���}�cT	�$����4Q���2�$Q��_�ߢδq4T��y������u'�h� ="d�(� F�� �l $UuZQ!/��c ���/lK�Z3�Um���;�S-��r���|���%�����H��}�'������1���v���ŋ3�{�sk�+�M��}�����lhn�H[�}������ݑ@�'x�+�Ff�Jn!c��+2���sAf�U��w(�K��+�x3P���h�\�4�H��B�BY�*�GH ��8�Fm��C�$�%��fvzJ<�Ƿ��m�����s��g>c|�a�h�y�f�K�/1-��,m�e�M��c��o/��fKTa�_�(1�\V���ºx�t�i�zm��qx�4�4l'�yple_�ƺ�����c��0[ꈠ�
|7��e5W
�7�NN    IDAT� �������B��i�l�44V��ʶcN٤���H�pb���GI&����T�hVؖ+<�;++�������Q!���#՘�JU���##�HKO p�%A���@T����@8�Ey�m����;yY�
^�<��:����ց�w,vJ���<5 H��(��^:�P�M=%L���26(J?�u۽�H�M�Ƹ�vܱ�����^�#�fg�M�����h���?�/�}���of|hhsss����O�w�������V���;��f~�Y_�0�+�����Rպc�t�y�`V�[�}T*�  ���*��!�@2��y5���G�m�u]��HK`p�:����b�w�&��R*Á�ZV��S܀Z\*6P �F�b�U�Q��0�_��WĈ}��}��*�#����V�K#�8�Ń���!���6TA��|[�L���=m$6��I�00�y�7���<���Ӡ����
�҆8RvJEYU���h�)I�2oF&*���cCY�F�3k�yۢ�n��c��J'���ƈ�m�l҄�+���9584���O��V���3�����\ǉ���Z�S�'q{�8���e�hTl����K��O��1�Zǂ���6��6v�E*ܣ�^ǔC�3�'@1 `PhH�m�(��cb�N=��@�r�Uc����ʳi}<cۖ#O"U���d!{�y�����Dp�q��w��5���VQ����K��t�V#Q E�Ԛ�>O�Z�.�8GL�PI ����K�R���_�G��c�ڒ=���4-��_��cW�^�'�^�3�vk�������)�n�ͅw.J#���+6خ�x�q1`�ټ��2 ��qsf h0�Ԃ�K(i�H�7���X�$��ج{,�Y��,��Fg�9\�.�q�J��x&FU���A���:��x�p���:-�LU�i�Q ��i�C��B���nO��Mx9��B�nm�f�!��<��H�2QA)�]3pH9�њV*��!.#@m4��	4`�ݶ��ZQ��I6��Y3�N�,6�׆q�yU*�͎�U������q���w��rL�x�ó��`) �n,�H�	t��V�&��3�O��+R����e+��0�2����L0P	cJ�T�H�^����^��52�����Q��X��1"�D���ؤO%Ե�z@���ʢ�֓��(<]m�.4��T��3�*(ilQ�N/�Z����g�/)ہ�c�����(�������8�/��<;RwBs�HBn˵���I�� sD���@7Z58hl�6/G��������#G�=�]U A����߹��W��[������'`7�w����T��r�YFS�����	�%i���t6i2?�4�%} ԛU�	X�ڋmŰ��r�ό��K�*�HA��7�-髊�)�����`���$S�b���c�;==+Y݈�����������G�偄��v�{-P/4M�D?�ؘn�#uɠN���4�[Z�����c �/N����!aG/�(�8
TyBJf�}2hOZ�
�z������!3��~s�Kő��6�=�S���cM���8F��#DZ��zY���+#�9B��jki�d��ሐ�ٶ ����x��()��`��
�8::2.�(�7���Ԍ5[��fe嶕E{RP� \kPwx�sU(�U�^Ӹb5/B�b����B����A xzc$N�j��  ��L���9^�7
�a����XFM�ή���ޛ�H�]�}��z߻�u�}83Ԉ����)iHm��E���b٦L�2b�NG��X�b#1���c�$0$ �mɊ֘�iqH�����ͷ�/�U�V�{��T��	�f��]���������9�9'�#j��u�Z���܋��sʾ���g���^Q�m �ͭV�;����O���uם*�C�W���ݝ��vr������~�������?���.,ܷ���}�)�s�r�g���Ϭ��<]�塕�K���i<��r��Ry���Օ����!0F��)C����1E�U�et��JQ&t��\R��1ihJ����D�A'm�%�����Q%��N��A�a+L��x V ��h��{�1	����#p�;��c���f��+Au�����j��ղ�t����m����Lq>({G�;��FKH�1,CB���g<H���k��C�Â� D`�<��k��x@��&K'ǥLO�̄@R��
�(��nK��Iճ�kݱ�|�սH���=�^�{�]N�a$���b��xy(���T!�/ ^�]P����x\9+'��}]�~Q	��<l�o�߅�ŘoRu[P���)�bx���R�O(c"�#�N?%<��=�o��mjC��o9�ɜ.����К���Ϡ
C�L�/&�BcVTϿ��!��c��B���5�z�ynQ@0A9O`=< �j���n9y�D���JT�Z������-5J�3O>����x���}�U�E^�R
���o����ɋ��T��x���ݸzSm~�x�v�Fy�����ke}cKTVj�EȰH��UPrz�Pӂ2������*�{lXY�Ux����(��_��\��֥��3�H�M� )�rjm�A���{@g(�٩Y�bmu]������ccL%k�C�eqL�]X8&d*��5D��r��A䮭����%�o��k=�{P��VA<�J�a�h-̀N$X��̀��!��}l�#�vdT�"�l��;�ji��&*\+�f��Fɲ��V@Q����qQhɗ
(1���^i��@w�k{�Ճ|���?���*�����p2k?�)��dǸ���\��^�s#��A��	ؔ�X��x�(��M�Rϰ�cu��s
�.�ȹ;�"{h��b���T9Ap6
p�j�1�P��DU�!
��@���`�*�Z�8��2���x8̫;�:�C�Ӥ{�V�����Uw�����&��DJ�ّ"����M���*0\N�>UN�>!R�u�\(^�x)�ˣ����ַ~�?����W�F%���з�Z]}m�K_��{_|����h4޺��>Mi��T��m�.].׮/���U��ւh���$�Gm&+���ů�^����<�f����g�Z!����Hغ���7Y�$��6%L�RI� �V'��%<���L͊ŷtsEx?[�P''*4sL��ƹ&���p�8}��^[YՆ�ú\^^��g��ʊ��7�7�{���-��6��>��<d(A�Y�ʱ[�ӓV>�D��c�W� d�x	��;���\+d�xA����1ĳ
�G ?U��cA���P�Zܒ10_Ε��NGc�x�Ͻf�thH�B��0n���"��w؋I�<��9&
tƫ\�VG����R��p_2�{��.#�+U	:���j�~�A����x��H���|��Ha@96��	Q�MS6TLusџ��n���jl4^ iؙTs�'0�m�p����א����B�+HG������:���q��v޹G�wح�HQ��J:8P������=��U��هN-�:44|���:7<<��O?��?z���9��W=��o	D��g�=��W�����������.^�p���N����NkW�P`��R+���e��4b��h��І<T�PROk��F�L�[R���e;�
.���c>@k�\Z����z���=���	�{�O�E>����7Q&�'em�it[[xӳ`��d�;�1�
!����m'o��D�!m���zη�Ӗ���TV�W{y$lL�9T�%����E�e��*)>�q���g��0h�Z�[�����"�y�㑢PӒa�DL\s0�L�pD0F���9�E�%�ٳu�X�Ϝccs[զ��1�S����P�n���E�S"��b���G!\A�f���Pekq�ǐ��ӛ�������M�F��d��](��<�iӹ3���D\KNkMm%\�	O�r�� �A;<��=;;mx���Z}Xs�,��6;$��d���H��P}�=�¦V���"�'E�s_�$����������+"X�7HRhwH7hW���(�s�m�ʜ��s�⭭�N������Կ�ُ���|���+(�o	�կ~�M/~텟�~�ڇ:���b)����l��*/^)7����@1��Lh�cI܇EK��Ee(d�'�����1+���$As��|�E��� ��MG����$��k蜃^�`,�IƼȁ(,������-�L&��J��yǻ��ó��_��V	��N���7֠C)f�17�n��KeskKTk��tۑw1>����w$���R�%$�pr��)����;<G,�H��B��� a!�R �Xȱ��H��W��B�p��Q��|t���I�JD��?TE�Oy�wܡ5�2|TB�F����kqn���%��V�8��RZ�*�I��<\������η���ضZ����x&�J�O�\=<��+sLO�nU�IL��˱�n����{߸���1�g�t���TSU�}�Zb<�@;�#��$�����1��{Y���@�۷b����������4K3E�F<t��nm�łi����kfp7�t��a��ͽ���=�Ѓ�����u�=���ѕ�^]����������7������7o�h d��8^��c�܅�R<�._�8�96,�l�Ee��l?R@�ڀ��To(���c6�o�`�C�p�B�5��X�`�������'X������n�xV�4��h(gJ�#�H�M�Oޛ_\������ �m�#2=��'����v�qݞµ������PI����{mT�^M�����BLLB����yb�4��������.{H��J����5~���1�BT@Q�I<�ɹ�V(�3��p� O�g�1ʟ�( ��0��+&#��8/��k�#,m��t_\��s�{��#�����έ�&xDТ�X�|�X��T�J�����K|'�<� k65���T��Zm���Z'�:p&�r>cM�������K]Uڸ�6%j&.�g$���3���>��޳�{�/�Z[ h,���'��#ʳ�#c��\�bʍ
�ޮ=��`�*��(��}qm�o}cU�'�8�y��^X��E	ю"��+R�����/�����O?�֯5�:|����
h}���g?��|��~vdd�V�5���.�̱��*_�岼�.K0V�y�b9��ްhd���F���LO!$p8�Eo��qj���fa8a��Ns����3�/z��5IqS.����",��Z�ڙ�l,��A��DL�E��8��a�� c��D#�0�N?�͇B��z�7��Χ�w�BH�i�ʊf�g`%HBL X�4$Ʀ�y �y=R�z�W��#���x2(_�!1��&_�bn�����Pѓ��q�O�+,R�/��!�0�q~��S�V�JZ�#9?�W��f˞D���P��hy�yԘowO
I��v[��ob��P���)��jX��j��F������տo�	9"�6�������3*9���ףS�h�
|&O�4e,0g�yF�Z{�+^X��b�L��;\���c��o���E��'�I�3�]
l���a@��<���)�Ѿc�=B�*%����b3�Ϊ2bG(eJB/kvj�ŀ�<�99~jj�����o|�}��o��}�w��{t[oX��vG>���xۙo|�on���{owo�}dd�<���j�u���r��M�R�D�� M!p�Ւ���̑3S*�`Vb1��u)O3�e��`��Z��U)�����%,h�"�ED�x6�U�v�HUɱÆM��6��9��I�( �M�{b��\Y��m�f�ז��W�'�����<��9)��7o��ׯ9�?b�1��d��>L�F�R��jN���D�Ͻ<��兗^��(
�xb�37@IO=��~��B���b�ǻ�P��E}��3���[j�q,�Y�cc�۾��|���=�}�ۜ%�lc��DԒ��dZ3��#�|x ��xy7�l\?늱]�|E��s��MB�UeE�	�[(���F`85���o�����-�����{��Wo��!߁v�|T5�����Bj��B�Da{V.̷<���������r3��O����~�<}� @g�N��&o����b��Ǥ�x��0񄔯
�W���b��	��s��Q��]#��zv���'N�d�}��%(�|>�S=ƃ���W�ff��O����o>��MR}�*�3g���g�������n���K�癙��m��.��W�������eh�l:l.p)�"��N���D�q�l6{:�c@����8�O�I q\}8��q�� 5����8.���Ԍ)� ��#��+l�:�y�O��n��>��s/���؇��脰lY{$VVE�t��	o:����c �yb*x��W�hln���Ʊ���=Ƌ��/��>�K�}Ծ;�ɵ����E����C T�ww�D�f�g��˘���.W�=����M}�|O	���"�������hȕ*�u��0��O`ީ��o�p���
4�R�5d�l%IK���3�Q��i��2E�=�4u:1֭c?�0�=Fƈ��r�u��jn����q�C�h������Q98rbi�1"���B�=���ZE]�$P�j��^=�O�ք!�%H#��d����$�Eb���K�d�|�l�H� ���R��s1�ڑ�[�吃��n?}��s�]=�
��[�_y�[�������ϽQ{�!йs/���W����/}tww�,�˗��c'c���kR>7o.�� ���g��b-k�%�Q@d�+�߄�KR'젚�c�Y�z4��������Y	Q�߁�.�ʂ%��3B"��7�I
�������uX��Ai��BH�	W˖Da���V[a�DK���T�- 7��3&xqH�$<��׮{�m(*)�P�G32��ӣ��`�)O
��핍�5�Z����l��󘟵�f����P�x6��#�	ٚ'ĺ@�p-"��'�]ES�?:P�E�2�z=O�Z�Q^xcQpj!���@Y{wGl��qy��[�n�)�z���(;[Tl>��LAK,~�0��&[�\��<�:�@��#�g޸��y#��)шC<Hⴍ${@1���0L��z�Y䕵�eh�n	�ǳ��1E^��,�
B���IH��Exg�]LQ0(�x���.��w�(����ʐk��y�{����P��;���[X��� n�Ь8� �Y)���`@&��!�Z"R�7>�0�DUָ	$������-���{������7"��S@����O������/��v��'vww�^;s�;y�L�O���V9w�b9w��Aj8��\Ϯ��L�L
2a���Kuk�iB���1|`�"3Jś�4dI��A��ϾU墊X���������4\�0�p����з���	St4V,�t*5r�zn|���:�B��X�Hd��aS�h��S��\aa�p��l�����A1��
fs�f�a��<�(ňFkE�=穠��~PX�j}4b0<��|�ga*h���u��x�,��S�^�X��E��暬�� �J���L.��f,�2:���W�����P<.,����29��
����ty�ƥU,�v���;�p82�y���fk�Ѵ�
�����=ø( �1�Ե�ibV*VL)��}��I���>VQD60�i��}�51�0/aoO��&��41@��=֮{�R�ăےBҾS"�ۤ`�%>�V=Om$LU�{���k{�rF�Z�(���)*�W�1	12�]�]����
�u����B-R>�Q���LYX�Eԅg�1���p�n����/�O?����7���M	����=��>���ml��P��8��3�����Ay���ʙ3���.��Q�Gv�#�F�G���M$�N�ڵ2
H.�b,����*�~��^�(L{���-4k3�*0X�.�o�c+�
(�y`7UI��{;�ǇH`O�^�W�Қ �q�A,@�� m*�AAЎ�0����L@�k6P�������f��2$761e�    IDATV��{���k�
�\�<m��[Td���ܐ�;�fs�ej�I�4�ãY\�#���+��~@���L�-�@R%ZI��p�o�s�B�X �s�uS�@iɪ��8�D�������=%���ڭm}�]`����mJѡXk����(��K F@��7u���W��0�Z-�tN�5����I��b�k���V$ȧ'ݚ�J¢-�~Rx1^�1�b����s��1�;��σ��QDXbx�������3K.��<U��{G�7Dצr�OC�2Tk�ԍ��U���C<%<x?+'A���_u�0jo*+'��|_Ŷ��n*A�]��ۊ�Pk���9Z�=G���F{CGGjb��{��a���}C���������KS3����c�x����y������;�7~�goܸ���>�5q�����Ï�V{��?wI
huu����ٰ`���P��������b��\�[��'�i� �!j�X~X����)YP�w,�R$u;h��V�l�@o�x������q����$�zYi�o:O&̨$�� ��P�k��cY(�����#BA��6\SL��#�@g���r�ޅ+]S�m��UZ��e9�
��0kڛWL��y�I 4\!�杖g��x��R$��1�as�Z�r�Ry�'�� �����u����,J��E������Uգg]�(�D�^J���r��U{��^?�\mmJho��j^O?Q�G��ǋg:l�<,̴~F�rn���+O�d��k�`+�G����ϔxۢ4ϐ��SЮ��Ã��ʊc�C(~h�%��PjsQ+�L�����g�'����.��R榖��b2���̺�����:�xR��x�1��' 7Z7����b�w�V�!�P�E��m�����PU`�޼
p�,ѱ�B�9�ʊ����}�R�M̎N�Ě:{�ҩ5�|ܑ�y�{��s�չ�'մ��#5�U@a����Ğ-	�ccc������������'��h4��� �7�ZZZ���?�=/����l�7�<<�qg�cev�xy��W��s�
4�ͭ����\9�����dfS���*��8�T���	�g}e�`%F�`�$�?В6��.P5�A`�_
���a@	%���VjS��`�7
J�K,k}���y�!%���3[����ʆ�(D�EX���Q|��x@3����F�=]���G�Pu�jmrc5g�1�a) yo�VX���5��k��PPT[���mY���'��p;C�0�8���`B*��� �Q(�� ��P܎�tG��`��W�k PμzVמ_0�6s���_k{S� J3q�N��)r
����667���S'��yV����K^�������☍�NK��R66���a�ӓ�q@�;� 29a��p�F�
�KL5����� d%�^�uȈ��Ԡ�W���wy(}U�o�J�3�{[x�=�P/$1H�w:8���P�w5��5<��]�{�Q�̯�����g��l��Tő`qV�v⡉EA��?�I����_��
��y7���,=:6�rK(�����Gy�P��J�#prb��Q���?��?�߿�m�~�@qo��v�_���>�{���ύ�5���K��-��;~��r���|�\�)���K���U�57G�g%��_=��^���*r��( Yy	t��(h�@o�ׂ���{GB�b�XI!�P�R(lN��[��@xQ��t�-'G?&0������~QSo
�&{@���l�CE��|�Gq�h��6k?�3:1�cQ�xfw�	�;�f�M�	� �˜���􌒼�{P�4���+;9?9:��� G� ��AJL@�����g|'J�k���r�T�f,('��}��'��B��s����9�(/ދ�V5�]j��8<:g╠��!�l�g����Q@S@=�S�܂�D~q���3�u1X,<-��O��k}��)#.��~}6�?�5%�g��y�õD���O(��kS>�q��a:�c�3ϝ�i���8��WG}�4&�o{�����)$"3A�66�[!�R(��RY���V�1@r!�J�%��F^��f�ФF���x������ZP�Q�k󜀆yN��Q��0p��'zv/u������>?;3�������7J��7����s���G^;�ҟ~�B��ٙ��j��������խ�S�H�J���B��&�7%���:0PĠ7�b(Ձ���VW�ɞ9:Nf��g�p$�؍�*6"%4� 1th,\y��+ܜ�6�H���f?y�����vГ���tS��&��M���D�y	V+�(o����.�J���"���9�N1���L��(x)���0�m�=�N%~�:�TXV�Әk�!����$h�F�o
�����ż ���{�('H	t�e]�܊0fN9�����#�I�H���Z�Tl�	Wi .D�CB)p�	� ^��nC�	��%}8�4��5F�������o�y�"��m�1l�����b�9�~6��Ԋ��[K�pE��j���N������V|j�� �K���q�
tj��Ϻ�E�Y������`�8�WC;οQԦ���NK�h�����B��)9+N���xn Q:ޏ�϶���pI�����>�ov����:�y�1MN���rǝ��-36����8<:Z������|�;���ǿ�F����W@��^z���n�m�Ӛ$U�+/��Z�t�\�{a$��ېJ�$k^��Z�`q�{�D1�Υb�B����}O©��}��b����,L�Ů�0T�*,`ޣ]��@0П���}��TJ��(�Ob=��,�,�n��f��cK0�Xe��`��QYF]2{q��q��]�A���l"�(��^�w���33��}mpF�*��R�&� ~�./���( �bQ)�5{06\az�̙��3w10zl���X�@<�(�T�F	�8��À�^Q(�{﹫�.��Dѥ<P#�E|�x$���a���u%��������Ӄ>�#�d�!�xq��`H&�^�ށ*.�}b��PLj�����0���Y���`���J�P��V�0�`bZ�T�oEo���;�#���[��p��.:����\+�x���
��C�Q�J-߁�BG�z�W+�w�}� ��U�A�eS�m��9�"������HS(�	�6gM�rߓ��IgW�Ó���9;���l:�뮻o����&�f��d|vxd�W?���O<���	z���V@@o/}�s�~��>�s[���k4ǯݸ*�0�V�S^|��r��R��$IoD��Y`&����y=�d��Yp�������X��w���,̐p���V�|л�Mefն��[���"hZ���b���+y��:Cq|������qL ����t�ǭ�G�x��8�N²Br(�4�b����8�k,N�C`���+ˎ1p��f�I�q��Ǜx�X�Ő"�L�$��X]��a����.�¼��<��<߮n�&朌��8G�2ʄ��/��Cy�},9����B�
6�A�gg��9�y�90Ox1.���]��@i0��6��,UA���5�W�ϼ<��CU�8] φ�6�����g�������5�^���W��X����ﭝ-���|���"F�y����gr��!
(��^��������_�"�u�PF�̷�>Cq]*a���=�u�;��f��]8�M	��%wD^ 	�O!���Yl��	M�;OD\�`E"���Z3��m/��S͡�Đ���{3}���xF��Օ5�?$_LL:yjQd�c�����Y��y�Z__��������q~��]��u��nܸq����?w��O�nyDq
��^(��^9��y�V׶���%�	�"�f�m�gc�0��BN>Ġ���̎՞ŕ���1b�-�Z:�!�ȋN��.��SYJ��w�� �	�*����b=�؍;��1���y�A�pr �U���\p�zRe��e����>���\�6��n?�ް՜J�\���#yq/�\�<VQ^�L�7���/+�|'�oCP#�����8�MO���,4C�f*�?׽p��q�$��,�Ikrʸ�,�*�&Q���;�2�̟!�y=3�B��(�=�g �x��?����!f�g�8P��6ֿiM����R딵�e���|Ě��:���|�r�*ǜA�¨+� &��g*I��(W*:�
w-�jcn��Ԗ��������[�"28�J􃞆�{G~>��+�fe�5�qH��`��c����) *%��1$ř�
h��2��r-�Y��s�����2�'/tcS{�(����)Cq�N�T���r"k5�������O~���ȏ�����$_g���Vu�/�~�K7���>������L--Sa�v�R�x�jy�ճb���'YΔ��6��_s3�=�d�����1+�~`�O6��̪�8��j��X+*�ߡ<Q@,�$��ݯ�iN��S~�qa[��k S��#��%�͈J�5���Ʒ�G��s,��;�r`s���XA��R�J�8��A���fc�Aؐ����<Q@�
^9M�rlX�17(.<����y�CѳI��z��G�I� �$��y�(1�jL$���QW�0e�J���(x�ͽ�D�'4�(a�l]t�X�Y2F\m<ωs���u�����Ü�XI(?��TY`\|�c�o�<���ko�ą�'An5��uO܆؞	
^$�*u༔�T�h���"�bD�.��F�#i�vm ����3�:9Mcu/e� 5;����l,i��tP�u��g��@�T�W�	��׶�6�~gWD�ճ��,�V����Bڰ2�sm��x#�w]�񤳯�UEI���q��ӯ����1.��А!�.HAJ`=��X�:6:�=<:<;>1��?�����o~�_���^�
�k_{��g?��cs}�CC͡��4	԰�p�\��TΟ�T._�Q�v�fn{��O	~��iYtX�v���"��0��d�4}�_�Ă�/�v�J2���Wa6��Z#&��=!Q�5�q�z�)� QIO��b9��-C�!\�]��������҄k������T��wv��c��)?�[<Hs!r@�i����<��U��Е
x!�mm7�\\����O�{D #((����p��*	�~��^yE�q~�ɉ�E2�)�(M�8�.�-Jz��8oj�,����[!Y0�(���Z(T��Xb<�Ϙ{�=�:��vQL�'1(�#�
��V&�!/< ����%܊���걩���c4�z�]}�x�x�"�,����mډ ��&]�F3�ı`)&Z=���Q��(�x������Q�E1Cw���H��Ab1.ݓx�b����7�}O�-Aו� /��^��Te�)�*�@���b ��d����)����76�+�Ɋqb|T
o��t��.?24�UJ�����_x≷?��C�϶�K��qi�/<��g>���ډ�o���$�LOϕ��ny��o���5��9����q�ټ���$��z�ƆU��es�=N���������p���N]���y)�Z��(�Ө�8c~u��H�bB����у&�ܓ�B¡���m��}t��
���NͿj�vJ�[%ےs|(�7!��w�˵�j/=�77ʃ:Ty�Ā/ߍ��w�^0
.w.�㝥�5si�s��}$o'P!c$c���a�9_bUQ̙W�++��q-������Jl/��V�ܰy��ؐ%b��%�`��'{17Ɲk���L���������ړ�s�P<�M oi�0B\����9>�Y�Z�A�x��I֮
��)�	u����q �#�m�t��!�;�ǆ��ks=>��-���]�A@�����@��.���29bq:�Ψ ^N�gTQ����<P@���?��keqʾ�3�k���CWB,	:��*XzH�p���9�
T�<��a��uםj��Z�}حb�:�����ԯ<��������I��߯;D��/~�SO|�����뛫�j̱ &��Jk�S�_�Z._�Yn\_)�fp9��"��cr0L"%l��9>��m����F�z��^6e�Oܪ����,�X{���xe�Y ���|�p��L9�2�J�-���,zJ�(�x��a�ţ�Q^�I�)9�ťMQ[9ۢۗ���ʨ�6{P��Ht9E8$6�x�"���K�h8/��9�m�� ���$d2w��2�����D�0�xs͜q��|2v��g���1�?�0��|҉3�/�*�!�?�x;������ƟB0dhH+^Z����}����M�w~OSP����8�ER�v�PW�{( �	i��:�
��y�##�G�W�Ɩ��i��{To*Ǐ  !%y������y5��8a�)F�G��b���ffL׮-�k�U����e������_*0�$��+��Ny��-���	AJH�+{��S{p��#�|�*	��k�����1�1>F< �!0/^��Q��t ���w�Q��n�	�������=*�������O���|�/�����뮃��N]����}�S��K��h<p����fsh�\��R����r��j��n+�/��f��d�E{��x�ӨചX�"�"R/�~���+�3n����D���e�x�);��[ݮ�FGV�_�����rQ���l'^�����LC5�P1�Z#�s��4	�TA��|2h����7��=(�7:غI(�TȜ���( �-1 ΁�O)|Wמ�v��O�!�=Z���#�# �F9�:��x%����f�GX�{��x�Q�|���}'�DMY�5�2ā�����m/ɉ���8�k�����޳ͽq�x�x@����rg����ӌ�г�n�(��a �Z���u؇0}A��U(p������x�B��RN(�\h�Q�WG��s��jA��.�k�s�ر2��v�<߬��T��0�k�����T��j�;�㘨-�^^��T̯F����|�����d�~���r���m�b�aP�='J�<?J��w߽�g����w��l�|����_�Ї~���7B��Ju��&>�������_��k���iNu���l�W�\*g^;_VW7q�e�C��0<R�.�/��@QQ�J��c/e��'���v:�F��
5qA�vr�2��Oۘ}�n�6q�c��[c4.4[�']�:U�α~��X�^��|.V�&�1k*~(K�kX'J�Z���=vL@0̡c$]C� �븏7�n��ڵh*�"�M����aA1O.dEiOɞ���â������XU^���Z!�=��X"�9�k�xe��3�ߌ����},T�uE�~1X�e��c ��vmp0<�����J��4�!����0�8(���1J�8_(�'���N��!0NU����f��`/�1�P!b���8=�ZKpt�i�D��촁�J;q_c#������GV?���!�0"��.kr3��kĤ�<;{����,1]��W)�i�@�5U�F��1���Ӟb<��ZZ�R:�+#^���<_!{p�5!-�mf�ě����-�H)q�#w_�ܢe��j����1R���r�=w���))|�Ş�p��h��v��������O���ZOc��x])��^{��g~��msk������r�Y�e��9{��v�BY^�,���asb�Qf�����XoR65�I^fb@Y�Q@�����˱��PJɣ�4���!���Ǔ�h��2<a�����N P�u�dI�K����M�֧�L���M��¨�R��vZ.uH��@ICb�5�ؤ+X3��$R%�]S&LD1�'���u�ÈR`lȱ�(s"�nҭƳ�0y96ʞ�ð���9]�0�t�+�N0��%s�X��5��qֵ�@B=Jސ�s���*3��ʑ��$.�o_�9��M%��!���Xr�=?K��@�ㄾG�(&ߋb�r�b(�ߓw?�xT-�V/$	�ZBg���g;Y{g1�����LC���LBA)�tR�8���\*�;�<��k�à�:_*�u��    IDATpmrsxfQz6;��f�t\���}{C�F�_�SW�$ϩWM��@�TqL��bڶ�I���Ey/
HhDO< �S�ϣ�颀����m~n������{���1!H�V����w��������Ѹ���u�z�( ����o}�]�x�号�7�>2:4j�5W��6�W��R�r�z��v�Z��O�dAOL��c�/��!<Z!.����� %�!��p�S���c�=,z�᷊��u2*/m�T������	»��f� *6�rw�l)^ʠ�1�=���qBV��ڦ����k3��6��!���AN�*�mUY=�8��;tv��VEFŋ@�8�o�tzr��mHX� ��_��Ĩ��h���Y��oVJ�>��Ÿ�p�74P���D�y`<�1�k�!<�Y|��s��"���sb�'� Xst\�()��q�y>�0�[=�j�s= ��]-�7J�U8�F�r�ĔN�'�ʳ�J�����Z&�<*;5(`�C؛�`��J�LK-���}=��1���A!A��δ�ܕ�c�O؝�^�`��p��m�W�W[j�EH�+4I@J�vm���s�>cH�y�Fޙ�x�����:_�m�1��jԼ�2E1"���nG��8~��I�x����p�J�{��i�(��D�S�g��7�~�� Fۆ�zP�oQ�i^������^�v��}�c��o{�w��:�=��B����ٗ�7��k�I{g����w�`�s{{�\�t���򙲴D��R�h�[1R2�)�y�؂���@qU�+�[,����b�
��"J(��nqU�d�ۺ2T�vƂ����²1��f�[�*�V6z�N�R�bN�IYλ.��ƒ��U����v�(��g�.�(0��TX+]�z�Y++3{xa��ڮ%y���bʟK�X��q>U���͂M:�Ф�oC��r�82���@��@��A/%B815���U�p�@H��琠<
���?s��C|&�+O��o�}6��N����/0��Q��&��~��<?2��?0cV>Q��RbC�3�EC��6��s���5�����܏0��Z�ı9N�~�"K���g�i��w�k�'�.1�x*�33ݣ�s�����NK��o���uW��	,��r��\N	c-/�==���k���\������su
6���N�d����J��)�@^�0%��=��}���}��n凡l�*�(2{��Ҵ�*M]�2�jـ3�
ȥ|v;{�����O�8�?}�#?��/.>��zPB�t�ҥ�g?��_�������o�i�bOL�H�v�b�t�F�����k蜩:5&uan��G��,Z31���b�bK+$�A�mp�'�d%a�B<�C.@�8�4k�X�x@���gG`b�x�ǂ�¯!+�7����a����R'ΞL�\�z��)�݅:<h=�����|�ւQTu��$��?�d�Q���0;=���\9��4��?��vZW�|Y�5ɐy���w���7<�xV%��ӏ�E S��܆�s!@��ƽC-�r@�ʨ������h�\j�u�|�y��)�����%���-*.�7�$�^�
����1�V�V�������0�!���x'g�[m�u���06�ս�G�>��)�	�l����5b����1�`�����+�Иnvvƴ{��T}�
�N�_�Dq-�˹R�4�hb�k���1�`yW�l�'x��'l3U%�1���5S+!p�F�ώ�)���~�Bn��	'ϳ�7��*��ǆS\�m�6���64!��Ow;��=u�Ա������Ng[m<׾	ÿ��w?��y��^����<�ܿ����������������Hhlmn��W��7Μ/�+[�i�=j�{�aR�y~~VL�`�dB��͸�������Q��f�P �e�+����6�k��*�$�Q�>�P`}�3,(����D�,
%:A�z(����mjae�2��Ehe�F���7�0�V�~�}qبW._.gϞ)��벰�B9�M�p�_A>-{s�,�\ฅ<�1�T�v�Ĵ�3+R[�S��-a%e" $�c�T��p���-�8O`8�U,(x�4i�J6�"�ܓy�3P�������ګUǳcnV����L	���3�`@��H�VN,�v��;\��<:g���-)��8���9�
{.�����A�s>K1R)�#?'#�F�|����F��c'�*ֵ����t�CF��^�\����W�0ZL�ܟ�	���D%�N�LAC�ı�a�����ḱ	>����l8����񀇜��ؓ=Y��iR�������zާΡ	9�ٴ�=ۥ���d1��Ą�Gld�k��8A��s��	7�^*# �%~(��KӺ�q� ���.��NxgC�2;;Y~��A����*�s�wZ��fs�'N��~�'���e�-�mn�r�_���s+�+k=B�tXc�����_}��ol�ｊm��I���N��	��@ �XDS�S�,n)�aw"�⌧#>��i��Ή@DwX�8#���ؒp��Pzl�Ъ%l)7Bhb�����Z�%p�E��X�!l&��N�M�� о��(-���p��e��E-2j�ݼ��K^�btXJ�VpW�B<.�j"���1)�Oͺq�����k���?�]��!roIȍ��@p�
x�x$!;�<"E�H�j��0�8�s%{�-�!D�kW���E��b��+"��>q\B������_�Ry׻�UΞy�|���V�ů�Z�η����H��1�(���x&T� �tX�X �R L1őa	}檵�zpj�V�E2ˌg�@U4�/�
64V	�*8Qt(����&���V޴.��@ ��_�yf�zr-y�G]11P�S�0	������TUs��L�����*��}wv6EZ���M�Y�M�U�;�5��;��ͳ�rb_�kt|�T�#�f�|imMc�]�[��Rn���8̀�꺵��(P����Q���U?��*�kQ^����!K��=2 \u>$��Ξ�,�lT���
Ů-���~G4w�dB�~�G˝w�.{���m��NGc[ZZ]���=�y�o?�ԏ<�������V@T���~�-_x��o﴾�1Ԙmv�c�kr����W.���JQ�~7ԞbQC�f��+�Zt����D�� �fK����$�ӏ1D����:�"�f��W[sã�!��W���ł2ع�q]D���WV� �ږ�L��g�(��Sr� "�	A\K�ME���/J�e�9�0��jA+��yXC�tâ\��n8ދ̔髼���,�Ѧ7� ܆�<j�X�I��P�9g>�3�1b]ո�a� �/K�V&Hl#!�2y����@��(�s��*�����W_z��hM^�G���R����O���H��s_*oy�[�������F9}ǝ��m�U�RWզ5�v���I��V�bF5��B�cc�-�ˋ��;�p�t�QA�ώ!��\<,)�Z猿�ڙŎhD��VW2"0`��3K,4U�]$�*��g(){�.[���!�t��w��kE}y�d���_����s.�˫�&urڹ�޼�"�e<!	z�fw:��j|�����cOh�I�Ą�V�C�A�kB�J%�B�Y�����Ђ�&!��7#����
%�=���W��rW4)]|��|���=�������-C�C) �	�iww����9��p��������߾�G�=�N|K+�k�^=�O��G�]��n9z�7�$^0Z�n�����r�vuU�,d]� �~4�*�I�~?��,L��j��q�Q��X�_*��gQN��O�:XtY�޵�ΐ�1&�h �#�@�!����:"P�vQ@��jr$�brUg�Sp{���/�N�x�\�vS=r.^��qE�a�-��2ntk�M��4����|:�B�
�6�h��@��
��-�<YH�����}�Q�z�����P"��@	����EUf� 솀�P�2.�;�xn_�җ���Dy��'˅�������\<�$Gn1	���-'N�Q����'>��𣏕z�]d���t�b���n;0Zc?��h�F�5e˻V2�!L /^�3bD���r1���t�hR���9/ʹr�e}������]��)�c}:�ckp�6@��@Q�H���wP@<["�=���@�9��mz�j��i��H�I�-`�/��hM���~�F�O���IQ%�LFU oveh�|H9�m�&bb;�-Fb͑��W;t�B��nX�f��k��%�ň�Pj��ףg�4��y1;!P���\-��m�7Ӑ؅��n/���27?YFF�К�����������g�������������#;�-���~>��O~������n����l̲!ǆ遳_.^�R���+ek��=���y�4��{(��|6<�R"�_q��X��Q@>O�aV�2��a
[�r�Zv0��G�}��t��Q{��+K�����25�$��_º�R�p�r➘>UI�\�\;q�$�r��7IMi�t��T����jU@@�QT��h����-U�[���x1��>��!ΓxY���s��xC�PL``������p �}n"��2>ϣ�&��訊�>��7陬./�o��J�|�<�y�5m�V��y�w>!aq��u%�nm������2=3'�09=�k���L%����iM�$��G 2{�����-=�4���1@ZVG�m)��n�=���֛k�FZ왐
O�#]!qG�]�0q�x�( fz�@�5�!M��z�V���S�gf��J��Mڐ�|{T0�呆a��਍'<0�N�.$��n�gHO0+'�^F��S���219ꎦWNG	���~�U�q/)���2AJG�-=��$���̙��&�@y6LS��b,Q@���u~^������J�'�I���d����˝w�*'N.��|#�v���Q�_|�#����7��4���߲
��嗎}����W?���yM}ۇ�ʵk7��s���s�Kg��|��d�&���z�6l�'����B�]@��H� "�*�*EH����q?GȘ/�m͋&Z����hhV�����5��A��QP�A4v)d+"��u`�$N���O�gey�n&S��A���$�)���Ǡ���S;T"@BB0���#�J=��� U�q\�#\�rXc@��bH0��s�iدg���-��2ݲ/J�!c�+��&r�z��~@����~U���^�����,�+��ss�G���N�S�N(��ʫgd��-,���'ʩ��(ͪ��	����LVV�2�E�E1��%�#HsȂ'�Q@�oxΐEXO��GL�ca�r�kH̤�}��LTYCPT%��hc�{�Ae�m�SE� P�?�<��Q�xZ=ϴ�w�� q ���1N*j�|6�\9�u#�������Dؿ����%>b ��N�Xb�՘^�ˠ�id�裄�D��6xz�M�iP�:�{�Xi�M����}߱;U��
��ਬo��!1+�/%�.̖��C�������S[��K_|׻���=��O<w���e�׿�̷��~���v�GGGs^�.M���gʕ�7���2�HO�i����
�%f`���'F-�Q@�^l* �H5A4t�@oZD�q&�7�����o����9D<"0l�����9/B)T�x,��+=�{tV]�Xj��,8��~p�Y�+����������f���2�&^� �� Ϩ7���?��¸JGY�5iU���z]��t�{D���cY2���$�k�Rϳ����]u��1���C%i�9����s���h�y��{-&{�ҥ���^^���}�����(>D~�Àzi����Vn.��G���=O=U6���0\`�ɋ�ޜ��!{ @�<�
��\%O�_&�U̮�˵�|��b���g֧��2��x�v�t��]}�eʽ���z�~jM�Ju��N`c +������Y7B���C#J��X��̔���1�^н�W�B�Q�)=�T
U׶���ek����)���tm�3��X���V QB��WOo3�����7
�ϞV�c�+e��\�%�wP�����I�QB�o�����U��M��T��{�?�_y���u.6�����?����{�,�sK*�����O|�_}�굫���<��B��������ҋ��U��l���P��LK �7�Z	�CSw�L��"eVI(�oR@�[W(+K^-���η����Y�����N�\s�
�#�m��)�n�o��h3:hi� �#BO��DKX7���^{�5�9.���R�$��:�P����Ʋ��
��8��gb<0�<˦p���<Àc����c��mmj2���MP��ĒC��M����'&�����?ކ�uyҥ�w�}�m�i޾�A����gr���ϖU�p��K���x'f����-ex��������ē�%&�b��H�y�m/-���! X�H�
�uBG�0�k��D���a Þ���P2[�V<���7Z��<�(t���K���ZgG��a�V3�̙�Pi(D�OE�V��Q@("�^Z��UF p�^���yO)�}�ʭ"k��XTꫩ�=�j�	�?�l9J�TR���9�$9Wq���2=9�8s�ز��xc�L�(!ŕ��{�U�%J����N�����Y�H�*��ӧ�K!���ږ�����ܓO��o���?��[�P�-���}�So��'�����v�� �A��r����g��`��`��SQ���"���]K�(�2R�&��F�y@	�V$J�@!R�ٷa0�۩�<je���������MJ���Ԉk��� 1�T�FPRa���W�Y��]f+�����K�*#��Y�{Rt��.���Rk�����F'�.�������Y���4֒��T�#!m�l�J"V�\Xg���B�:��2��MnHUڂ[-�e���8��BN1����@����������/|��-}�+_��h�TUb|��Ϲ����w��	ZAw���NYX<F?�R�G�#�=��B�#&!(h]�X��t��G
j ����|�<7�0,�̢�c��Dꂃ�&3�{Ce��V�(S�Y+�.��_;���6�A����Z�M�_�/PЙJSϩ!�����<qjj7���Kc-�C�\���01k��%η�I��Ʀ�ѐ= bK|%+�ƾ�8U4 ����|���ň!��}C|�	�utx�̪I�{@���Ao(M�b�"Bec��{q�&���'����S'��DϩS�Ծ>� ��}v||��}���>�����2�n9D�������_��CC��.GC�p�=wQL.�(N���@�\Y��;f)� ���]AIЅ�9�b�;���h�u�$���fB��ɺ�>a�m�ϱc'�B�����OJp�Ŷ����?�(�[���
�[ny�,y�P`{����M y�.p[�f��27����j���#�(���X��'�l��gh3�^���.�B��W�����8a���Ay�ٜ̹�t~�i۵t�[G0v��Ą���o/O2�"=���c���%�o\�"f�n�8>��g�k�/���f٥�(�J�c���(sӣe~a�,�����r�����)�{�&����U���"O� �n�I<b��Ъs_yV<Cbr�	s���j:s������\�5����5�,@{F���w�q	�{�Q.���w�5��PO��}ŋ3�D���Ѐ%��e�gf�¨P)�I���{&Q���_!��_( ��X�Tg�a q�)(NF�R@*U!3Z`�qXaq�	#&Jh��V(���d�>�[P{:I"����H�.������kmA����7o^׸E|8�W���S����߯B���t��X[[���~�����}��v�h�:�[N}��g��o��/�g��\�UGɴ���ƍ���ū�ᄩ�f[��N��'M1%���Xނ��M[�;��Z1D%d�+B�`��F��`���(
&BTVZ��<\P
�NO��H�LZ$���G�X���(�;�扅��w��p�WV�H�Z����6j����?
Jb��{���9�!���H۶�    IDATc�ŕ��������0�|��9��bĘ�h��)��U�0�oMx)1�g���I�db ��7ʸ0�zq�ZOM�����;�T�"bg�7oX@U:�|���3e��B�2~�s�=w��q�"�3Eo����\y�����[�V����*�vmJV=d7j 9m�V�q������J��g�3F��V~M`�x�mCƌ��$��<� 5@ʿ�/��c(��l��1��86�J$7JYB��0\�{j"�M�gl7��1�=(���j:�:�H.�G�?��i���u^ۙ�J�����M�>c1PDHp0�Tk8��ȏ�z�4��g,(.�ȩ&����c(yH�b�婕ϫ�ދ-�����b�3^�y�C5פ2����Y�+^�=���уN�����w������Zu�[J���6�[���?v�ڵ����>�"����9,7��ʅ�W���7���:��V��B�d�bU��<6,��P(ˎ���
�����¢���SQ@�LI�X��P���=�^�i��#�6i,����3�t&�wp��c�����.@�Pb(�;ɥ������e��/���?��BomnhSYZfc�Xǂ{����|�Jæ��~�t05�^�M/W�8���'Hf�P���=ӱ1�����\Ý��XL+v/��B��.�i���e�\�ʈ�7 �k�I��+K�ʍ�N��6;mAq�?����j2�=��;�n��թ_��2Y��7ʻ��{ʣ�}�P�`֠�<���rBd�1)�I�8�dRQT PǶ̐��b�݄��q,@�鹍��h�Z�[������>yU�#ʍ��g���I��T��ë�kb��뗲T��+܃���1ɃjBƐ!a�mE���:�xR|�8�Y��
�æ�A���_�@���� O�����d��
n8ׇR=3Sxh����̮�Y1բ��{���"s|~�M���^�&H�
���T�����|��~��j`z�Խ����������'���o�J^�-����������?�:�S���I��V�\���rYY]L��EppX)��� �^k7 �ŦO�Q\W��G���`T�*d�tj[d� Î��r5����*A3N�r��Z�ZUT(���Z��V��BK�]�s᷼�ξ?,̛K�{A�Xd�5&V7���2ā%I����ٰ( Ci��\-����ppy�)�جP��'���)�I�B��v|�o�8�k��Y6O���xC�7�Ɯ�CY��n�G]���;�쀷��͸����7Tjgmu�l���au�,/��+�6>)�x�}�K`-//�!�h/�2>1�+O��=J�<q�d:Ҽ�2=!� �F�p���sP�P��6�h+p	���V���ߚ��S�	)&9B��ojrFFP��S��8�����g��(S5���㱧�)J��u�qx�&CP[.�X���x�3 ��N�����]M`�Z��z( +y�_�`�h)4�E)D��<��P?�e�v��k�o���4��}Ղ�E:B����}�����������QD�xb|��2�VLF���*�-Hú{�{�������<��#������ɓ'��x�n��:�+��w_�r���[o�R� ��~���m���+W�����(���n�&W��#^p.0�,3S�Fȍ4���XQ�,9����q��ԯt=�ys�v\��ּ���R�e>Y"�Ŗ�R��xe�����*+���uZ.l�r��)�Pi͉Ǥ3f� o����md�ŐALŠT��EHm��ͅ�%�@�{贮�9�eH��㉛��sp$+;� � �^P�P�P٘|��d/��E�&Q0�g`<��-!C�f��r�`Q4�����NkKɈ����8u�0h�lԍ�k�,���+�.��+Keww�;~R�uh*����\Z��.���d۱QC��cY%�L<	}^;�фX/G�*sAH��h��8�H��(]7�0�/�����DMX�rTO���ya�TꩵS� �d�фZȓ*�����ҥ_T:��;����a��=��X9v���E�!n(��&r[1��V��^*�+ި~R��u?�Ն�=�~�x0d�������:a���Qڳ�9qj�E)$�� �����Í(ޡ���WRT@Y�� �e���i)Arj�?'O�(<x�B�i1����n)����}�������-�{�o���?��m����������CC��XV��~�~}Y
hy+tO�.7��0c�TVs�P�<dɏ�i���PS,,�oV@���U�y�N���XS)Љg`�Ʊ����wF?Z�a)��W��{c�l>,�`�X��� ����b��~��g3#(B���2�3H;w�2C���^)
Gc54�BB� �,P]�?U�-�������Ӫ�a:�P#�+�TT>l8�����$�^lA.��*��(h|`�T<��{!� ����������,�,K7�I���6��tvfF\Pᶋ���/�-��[es{�l�\���L�ΗK7������*��6�sM�nm�k� ��Z�)�ޕ��p�+P���#���"�2*�N�\)`]�7�%��anz�g)s�W|���8F��jĩ�0$�ڇ*���j�ɜ�a���ܸq�F+$�l�Ee�A��##e����`�AV�Y8����e(��N�с�[���~1i��-��
�{��ӶH�8R�'c����m'��ҿ'{jc�2D|-����Y���=:���7�>�o U>wU�~�,Ў�~�I0ܽ��-Î�_��յ����C���K�l4:̯[Bu�ݡ���_�ί?��_X]^�����i�{l����r���r��M����|X�ѷ�8)����R�
�Dg�(	��m�����ܠJ.�L�P	�8�HU��2U0��i+���>����؉^l��y��#0�z3Ff6q�,D����b��y����s�xK�4w~����Xd���'���?ظ<�Z*������޲�}<��9�ł���|4	����j�	8�[f�͠Wh�˱3Ɯ؃XO��=��C�֜3�F�̱�W�Zy(�Ak~}e���Q��ޔ'�|�zY]^.�v�_X��^�V�e||Bׄ����.��2���H�'O����}��/�A:i��Q�0ǘ�Yc.ؙ8R�@�ژO��v�E�q�����=�!r<���'k���b�D�Ȁ�ۗ�f[�׎eXp�Ҟ�M5�l����B��P� �b�R�Mc۳�)Ȳ���Z�SjGº��ٟR$�Ӣ���^�w���Ȅt���F)���9����?��*��٫��R<��������G���a*#�& #��'�m)��Ad��XU��]��t����L�BR�5����k�pw���P�w�qGy�#)nҍ�#1_�u�/������CoqQ�?��-���^�z�W�?���������,nj9!,i6w���r���rx4��>�0�mt��<a�G��a���W��!'���������.;�6�^���X����2��K	L��{� �s@�RI��à˂�5���'��
��ի��`���}�DW��'�,H�e��I����h�R�X��ڶ�%$L�؛��f!.��H!T[��{�q�	��p �PPA 65�5g�l N	ʁv����sIQ�+k�g�9=>��M$0�W�R�S����ofr/h�ܸvEI2ă�^�ҫ�W�osD����2F zf�^9f)���[�Hk�j�{�R�q������X��wE��<Ӱ�S
�
Lڰ�Џ���`�cdnnA�ۛ�¡V>�^�A�{L�Z�����:�R�	�ێI�X�i�$��0�״[���[�ϙ��o.9V�z@��HP�"��3cýUH|o��q	W�x�B�vրi�F�g(�
[S3ӪjN�:2�5�S		�;�B��jK�{C�e��KG!8v�!]]���q��0�,Q���7
(^k<��z=�jR���u��n���u�*��}��{�ч��w߭����b�l߸�􅷾�-������By�[B}����Ͽ�w�[?4::���E��ɲ��*.\)���j9R�����kw����Kc�*�Z��S9,c������@� �n��r���8*[�ۂ����D6<%4���
Rc������D����]qy��L \��#h�%���F��t��%�����;�BpS�]
hl��� Ӵ{�r��s.����Q��[�p'��1A���b�i�����:=،1ONM(�BH���[�{��a~Ef���l6H$�}$�k�>~℔ FB`GƇ��9(ѱ2��p;=�d}s[��"8���W��V0����j���G?��Ʊ25;�g�`�8���w�)@�'����QB�'\�O(����ٓq3>�|D�����G�$�\Y�̹�!��s=<è���t�(�e�L��ͱ�Z�=�`�h77�'�#!|���a�y!�U�������U:�~ ��-��9��B��3JA�I���b9v|��gc�x��e��H��j��]7�c�2P�779�����:�޳��+S����ey��:�혢�Q�߁��,0�A�)�7�	�D�5�bB��'Tݯ��2?�ԁ~	$���Ƶ��S'�i�>��}�M�RXƭ���F�Bi4��~�����?�"��
�۽:�K���?x�ҕ��h4�cjzr� (����y�\�p�Rj�IG{
hddBm��{լ�{s'�(A1�H.}m86X5�!�͙M��j9%~�*�H!�{R�Q������͉����m�bu�ʪ�X��3NY�5�����-0�x?����q�L���Q0Wv�r_��E
N�n��4�TXKl&+�Q-쩙�g���ǁ��\[0f�܇Xj5��AnxbR^P����ac�g�{1����<=3�h��J4޴N�M|@1Q��}F������	⫍ؠ_�l��zU@X\�z�+�Sʔp)���r�}��{�%�Տ��bX-F�O飬���6W�	�n���)�8.��6Uu#π9�g����q?�@S�7���r��e\�m�v�t�L���,�������&�C���y���8����N�u�@<0���/�X�Hx4��*Auy=߱a)y�>0�����yo�צ�[Zg5�WD�B�T\T���c>��9�IC��T3��?���)On�`W݈���mӅfT��,�����c���;��Y��f̯��A�v��RO��QYY��^c���b?��R럵���햍���O���'���~���a��z�/����o�\����f�yZu��ȷ�W'ϳ�.����22L&sSA;�%�c�������0z��	��MG�PE�i"Dm��
��j����֟��\�M��U�hΆw��!s���p7\�o����Z�@�ZQBasi ����q!��9���q©�.T�k�����9�80N�c�,�,Y Ծ��e2s��t@f�,C6F<6��+q+T�wdn��9��`9����?�Q��	
(�dޏ��`�ޡk��B�a��<�xyu���u���p��lImm�� ��W�Ց�_�iZ��#����xn{!�|ϧo;)t���a��!��G��lv����1Y"�d���}�WK.�����+\:�ح�{�V@�6ֆ�ў�*���'�X���#\��ƫ����G�l�\��!\�zY�䡇�W,b|bD���s%v��C�}��S^0~���+%��Ѿ�H��;r���4����GZ��'�ƽ����7"�M	�l����J������ֺ�=���u�Fim�ޜ������ڭb���_xA�lR�ego'ΉamφDP�(��~��D��u^��-e{�Un�X�!������Q����}o@���x�=������7��5;��v�9u�s���ݭ�u�$ґ� ��,� dc��0da0F�����2�+�B !"	����( -�R��y�|j<U��y�SU�ş}���:�S����o{���>���z�ѣ/َ|y!~��
h4�~���W>��Ͻun~�+vww��,l>�3�����c17���	����]q�)��b��M6L\PP�P��j+ދ�2�+h���=�\�.�ȩD˹&��r����<�X�k`���c�l�e��r²��ɍ%�k�J���� l �-���Z���$�9�kؙ���(�k5a�{@��B9t�0�f�ߡ�ƥ�,|�6��3���Tc5�-�@1�Ir%k𬹿���c�Jy:F��������k	����n�llm��-�c������) �#���kbD=�Z����/zѽ����q� �ʺ�z�	�ôR��5c�s�0��lyq.+o'�Bz�1t��Js����U5�Z�hK
�
�X�Qⶶ!(8Q��6}�{�����=�Wʍ������r�ʥr��-e��{��e�����:�������o�o�U�\��p��ù��-E2p?#�<-W�sKjCa�3�ٱ)+�x4i���T���T;���j>�3��<9���Dӧ�]��Z��s`8��8pP��0��1V#
Ȳg�r�Y �ȥx@��b����՞fk��f�6d�<q��8~���e������5_���K��U^œk��
��է��������_|p}}�,��iќ9{�\�|�\�pY��"���ȑ����k�������e�#�VR�# HP��V�J����x���u��M?�L��jyiM̨�ɉ	��p�s	����<b���|i%�l[,������a�X���<Yƣ�$���O �BP_�s� .�M ��D�[c�&E.Q�a�ɓi�HaLS_��"��� Q0�؀%#�<*���nc��c�Zt�2�s���q��s�3�|(j^�e�׬s�q��r������;��IH2N�#�t
,�W�h(,�S�N��ǏIP�S3IK�
�kЖ��X�7�ڸ�J3����3��=2��V̺��sLQ��Z�-�2�-B���^���u�vFy26���ND�ef��@�d$2O�x���e��ѻʉ�G�m�s��oWkygӞO<��OBS�c%��X�C)փ��(�# ��Ż�Ǯ�Vc`�#�����x��4���3Rm3�������@	�nQ�J)�ĳK-;�5�/'��7����j���������T	�۷5�<_��^�MF�y�69bo{f���}�K_����oz#���_����>��?��?���F��7�Ctk��	�>��J����@���¼�0�hZe\\�\݉e�^�Pl�-P6�~h��$T�t�( ���
*�	��j""<�&[XU���	=Vp4֮��R.O��T�����������l���:.i���ඤ��ʰ	�����$r����6Zv���KiqQ�&�4�M+��0=�����b�U��j�)�m�+���P����3yN!�@�μ�c�(�d��ge��d(�ĥ���Z��}r�lm���*��a�<�`9u�x��y7kl�cYs~Z�JM<��Q0�n�3�Z��,��Q:i9"X��	�x��(5�Y�K�x7)�K	`8��/��@K��K�)�E\�p8/
=�>t��e�׷\!���n{cÆu�6���W��)C�(�`(-��`j	�U�gש�_���})�G�_Qm�ĩ��Qr����@�3�m?9C�ާ�o��*cJ���T���f5NF$P�+� Ԡ#�����v���4����k�
(k!P�R1k�z����B�c~�hGcz�Mə�~�<u\^��t�r�9��9t��������˩S�o� ��2����SO=5��O��W�?{步1|���^��Z({�A�X�.�{�ɲ��#&	荅���GV��	�b"�<����5؋�;�,�z���a�<H�7���b6�, ����aiU��s�v�qT�UO0��
�A��i�(V~,P�1�5̖X��X|ƴ�M-F����\��pg�<����g�Rb%��M��Iq b�    IDAT@�4��"�Wכ1����i��(V2aq�-U�!*�T��>�jl.�b6�Ҝ��=��keU�J����t߹�[�9)�k�2��r�I[���\=-�p�ȡ����V'��͵�7��0nL�0�/k�v�e@��b,\U=�b��s�M�B�W�l�,,��-��k���a�e|i�aC�a����޸��zk��r���cgaq3��+׮	���sߣ��N�UC���;?��1W]pu�b�g�<����k*HD�R��WRg�7x�X���c���d]�MY%2�!^b�����S	��)��g�f�)�?(s-%XG	i��S��K�3p��&�ɘ��x��ŗ���n�;�(�	���zQ%�k��\m�����_RN�>�N�2lG�+������z���|�[_��>���>��Ї���߾�湹��[ZZ-W��.;��r���r��aoX2�a�A<��8��kW΅yCoQ8( ����X�q�#��yA8��� z����qP�����!���s�	���9��b�G8X�%��y*_,lcp���zJ�>X9,*6Ft6M��JJ���2�͞P��(2~>��?/W�\��Nb���`��7
)B3Vy,����[J�T�x�W���1|2�k*�V��/N����`�7^�o�'�0��B��b��g���Te�w��z�[y.#bF ` *0�wM<�Z�Yr>����o��E�-<1^�W��e��o�G�ssNg����;9����e��9+N�M~�׃+2$���?x���-�}nN��X��h����&�,�,)�
�Qr���h��BWFر����<ў�H����~���dnnݾ�9��9Fp0�h�y�I+3Z{�j�Q�֤*��)U��V������=|�.�e��c�zuޕ�"�O� 	A�f�c�=�3D��qi�
�VB@�)�A[-���g�Vծ��ȅ1ZCک2R�T�APۥ�+��8ǂ&J���a��c��|��y+����C����V:�i�>ܹ}��_>����گy����^o�����)�|�]/��O��/�z{_7�1Gf��v�<���r��U=�t,5�9[��ᜳ�e���D�t�`�$ٕI6V���x�Ͼ�x@fm��V�9���8�w�X�,h�\4�9q�X�^�!y����x�m��}gq��fa��h���$�$\#1�T(HB)�ye�$QwUh�|/S)���Cіg�sd�/�!X�A�<2��.�1_l 6X}���OXX+����g�5!D��\UŢSL{r�J�ga.σ�1#
hZ�G�ċC3�(�.qj�1~8�a�J�Wzn�#�(}M�V�&?@����`0���M�X��<��1�q�b�Y%(� 2!�g���q�ԈC�B90w�hҼX�oCN&<���ۑU� Fxs�\+q��ex^�(V�e�[�a�J�|�re�:D�bgwS���X(7o�*g�|AL�x�~�j�=?�5أ�ª�)���Q�-:oO#�O���b`���W8��z�1V�J���7M�Q{�Yyx�~��2ا�-�N�۵�����/ԧg�o�8�k*)���y�iE�<J��V0T��Y�x�0:7c��>u�����EF�A10u��wv��������/yɣ��gݣ˽ 
����+�������6t��#��A�\��!t��-	9�,L�,��r�Ǌc����T�$
H��JQ<c����d�
��lm-�V-VZ!"pZP����ؒum�@�@,Yr�����dsy3�~�j�`�,YP�����������;�0jc����8�o��(^���O�3g���dlޔ4>J�~'QQ%LZ��U��#1��UV�����WːXbA��i�'3�Wb�(���%����HԶv?�QN�7�c�5p5	P
a0���ߌ�0��xX�;{�m�Y���W�
�T��P�Ki�MzKY�nܯF������Y'Q��VZnaK�prbT|?���#�h��#Ǚ�5ʵP���R5j�Z�2	��sLR0��E᠀ҟJ�b����T�zP�3�Ey/z>}�^ټMQ\�	�����[�ek��ʹ�6ϊ��<I�3�44���=b���s�8%��\'��e/�
�=Ck�w{]ׅKE�ž#�Xę
�e�.ϼ�l����3w@Z�0�lp�H��̺q|:h���-�B*�RD�Y��e
+�(�w�B�|SM��Ԏ�ƭ1	F������+9z�e���Y໲���������g�������Q@O<��>��?�o7�7��tOJ�Η��^9{�R9�r��ީ94��َ9�����ģ�jQU��qͭ( �	ZT5�mX�Z׭��dq�}��e^�i�+v�Y��v
�������OZ/Di����۰p��F��x?�o�Et��sf�bJ��j	E����v����/-�Nݣ��J΃]�"����ӗ�hc\O�j��t�F�a܂'��l&Q,6Y�C��J����	��#�{�Y���gyU0�*����(Q�>{��Q �@X���<��^?�$'V���s���V%F�@��*9.!��,Ar�5�qE]���Pd��{� `%��ēN_$ϣ��76���g�:Jr)�5�4��̵D<	ك��xu�N��g� ���z��d���FĂRϝZ�l�{?�yN�,��Ѝ�X�D ژ�ࡄN C�*	�[���S%ʄ�ͱI���hC�W����rE	b?Rеܐ��,��T��ҡ��!���vL�d��[<3:�Ż����cbO�	��(��J�F�K��vw\e�gr�[5X��[#'���Gʁ5R\܆2Ű��p4����_}��_=z�y�	zA<�~��_����/��请��eY��Y1�>����Xp�{Ii0�%�sRб2ހ�pj�dY�M�7Q0>�@���r&�@��Y!v�x���idW�At~ب��"��>�!�X�ܒp���'ǲ������G��n��cKq3�g7���P�l\P�޻�W��"�>.긼P7gK���nlt�]�0��h1��XR�`J�a��UhT�����<�xp��,�$XZ��s�X�3Е�W5�w<y;<i��
ʕc�$b\��l�����{s��wم�
��@�R�m�*N����߆m������d�/�b�ݶA���"
��Z���p|���vv��6�>���l�sb<nD�+���2{�������rE(��=֏�VǏWfݾ��z�񀺥�v�\�����Q���v�e��c2���-TRQݷZõ�BM"�S�k��9VóF��84�w�^�y"/�����#�D{q��Q�̼=��a�0߷n�0�V�:��F�����S��1��C��]�^w����K_��� N�ʴ�p�c����f�exu���{��#M����(4Ku�ƍ��������o}!r��wt����|��}�ų��Q���2J[@����+7�O>Un�o+v"�X%<�U�	D�E#�����tGS1 �K���GOo�"���Q4f]�V�� :HqU8%
����3�U����9_�RM��c�dCI�U���M�K4-���Z�5�;�X�j�dK�D��Z���0k���
[,̋*�7��%[�����3�����&��XL9E�1��:V��	 3~	�����xO���0V�Ł�@E�c��i6Ppp��(��
;��]ȓ{�_c� i<,*>s=<�#='*�e�ֺ��gՂ}��-�ٞ�M����&,�A��0)�����������4���n��+�0/O�qr�I�Z��6ַ���8~J���U��~���<�=�Z!�V��1��whO��{�2D�ϕ�^*l�H����v����6��/.@���0A�� �9�-%��\Y�
���=�Tep֚w�
T�U�3�\�Ҽ��֪��?G d�ˮ��22RQk)��y��iߵ�J��3����8Ko����YX^W�9�##r���$�y�ֽ���qq�x=Yφ�ȳr�7I�a�m�o)��ڦ�	m20�y�Cj!?�$5��C������[�7>�_�?�������6���=�
����{Ϗ���~{����NO��p��^�TΝ;��s��u�4.�"��~*<�Bm�#f\~�X�ԓDZ�^��WU@`������R��	5����B�k�յ�(�2��E�,P����d�SV�zs
hzC���~��b�����Ƣ��?�����T[T(��z��Z/��h�pO��I9����b&&��^^���U���Hc�7;U�u��.p�	�\��on��s��9�"��}�c�H�ѣǫ8�u��&#��*h_��/�J*7X͔Ƭ�|`�q?��M\i���}�%��fJo�VL��[�'���XVkRYÞ��V�����RJ��+�S=��|޳��ă���.�8��X�0��>7w 2�)�����B��yq���*uWL��J��6�j#��2�b�6�u�$,k�Վ�����:�z,�iV�!4�ӢD�'�Q�^7��TA��H!A\�<x�ϋ�����sy��q��z�
=F<zƲq��-�LϽ�'�}���6I�Z���'��=6�0�eؤ:�8�k�CQ�g���i�#��V�U�������~+�eG}�ӧ.��:X��.�J��ٙE��<y�������m�����s���z��{���G?������p�53��R
��l�us�<sx�k���.4yZU_����ǃ�"kF
����}x��ȨN��R@`�( S}����O�`1���-+��R¡[ALZJ��
����uVo����|P�͒J��6�rL&jm�}Yݽ��]mU>4�I���x�=r�	yu�r迆ߎ;"K�x�O���FIՆ{�m�PV�Qpm��l)��S�XD,�$�ɦԃ7��ǰS���[Hb#�+�m<P{�fE�9nC����啸���.x���y�}��^����DU��<A���Q�̫Ղ!1s�-S����Ev}ou=Ԏ����8Ob���䣸�٤m���ZN*���jӞc�:�}+B�2
v�4�Նf�b��2�m���O��6E���o
7c�9��AICR\�6�ڽ?�7�¢U���ޡ#go�ƭ�k�8%z����%$y6�2��>��P�<w�Yg��$)�ZK.�
��9�is|C
ʕ&ġ��{�8!����[b���P���ީ��}3��1��E�D���9��~}�B�DVD��^�U�@�j�P���"S�`����%����W�x�(����Ӎ�ٙ�z��}�?y�k^s�y�=�+���F��k�����_l�����htZ���F�t�jy��g�cE�$BM��Z*�N]+��Z��7��d��y
��f�����h̭jUz��.�[�-���A�o.���5��I�7p0g�,EA5p�%����Z	[l�J��󁡆�$��fq6����mWV���G�� q1c
��g�e�a�[��3�*0Zk`1�iJt�Y�V���=8<��@!�\+�1�����PQ�w�)K�G�-��`N�'粷iEŜ�`����=׺Ch��yggKpY \�v��ē�j�����^�9�؆�\�}o5K����r��.��sA���U<rҼo\j�V^��O,k��B%�C�i�&��s��+��a�(:��`؎�K�3�+��[M+�5]�"����V��Z��k�A�ג��ˍ�(	�j�E��LQ{枽�>�e�O,�,U�~(uD;���,J�9H�oyц`����
<��7��ǽp�u���#�}���l��IBq�5����5�H�Z����'�����_�]���$Uӆ���r\xWQ�x@A5�w�W���k�Z&�5c��"(} TXQ(���&)��"
hyi�<��呇�Ә�
�� h��7����G��ѷ~��ן=�:�yU@�����y����vw��u�Q���mcNx�ŋ���+��[n�-��j5a�ЙRpO-��"ʆԴO��F�V��X�T�MpWV� &�)�v��7��u��������!,f�tx�J;��"����R�e^%?h���� j�I��8�~��q�S�4���k�ϻmK�f�^�q9��J�59AU�gP�"E��X0��a��l�f�P�(BJV� 
2��I�a��M��:��U!�5b틥T�pN6uXV�-HTă5	���[��A᲌P�iɁ3�1#EQ�}bK�>���g��1�X:,$�u�X[�>�;^X���w'�,��:��`pE��`G�3��**�4�R�13�aPƓ�p��i���d�k�,h'�r��)d�i�9���XG-��]
����3 �,����8h��9��O-�J��{�`��Ȋ'�'C�V� �b�VU���-J��_��_^�����|�D�(�_Z���ҕ�S�
s��d�t]�I���^Y\���S������g�;��	�\r��+ce<TQ�Æ�?#况lhT��(�a�x1�aC˨��ƶ�r���&5(��9u��]�ŏ<T���愺���}����ů��o~�#�<b��yx=�
�����/�ԧ��6��"�G��B�z�F9w����v��JRV�D�'N�C\߈M���Z!7
���iH��w��|�֯	`X�V�3๳���$�*�C�y[f��ǒ��e���|~O���k�ɚ���X#��j�]�c��Rc�zn���@H�>�6z��
\�x�t\(��k_IQ�>���
%T`�����'��*�=��Uzx�%ץGL��{�'ٰp+�U�f1rP$/F��ĕ���]��y��J�|*�j ���7�S� ?IA�x�I��(8��Κ	������,�[JgM���gV+<�~�{�r舡�P�ܦ��ُB�3�j_������3%��]&���,���3�);ۮ��XG9����L�G�x	^����=\<�S1� �q'��䓟�<�H�moI����[�{�9�!/�ە�0����\�i���F��/8�+_�J)C�V�5�W�|��t^TYa�^�r����r'���Tɰnj��U+w1Cډ�j<y�P%�9\]^�Ƙk,B�3+^�e��U!��s�LW�(�g��0�<, 81|�Ϊ�}���r�ڕ*K��L�C���/~��8qL����j�ӽ�����ox÷�򣏾�yKJ}�Ѕ�����k׮���Ly�p8lJ���r���r��m2UD��x8y,x@�eA+s~^
(7S�J+���	$d�Wb��x��2�]�^(AH��*��YԚWae�e����|G�G�YV$�����-��Ԝ������m�F�<��c
%׈��e��Xo0�f�O25��0?���#آD&�ҾcA5���( [��+���L VR��
@m5��w�<
.�P�>C���2/<�ĉ���z����B���?|��F�O��r=bv���R��Z��p%��M��+\Ι�ᚁ��S;/�F{���@n��!�<4A!q����-��j��?�Њ�,�uY�Y��=+�c�Nrl�yp��g�T�O���kӹ ��-����%�7��u{ccL��bOB�o��k���+`p��Y{�1PL���⧔��D�3��Wy㺉?=������3"�X��k�1�t�U�xwGƮ�g���ʯ�Xd�Մ�$��.(k�H�mHr�
g�'2��S�z9�'+ ���q��FI��7y�/]��@���=����Қq��Z��������z������7���U��_ϛz��O���{������n��A��5�3�|A
H%�k�r�m��y��A)���r��m�x��3lf{A,Y��T�E�
ێ��73�gญ[������?J� �Q���t��C'gA�#*trƇb��{�w����� J�`ey��c;��߲Ql�Z�u�>�A��t�@
Kt��#&
��LCP�KN�e�(�(�l�2�Xɺ�,�T���TŌ�q�\a���<����YQ������5���)��Y��0jb��l�|x>I�<�fk�0�oz�|N������{�\��&2�    IDATߊ��~���P^Z[��z��ū��˼+��i�(�\�H,���[x��c.��^!�x�QF�&d!���87τsMWw�=G!��X�|v%����K�� c��6�Hy9��:�c�a����
����U3�BP?��/H
�����Du�P�/����s�Kq�O�؜�ى!��B��%C��z3���m�� ����(�u�*��i����K^`������g���K�T�� 6@ɿ��Yb�Z�=S�w�.ͳ��J.6������5�U���Wz���Z{y���W?���~�K~⫾����e/{���;�z��?�އ{������뷶n�u���._x�\�t��j����0Y(���>�u��V�C��������%kr����ʾ�~��� ��Աw�~94�r?>���7g���p�	�=��6�C&zI�V�$��a(ڈ�a,Z0��:.�Ǥ�
��k��\z&�+`�8���%f�x
�'O���U9��D9�����BT�?��Ը��ʝ��C�e�|�<��z
__[+�{����K� 'W9���o6r�g6md����
�1'���r�����%��-Q�9o����K`�<ދ�,�Ե��X����v�U�����A�@p�^X��e}4I��hˈ��;��3FQ�w�j�{qb@���'�4�ň���^�ʇ�@,��mQ��($,ld�#Ϋ��F��T�~1���DyV����A/nX�.��-��Y�~�P��@x��5�sP �3�x��Y�:n+��;��ƺj±G��:�8Ӱ%ľ�w]?�d�����A�~�19�N�F|Ƌq���EL�%���Ɩ	)��q���:�=�C=X��uX�:�p-�����lk~�}�w~���җ����=:��F����7���z�s�]�Y^��t���+Wo���!�$I1��| ,�z���Y� ix���E	�r��� �9�Ɇ��q�\���=l�(~���z��l��R�V�E���.�B4t�,fY�6�2��f�<���YU5�"� LnL0�X����'��=���!���P�L^Y��"���/����g65ղ�pY�S����z^��(�GB�o*0?Q~|α�'��/P��Tˆx+]uQ�QR���U�IDQq����N8�b��\3��<�[�<��(�@����_gL�0�v��i�VJ�����P@"Tt��U+9�v��1�"�9?1�*�:.c��L��i��쎷�F ���Fg�)��-@�>L�1˓h��xn귭�f�<QB\�[��I���8��1o���a�\*˕/x�9X�mX���7b�q�o���W���r�#ǎ�=�@��G�zp��O�&�P�#�ͷ���7J���g��ɵ:m7�6d>�ոԕϣ��@�Y�g ��*��-?�7�U
�t !+�S�������p晧��
�����_�ѽ��e� T��F{��~�w�������y���(�?����/\:��ss�G,Ha�Q��R�~��8q
� ��H�����F�M8��ō��.�4�&�6���c ����g���E�"�&�[TG�-[#^ 괪<׉k=m9��eC��Bۛ���apE�f�E���"%U+2Ļ� t��8a<���!%V����򳐳�%����bD�s����j�4] 3����U�?)�j5s�ľ?�b�R�"�dc�z����F�eDiң�P �x�!I8LAq�
�	ղB\+�a�5�c��m�
�֭�c4��R��1�NPxj1��>�D���������&�	��qt�Y�'�1�%�b����9g*H1/͗����EU��#��-!�K�3�90�%ϣ1��Rǥ�4�h�㣜8�p�P�f<k��Az:���DX��s�:�1P��@�@��+�\p8�����N���R,��[r���]M��%��|�0Ce���Zv<;�*ʕ�����56�깓w���TmoWH����@j�(�r�����?�<���o����;��G��+��'�뻾�3���{�{?������W�t���]ތ���/��i-T�,���w�������U:��er��Oڴ��k�R8��d��J�ł��&ã�e3i�k!���<�
�lf	hߜ�QBl4m�������SKiH)�k+�UcV�{�qm,6��@{�x����Qh�v���R7c�F��1V��ꙓ����"���w"�"B%���|:���?� w�(��=���	��yC�^��յ�%ج2ׁ��YL�W�S�,�;�Y�`�c�rҪ9B�S�
�(�v�1��e��C�k��}.[�( ����XB}v187�ǳ������;�'�֖KM�&��<�xH<0��.�%*��V\��<t�{��m�%��<�5#�ȊtIL�c<2�����k��+e,VĎg��9�?k��Tj���Źbگ�3O�+s@-���9��3&Ρ�2e}���N��#xt~�=����w�ew{RAE����J=@�g���Z�MǄ���ˁ��S�k���P�S0�i�H�[~3/Ġ-+\/Ň1���t�=��*/=}ZE��]B�,��^����ş����w��.9r_ϋ����e������p�u�����iQ+7�_���J��}�zYLX�g��|��(�I��+l*&,8{��œbA��΂��%�k�*Y]s�Ei�Y{`�Xb��Jb�v�R�H��ʞ7��N�)Hі}��[`<@l�x|'����(0`0|�����k.Cb@��	��#;���@w��p\�-�f,m�9]2�D��\�(�t`$�Ch�?�9Cp"RX4c�@��l�m��~",[�X�z��x.Q�^S.fI%�x���.! �ur��b��b�o�-�h*��u���K*L{t�����(�:5Tb���A���W�����*�
v7ݺE$
r%XP�fc���mT�5���%�Q�z\�cjn���eD5�6���e8VE���o�b=��`����8pl�ܢ<s�qksG�&^����؛�a4빟�������$�<O��{ܓR1*kOh�� Y�<	�RJ���9A$�"�)�A��+���gϬE����(f)��U���}9�MI�$˓�=���sm���2��
���t���/���D��~X���s���Q�y~gw��������x��;�{t�;��Μ9��=�'_�����F�<��4��`��*�<}�t{�Fȱ�V��D�>�(�<�YP<�X�$SF�J�ԍ�!�,xA\{{ǹ6J��mr��mI��I����/3������hI�b�����+P���~GծQ<fθJ�%� lx�Q��s 5d"K]��xRx�;x6�V�}k9z�C81�x^�<ᆀ@�p�`�Q QB��C���ׄ�O J��M�+1*>��3�3Mq����s�i�r��kG��d2���9IC@�R�|�Z���E�%c�*5_����V@�G�Wr\���z`��9Wjo�g������s|:k��xj,w�Sf�'����Q�*bJ���p�@S�;�����y2/����QʁյjP�~�a~Әx�Q�\������$��/%��~ .�-]	O+f)���+���ƺ�@ԑ��iQ:��@��xK�`�d�}���uj�j¹=H�r��+9M{�X�{}�K߷���Em[�F��D�6c|��G5j0��,��f\j*ϟX�)�6��D��fd��Bd�q��'����ɮ֋P�Q�����o��7����Ƴ��+�˟��]���w��ׯ_�{���>0�X�t=�p���O�@WU��Ç��Ynd������.��=�5�F��>0�-Ŷd%�~���.��`j�R�x8w��D�+V��ڂW�G�	���*X�а@�L$�ʪ��~dq�k�Y�q,�E�E�dRu���?]���X�c�����0��q�Q[�V~�8	�ʒ+�y�5"���7�˥����Hq�����*����+�:�c�f�]j��(�X�!�JL�@Qla�q���5�c8e�Mb3w<V��J��fj���3�:q�0{��Z�`����ި�e�3�k�8g,~���k��Y$�-�Q֚���V�u�1�"6��ժ)3���!(��}Ce���?�*Ef���@��9�< �NwKr<�6�����8��R
��=��\�!�AS C�ňP��aMv�s5�x�T�HNX/f�ΫTN�<�no��l�>�Qy�E�d䢀����Z�"�fPH��x��O�uV�#�Fe��8�M�U�f?�+#{��{GΈ�#��-b��������l���,���7�������>��?��?�ؿ�
�������?x[�����ht
��`�=wI,8J���eCc�?vL
(T�@J�H�@�4hk�4��l(g��|x�EIb)��ֵ|K�ސa0CR�~bQX+̻�=�RG%��

@~�~�4� x1���^j%"���� ��=�{#C��b�'M�8fڪ���(�L>
#�V��_=ƚ�m Λ1��@����2_�,y�(!��R�JO��Z�(֨����'A�ڨ%�3�A���R@|�3dbl|҄@U�#
;ߛ��(�x�(�@f��sR!�{w=�I�&[	�dmN
(�$�,�U�{q,�������E�ū͚�0��po�p��a�7s����^.g$��5	���Ë����塀ρ�%��GȘ�����d���jO�^����y���� L$��5�g'�o4�QY^��1�W,,�[�yk��	�2�+	Gz��"�͠mH���t��23kc���xh��M��V��Y�~_�5�b�e�z?�"�3��V��7У�q�.c���ԅ#��f�����G�Ï<X���!���b���>K������s?��w�:u�����Cp�}������_i�6^ݜi.�u��zy��3ecs���l9�G���G���w��0���Q2�t�8j<%_��V	μ� 	L���C�5|d(�E�W�a�j�������f��3E�[��6�5@�y�H�����6#���� ���`>PԱJ�M$�B"Q��IYW�����ЊWA�58^ɀ�|�s[t�<Qnx-�f�Z(���8.0���N��p|��\����>J]��p-C�Ÿf�;��8CsF�Vr��a��C?{������5[BXe8�Tx���x	Fǒ��>.�O<�io���S�̊he�-�/�Gm�)�9o%/��3'�p{Tq�YVj��^`;{+.���N�<3�(�(��s<sRxy6n.�C�2h�|$��o�1���-�5��ȳ:�|�hS���:�c�����v��;�������i%Xu[D�6Z)�iSlk�/��Z�#��AXk2f*�DJ��"s3ՠ]ei~gG�а�&�n�BaPɷ�`h����kP�ݬ%�f�TQ�A��֡�[k�����B�8mc�{�:|��1R))lL=���������㣏>z�����*�х����{���'��Gò�
A����7˙����F�tq�j�:���)>*��o�k:ǅ�d����z��DC:ӏq�y�r�D��o��M�i���F!����z� ��(�\��=_�Da�;w��GJ@e�&�*�� 0&��fHp;?tj� �ڙ��>D�Y�.�8�|%�c,�x���C�p]�G� �D�0e٥�}��+-Jϩ�8HM�B�4J$0f�#����b����
=Sj.*mz:�o���E�� U��kڛ�@����%��Q���yL�-#㍂�!"h�O%�-c��k��πL�2�J�|=�J�ē8G�X3v�cf�q|bmxYkQނ��䳘�������DR����s��~�ŀà|,Oc}]ϐ:���i����T�0�Itq�o Vs,���s��,ϊ�0.����S~.(��G�`���Վ�5}�~U��sw:JX�5�7�0�fp#�����+� �̰,�͋��q��E�����s-�q�T�9]��>���>���k���H5rɎ
݅�#.^1c!;$����r���2?�R�-yd.�{�K��ƿ�m��7�鎶g��
�ʕ�������?������v�m�ZT���k����es�[��7k��k��
��c$�`��4�$��J6{VLnpr���^�j�b�2�&��C�0�y��( 6V�\���C�w]�A�m؈<^H�S���AΏ����gΪ�S6O�D����*(���w��x{��4|�����yD�����V��Zf�� �k��(t<g����Hy�����7$dhK�c��8גe=�lq�!b�:]N��%63-�9O�/��`���:mr�Q��E�����[�t�z�7Tdp:QWVd�U0�@o�B%�R�����#���>c�x�I�j��X��l`��{X���|�=�d�Y�yM��g�ָV�_kK�S���PX�i U�J}A��
�L��d�T��㌡��YY��;׵���@��-) �0f���ƖbO�����8Rv�%#%68�͍c@���ǥ���li���n��a��m���3��ćPR��H��tfQ�K_r�?��(�>ރ�����D�*ԛ�oT5�k\N�y�'�.��EȵbHݸv������S��C��W�Z���[2N2�vw�:����?��?�鱕~���
�g>����������vw#�Uƾ�+_8{�\�t����zJ�80Tj��{�=euiY�������،�<vW��ZJ�}x8��yhX��C@�`�Y�YPI�7����9��$/�VN����Ư�X&��vzb�`��C��_R����f!��S¾�nf����j#�x?,R�&l�i&�HS�A����ř^�q�'���yluz�YX�C��0�y�9G|?q�X�|��(9��]���=qe�7�-�h{����U��+���qn)��i�*uYuH�8{��<�r1^2^����0�r8�_�O������|�G�	[�":��V��FqU�U0��{�f�Y�� )9&�E�V9n�ƹ��ch�*�Ԓybno޸Q���%X���R�+�#�����k%�nJ9��Hp�Z8�r�����IJ{BY��g��A�^�N�&{���rb���oh��Z(�n_%pBJ��;��L�	
����Y�Ѣ��~h,�I�e�HN<�>^2F�\���˨����.D�� �x.$_Fx�Ff��^���ʺ�[ǎy3�(��(�ª�����~bJOQ�1\M(�Q 8��q�_�$2�c�>u��~�!1�Ő��(
�(�O-����[��=ￓu����G�s���{��[s3_�i�����-�������ϔ�7�K�OF��iؽn9u���"H$�k��,�$�F��0q��0c��	��>�)Ǒ�;m��r^Z����<(�#���z��/������rli4���q\�0�ŋ�yؐ&ԸQ^�h���ne�o�JJ�XtqG,�%���x��|�}T!�+�M�|Ʋ�/a����ɱ(�(�f{������DJ>�8�I�6=2��:�w�<��\/�u��}�HC1bJ��@%ݬ���l`&�`P~���ؘX%R^��*����33�|��:��������A���@4�x*]ʾM(��l���p,_<A�U�F`I9ap��*1��!]?����n���!q��_[;dO�V^N=4�� c�o�K.�4�'����w�}��e��k-�n|��ܰ�כֿu�#Z�˨5ji ���Bg��:,�T�����s���Q�{��E���S(��E	r�(b��SUc���y�k��m�nk��װ��3 8
��8�ߵq�v��KĞ���.�ߜW������֢�7d���#�[/�v��"C��ٳ�S�{�С����)�[P*fk"���l��?|���;^����}�˱;u��h�x�;~�5O|�o��m>���M��nn�/|�\���]:@lkɑ{O�>�Q_��	�MD���!hq�Gٯq �s�TT��n�x�d"����ۏ�	���
�Lbmġi��b��Vٜq�ϟ?[�z�m|\u�����f��4�gԤ�檧�N�    IDAT��j�g�Tf��i����G�Y�9��,q��S,Y6�/��LO)�jY{�����B/k��#(cy���<O��\��o�+'ƃ�
&���e�gᒹӲ�Db"�C��^_}PP$(0��o����b�4���j��H�X<`}�`Jr�((����R#���9H�T�0U��a�($�K�2�9� �4
��+�̆6�h_��h��wwvvǂ��<�vX9-��+�!�=5�b���M̸EWR�<�f�u��@�1Lr�F"j;�Z9��������Y0�aeb*y��ڕ	z��q~�M�i��5Ys�H�D	�t��5����f���X0Q��{�#����޻Y�;������-�~[�J)ն�G�ld�]��Ү\MY+��\�Ed���T��\�p}_�1L��� ��uʹs��̓���@X(�O?R���t��D�`��\m�f����㯼�o�c����u�ց�/���;�?X��!���3j��Wn�s�.���v��m��
�`��������"*LZb������0�$�H�K��\�	F�N� ��W8��E�����
�`���s*�j�F�H���=�e1_�|Q0����Vd��;�9��BȌ��Y�)($�͝����Ԣ$d�U���ě%������P �O�{�~ͬF \C�ǭ�-�Cx����Ą�9ED�7��9�=f�9c$^��a��4���@�p�n�s�� Reh��ݞH/( 6�N{OJjq��U��a�� ���濼�؋`Йf�S�z��Bs����}d�K�VRB���G�5�9}�y)����˚�#�AX�"l#�'M�:$A�P���l��8�8T�s�~����86����WF��G�J!�x_>g�|~O{�V�n+%��m�D�S4ĝ}����a���8��񺞃�m1����҂dU PF�l+5;k���;|�\��1��H��jL�x����b�tFU��N[
��v�䃚-DL|�w<o��9+ H�t�����"(���9�խ*�����y�3'@�̕1uh�Gy��}�I3��J>�@7�����W��g���~��;��1t��gO�����ϴfk0蝠DB��+���k���+ew�WF@�ҐP���m��Q+sO�)��h���B�
�־Q��o�����j\w赜A�9��DV��8�L
�3B��8e��,|�$��d˛7�kD���&W؅��~�/	+6Ag��j5(�c�=9%|�s�;��e��\X�ɤgsL[t��9a��]���9���X�S�&�2wy����Șt�1�/8�j��ל�Lw���?9N�IwK�����5� Ci6��[�gī�Ƙ�G
��iw�q z!j�0FHn%i�1���g�>
H
\~��k�@��7-X��RVY�ָ���%�ůxZMH��آ!6����O^��k�v2r�UQa��v�n�]م�^��P��	d�j��D[��b;��n�1Ż�ђrL!y���P{�:�,��s�P@ɥ� ��M�J6
��B.����8&%4h9�/��Q����>��E]�����,ϔR<Rt]E���b+�9���<�n��m0���8荺����������MJA��^��w%�?r�0~u��I]�����"�#�1���v�����~�?��	�wL}��~�w~�wy�Y^�����^9�r�r�* ��/�v���z�&��Ury���S[Dg�B�4Vl����%�VD��7�D:����&�CY�{�)��Ǔ��r��;���gb`Ѫ��ΎX1�,l��p1�g!�Q�i�Z&C�*�S�a�-�=$���H��Q�6P��!0pK���c�Z���Yln	���6l@�+�X\�9��&ev��Da2��@?����}�(p�d�ӕ��Аlg˴z�}L\ a�
���T�>c@է�ଡZb@�Wש�ǫ�k�YZ3A�( ��i��Y�,enV�!�GyX������s���}WV1�+����9Ф��yci'��c�%�1@o����k�ޥ����5p�������SN��V�`��p)�'����@bQ,�=9���&�� �
�
f�jj��I�}^�<��,�đK2��,Ϲ3�(�x�( dF�ѣGT��<�i�g�5�>j��5��g��YpKtb@Y�%yss3���o�)/�*����"��h�B8���Bk�Vk��~�+�fVF+�����׈�`d��y���^�
�D���z@�� L�<�9����9y������Cx�R����{�+>���x���u�����Ɗ��ؑ�q�v��Geva����iëyԑ#���5�r~N ����P��,�!{ɘ6�U�;�]y@��]c�s(�˴�����,L��X�|/�1F��Z��"�e�Z������e�s�a�h#�n6��\�U�d�Kf>E`�
���y�jm��e؀�v�XkӶ4�Ҧl��a�1�[��شl>�KI�E�f���ww1幇D��j�g�Q�+3��1��'�(τ�aL�*,�V���� ��FS��ŕU�(b"P(�Rhx����īr�4v�w o�4��3�=��7�4/)���8ȑC�Ǭ�(P�B,��O����(����-/��k�y�lcFB����bTvb"yFa�I�W���m��l˳B	9��D,�
(���g7-�e�7l��0��^����Q.��+2�v�����9�����l$F�AR�Y�ϲ�9ƹ}�es�z9|䠪$���F�$�������Y��l��;j����{2`vv7Kw��P�AWqF�vxF�8�j�D�AQ��kܩe4��:^�cQ@AP��أ��c� �Ⱖ�S�����SaRB4�����Ϭ,���w|�㕯|���B~��#
����K�z�;����??S���U݂�]ʍ����KescW�nsn�l���e�j���S �@��쑈�Z�
�-0��Kӊ�"̕]U@P�Ě����<K�+XK��-E�岃��ѱ0b�Ǫ�Z��������H��ax��k�A����5���p��΂�-r�S'�6����q[ ���s$H�<0s�=Be���0q�>A�oMN|��#���b�r��M�³ 2�oFsXZ����N<"��֦j�F�	�_ӕ��Q@��}3��ǣx$��R@�O�h�^�~H����� ��賂�/ʇ=7;N`�+)���3�4��n`�;��Ʒ�,����
쒎�a6E�1�|D�uΝ����߁:����م]�g��m7�È��#ܙ�x��'M�@���8��+�^�2����GP����˒��/R.�ޔ(��eԕ��58&���� Z(�Y��'��]\j�~w���r��b��=�ƪ�����TV��*�ԭlNP*>p��/FL���;�*���Xd����:�W3Ǉ���
'�\��S;eV�NrB�GmD�?�ठj>sv��5y��9�XVa�#G��aOb�tڽk�f���-���׽�uw��pG�ŋ���o���v�ڏ4��i���2��˗�K��PE�U���RlD�o�������K�s-�)��I����������e8��`�/׷������TL�f�L+�	�ֹGr�eY�� ���g�<�/9�,q~�(��L�Tc��/�M�c랼�����jBR©&��E����D�l���d��T�QM�I��&9so�ݭ��b�G�r]64�=�/��歴�X\��k�Y�o�1��x�z�6�#AT��|G�k�c+��]5$5��T�7 �-B�&n�r�k�c��	ށ3�U!����������5��������Fc\u�J�o K<��x��~#g�����t��GP���S��3�̫����O���2��p�~S3q<�쳰+�	�9�����Ϻ��Yl��̲>�u�?�R��FX��ẘب���X�ǲ�Z�1�<g�E^lkҶD�	jq��a�,-ϩPi �<�x�Y��;� ��1t��g�t���x��C�Gm�ĥ\�ΎRBJ�?��G\��;�v�oV@ AY+�
��̼��(�(`<ݳP�8��^>c�y��>�Sc�X��+(�1��a��~�w�����x�k�Mo��;R�(��~��'����nܸ����� ��% ϝ�T.]���hG���N���y@�$"p*�� p��%����]�>�ެ|�ɓ�d����t�%�iaԚmX챸Y��(*J.P� )�e������X|q�m"���L_��X8F��zzt�X2����A�@���C1nm��g����#P#�i��Bp`(��x#^J�yV<�B%l�TF4��ǜ�Cm����V�N,��CA��ك�����a~%	�M��'���X�t�y'�`_��y���Z'��#�ô�&08d�j^���!�]Ō�(D؞5�� h�͖F˱�(� ���K�Qe�c��q�$�F�L<"�8�a��]	�a�l�o��Օ1	"���O�P6���,8�%
�gb��:��2ߩNd�s1��x�\7	�Y�̴Ђ�o3_�����=��%a�Əb�vl���ʐ�<���o�t̒1h�7L"���mΌ��#����ZC����r_Y�2���� ��)U��~�oR	�3q&����[:��b��Ȏ!����lp �����8?'��<F�]CpkmN
"�C�>:�J�-�.�8?�$�f�r���@� "`��s�r��q�Ejj�x�h4��u�|�W}���w��Y����;��>��O��������q�o�6˚,)�-���K��嫥��h�E�v>z�.)��*��%8Z�l��S�iQ4C��"�U�Iw�đ�/�җ�<b���ś^?����A�Xc}@�`QǪD�ZM[���b�ŊҢ�t�|/�x(Zd�+�[����g�*��g]�ŞOm�;3�>'�>��X��6c�����H�+��3/l����3��C��(�X��Ǝ����-96f�!VzbG�ω5-��*��(�@u���J3�95��j8/��`���<�
���=<h�]m�҆�6��W喔�f+d{f��G����+%&�$s��y��-�I��r,q�1�ŸA����\H4��q�4�s,���Ճ��V�<���z��,rMy啰���햗u^)���ޕ�]�oz^��8���blQ�����
O�z�U�96�|M�^��g��?
(б�{����e�$5�?蔓��noW�-2��|�^s����ZN��p��&(w*�=ja�ɾ���R@0Q2`3v[y��K���jY"��	B²3�HB,y@�]Vz�m��A
���+�}�ƪ��f�q��/a�����S�N��*�������z�N�?z�K��e?�C?��x.O�uGЇ?��|����;;ۯ��m.ɚ�=��|�p����鐖��~9q���*HI�bᡀb�O{@�3-�	�1'F�d�e4Fes�=�I�j �9ppM��s�&��~��i�൱�d�'X�$��C�mR��L(��jГ�٩U��ֹ� ��P"*�p�!�0��< ��2I����Y��q?)��5�D�ٓ����+<�D�w{��v�q�a�!�qlF�?�zPi����b�$�	��EU�9>�΅���8��
�K���7��V����PD���H)���A���$��P�X!��ABHU Z.�3V@5aKñ(��:
��޺^��x�
7�~V������/k�1C+�( ������Q�c{����xᨖNRY�����g~��w=m����{<S��a/#��&�;�˜eN�.uL�@qD�e�bĠx@&]ζ�&���X���Q@��̻�{�fs�G�r�಄4/�@1���0s�u�E�*�U)�YI�q�(�^�������QB��H�r�����/�eei��4r%#y@����h�F�>P)�T��Q�p�쵷J�vQ�n���W.]�Rvȝ��V��K^��
���亭b�;;;��`����~�o�w���(�sGл��ۏ>�����^���V�1+13[��v˙3���k�������I\'���ZH�N�5J[pf� ا]�( S�cY��4�'1���s�f�n����8/%uظ( 64�IxU�,<�i�O5溰E�Ebk/�������ʦ��2�Y��+��4�!�uL��?��Y][Ӽl޺����*1�A|-g�d���)�(����j��q��l6~��i('�*
�Jx�l�l��H��;b��2]=[���-��t��`>�s���h�����2`���jm5,�I�~�i4+�_+TRA��x|R4,����{\O& ;0�Y3��V�3�K��( P���t���RBu.��eaW��2F�alAN&�dm	��h�����WYfZ��
�k�k��@��u���(��2���9����cl0��L؟�ùV<u�+㮶��|�����>?�{��2���c��2P�����^�,/��>(�( U�*��c`�������a���xCPg�V��\O��]
�Δ�>e����֦�bRb�P�wZ��Օr����oLڭ
\���Mƕ�h4SF}�%�<T���l��}
>;zg�S.^�Rnol;9�Кa��w?q��j�C�T
�1�=��0�/~�G~�7z�!���s��h����}�k��3��R���2x�zQK��V9{�b�uk��4D�4�E@��i36�}Ge����H�Θ!�EN�6P��;��(�>��kR�r}Z�57��@��1�N��}9�
�#�)�k����%�D8[�3�����<��V!�����Q�˵�-���� ��G`Q:\ӊ�I��,�%��}�Ԧ_�[�s$���Q�H�4t�=G`�g$�T�|�8)��y� �p�c|���{�.�á3)pK���No�Y{�
fw{R@ؐ@�`���@1��];�f��C�R<��6�4��륆��E�$�E�qQ��㢓���Q%�T�mD������̱������6(x@<�%�J���d}EɄ�C!k��B>IQ�Ύ�c�`b�Ns"�W%JG�x�lP��B|��Y��]^a����be�)~*��Sk��[���sq�8���4O���2�+������x���jH!'Wbk(�̨(�D�Юs�H���q�ϑ{�R�V����H&���:l@�7�{_TŎfi죀eد�����:}����)�._/�o��P�
 ̗�ww9y�H���"�"�m�_��������;��9W@�Ν;������̙/�X���
H��JSe�Ϟ�\��pK���3X�!E �UK�M�t��d8F0v�����h������m��-*��cPg���ܿd�e�-B�I�R6�5�3�x��V-4�l1����R">�M�	(��g�ū�T�u����y		�s]Y��s*���wW��b��p-�-����t[�$���Ë�p��[��K!g�֙-O^�h����5�M���?I�Q^���e�w���s�pP� U8�����CGx�Pg���%ŀa���듴�RF@��HB�B�|O�Ő�P�ّw�WU��X�V<V:���
c �8Ƌ�Rmh8Y���bTQj*ʊ�e�ēc�2�t�)��%�A�����ѕ8�Xe�Ͳ~��Ǚ��X�W^c��<^1�<�A�ڌsbPLj8F�H1WĹ��+�Z�'�#����k����w���Z�5#6�J��V���X'5Ն@����5�X��T�z�>1�05�a�1�\����E�ya�#6i!]�^g��	�~�$�.--�+K���RX�
s�
���~�!5��(R�߫��>�»�?����h �W��/W��,W�R�g�9q�RN�}��s�	��Ѐv����v�������������:?6<��>���'>�G����׮_��>�.kxXT����+�K���Ù����X�9u�[�8�"K~fbUق��H)���q�'�)�m��-�a�y�"	rnYP���A\����V�Q\}Á5v 	!�1Xm�m�s~�ڒ��D���QX"/��|�v��    IDAT|*��E����D�=K�`�W�[b,�1\��(�Ă,�@K�E���� � ��<(���ͦ�܉p�>I�mVy��8p�G�t+�U��ā�4�xQ,���b�З*\W*�^{NT���"&	uq�,,��*l� ����Y��"@��&)�jL��LP׹���]	��$�^���``:NÎQ>��P@Q
�t�
�C���()�ϹyKʩ6rK�[�͋sJ�F�D�J�RZ57-�&�~P�$+E�&�Ɠ�gkxu� )@ֿ����,�CLnZ�%�Ź�_���dl���[Y{�%�;��Ӽ��\�s�f�ɏ�&��m䰎)ѓ\���߁��q�+�Ĉ�s�B�VrL$j
�H�-4b�4[�}�
hqq��./�򺛄�G���d���q�R{�a��ۥ�߫
�k4ʵ�˅K�
F84J�ԩ����)��ʨܼu�uw����k��o��w���=�9W@0�>�������7v{탨]65�.��RΟ�\��Q��1����,��/z�&��O����r��Q!���U<�( m���K��ϚR�w�U�����oss�en�\^n�m���������9�Z��9>"�����뷮��N��޼]�7�Z;�!�$)�~g��*�W-�/���/��J���}�-������ ֦�k=��� aN����\'���w�C��%v���g E�ᡇ��:��ʵ�'��>5���1ߪ�����=5���C�0lb|?8�'��덭My@�ԍ���#XCu�T̩�^1�$�7��A`-_ᨱ�?��,o��c�Sŧ(}�u\��6J��2/��s�������U�Ј�Ըs�Տ��G�9sŽM�$�>Wf���[����/��҉Y�Hm�����j|-��4Y�{L+u�4Ǆ��X�>̵�ɤp���=��yT!ZBR��xO5���>�W�V�C�/�I�6�L��Vb�5�N�Y��
���x���g�,5�=q�([�w�Xpy�T(^����As@3�j���}`��aF&�ke��4�96P0zX��Ƥ+9ȁ��ʛb�"�î��v{���!2ܸ�QΜ�`d�/�X$��~P�"fg���~_��no𡗿��~��~�Ǟx���\}�#8��?��_�u��_o�Z�r��B��ܹ�칋�Mh���YxC�?z�dq��ʪa1 �pbEn
���j�,<[;Cߣ/���& ���Bk-h� $�^���ie���R!�)8���P̌��j9�8�lo��ݭ���V�V��B�K����-�Ɯpk�S���YXgi�����0L6:�M����p�Ac���$�	���X$T���x��ɓc��J�1�-�3c��X���p,��{i�����2�6��}w�S +�U����jp�B���-b` `R�O5Bm�^e���X��7n�k�	�����%��ñG'��G��2�U2�K�8/�1��P��/'.�I�`L'!Y��0Z���kk��{DA��zg�j"p���5q��}�s兑$(�V��8�U��yց��w<����mI��Ŵ�b��}�9.���"cb#ώ�1gi��}�9 ��\S	C����y70?�c��x�����'�AEE�1FPgR#S�/Ϥc
7犗)�t8�zc߷Z��}\ge����8��6�&ygi�f����u�TF�zJ�p���L��E�<Px��Bi(����m�5;��t��;u�O��/����_��>�������G�����W�Z���Dϵ�xz���r��U�� ��f(�r�ır�Xg��A �5H����}~� b!�*�Ŏ��]�`���B�!�q��ȴ�i��H���
����Ò�,\p����'롌���:1-$,X���V8��R�&�*0ZˁDh&/'��@DQ�QбR��W�R����!B�1r��8�l�a+w:v�u��Qt���}����b������IY6
��b�iW<)�(�8��)WR3�+�e,�(o&�.-Y�\_&sժ�����)�h�;�Y��� �p<�f)��i&K�ƫpc<_(X�r���i�B�T[�{]��(��c��Pk�A�ye�
~�l�g��+���"V��Q	�T�J�g����>R���s�=�=��P�*�@���)�,��$�a�#F[Yv(���o����C��N�����5y�%6�6��X�Y�Œ�<yz�7FT2&��������j�'����g�ǰ�M�Z�z抽t�v�q�Иj2�TL���{����9�;	�ZO*dc�=~�	�gw�"��v�pd(���,�2����i4�~����啷�����?��#�>G����	��������'{����_k�ZpT5i�~C]�~KP �/q��(w�}�9��M��Ƀd��N�V@��,0"`9u�k�n6��[!<�/
���HWB�ܰ�l	[9�HX��D5�^l䜈��-Y<|8����Ŷo���D�e�l�T�B����++��j�x����������9�׏�k�@�3�����g}�y���/�V��5�f#��<b�Ƌ���#l�8��B^��@6���1XH �FX�-<,B,�����]{U�rk�[ޛ�3����������謨��f�<�[��]~�Ƶ2��s����.�on֟ߙ7χ������5ᴉ��o�~�,�Y�	�H�TI�^�5xI��BȺ�*�L��
�j J㥓ei��A���)\	$ID�r+���{���P2����W|R�	oe����R�"��/7T=���7s��k
�ca�P�����+-�@��֢�@�Vh�,�.�([Q:X_�M��ю�/�k�U�s.Ŧ1h�%��BYLU���9���^Q�N���X[����9�
A�%,%�m0��5� �AϨD�B�&���>��}f�y"J�s[�Y{T�@�4�b�%�����KôhY��Rܚ�z+��)��X��4�݂��g8+e{^!�u����'t8zm	�cG�����LƧ7��~�����K_�Ҙ�w�u��ǖ~���+?�?��í��+ӵ�v纫�nGT"FL����C'O� �&�wЊ���!Z�Es�3�H4^	���b��hM}�cZb-�%ϩUZY�1rMJ��b��J�<o���~R�ḓ(A4u���l��3Lh)��p(��ZA��|n���
�u��E��Z0���E;��w�����W[��@�<׃� �\g4�!�E�����O-
c&D�u�r��-��>|?�,��"��5��<�\���Z�'S�z-,�W�͸��H�����j������N-�0,�Z�j�Hu���x��ǜVk�����3�Z@-�-��-���cTJR�rXC�wyu��C&WTZ��O0�kJ�Ӎ�90n֛�|���C+I�� �?
]��B���*�ڪ{�tDI����u]�k���#A<**�����_'�nV��(R���(�|����֖�+�amma�\Td<?@�"
�@��g@M��\ =�:!8��J��&uދ.�UVհ��[e�3�Ӡ���ܠQR\���芳q���BR�#�i�p��RB��-��y0���~�}�����vU�*�.]������k?���}����KX$j0�hW���=�ԙn��F	 �3�ç*d�i�)f�+\�'�d6[�Y��A=���}WF˲�y �?L�k@#M[�$r_�q��ދ�lżv��"n�o�BKS!��b���F�VA �hPY9��:��U@(b�V�P�'D��"�(���za�bT��˸]K�~91�6��Z�Q-'��ԚѲ1��l�h�}?ϊ H	^ٛt�"�t|����>���sn��wa\{�1:F��ڃV�\��5���@Ţ��,\�;)eO)��*�cݗ|4��p�+W.��9�e�����!��[K���	-�Z��e�a"Y��_J��:Ӥ��ؠМ+�W��Y6�`l!��o��1��=��*D���ܚ�7�3�����Ԭ̽�J�������
�A�ϰU�7��(�ueI䃵���+%K��8�<)$k.�	`o9�):�$1�Z@P@�%�>���*�R]}f���m
����nW�����(!�f#�
�F0V@DcU�_�d9���,�#���Z���wv��
<�s���Toa��,��^�Y�ɭ���`0.�ߺ������o{ի^u�I���
��7N�������?��wv��CaL������W�'O��nҡ=q�D���Ų��A[�&��<8���o�&�W4�@����H�T��!D#c�&����!��W�4�V���a��蹃����q��q����,!:��̵(l!���0�7b�T>�j���5�"`�h
f�0Xt�h�
m�A1�V.G��p������K +�cMѮ��^���%���w"䃅�}dv�'�A�B@�:�B�5��Bοo��\� ��s8
�S9�G��8�ˍ�k������Ș�;�__�>msX(��iU�x�[���9a�����a���e�E�B-fӜɬL���ܻ��f3M��ϺkY��hA2�Ǻ4�+�SMh�dw-��<g*;E��������I�FĿ�(� �U
�\Q���A��,����ٰG����}�!cע�^YO���T��e����܋����iqQ��$=�rO�"�37�PY�ʎ���UR�k/Sq�#�����3_P��f�P�/�/tB��~�X���/_�X�rځ�e�#�>T59�h+߂N��quk��ӯz�W���_�?�նwU ]���?����ֳg��[���

�G�0�`]�x�L����<{��PZm_���t���=�-���C�[nN4��
 	�����p��8���t@r�ڔ����c�-*���8��|�JklO����0�f)=t�vw�ҥB��.�J����-�	*�y6�2LrƎ��3�z�RV�)��MeQ=��R�|ӸKp-Ŀ�K�5�aQ؊�*贒��3�~��@#u�
�0�Ya���p�ܫz����U�(95��.��h�%�9�%�~e��5&���o�1��'��l���&��˒'Z@�<�vpqX��혐_�H�bD-���P��t.�┨�-/J8Z�A+U˕`�m�0��%�2���HQ���936�|�����F2�i9���h�D���� �.��[A}�GzCX������1н4��[,��>�����	�RXp_#�Or�w��
�o-2~��Q2�sQ�E�c���,n�0'�QH�p�X�A��G;��@������$��H�řdmJ��,v�^�q�/����4M$JF��|�V Q���|����"��;ׯ_5D~}o���~�|߷}�w>�W.>��� z�?������7\�p�5ˋK�J�]A���Ϝ�|�L���[��yֱC�ρ���D �����B�\	���`��2�h��Ւ���ߵ88ߕY'h����B�Xr��{�}�W���
n_>��}%t�VRK��b�"��`��L@p% �gZcu�X@��U�\b�Sa[�+d"$�5h��t��OBƆ�]UZd��g��H���V?��,9���î=����(��C�����V��j�<S($[�&��-P�����>}�M&��P�0%\xVY�i-@��h�s�D��C�Y��y�#�΁����a	Ֆ������ۜ�f��G�+L��3Q(TV[���$kZ/}(��cOX����n4s3���0.�Z#MHf��R_��M�����=�s]��Z�[�s�(���e���^�+ S�M��� 0��
Yh���s 6E� 	-.�>{�₠�:^��3�܁����r�@ &��]aA��?FAa����VRF��Q&ȃD �{	�B�p�X��Gn���;��u�/S���`*�@����g�O��<�N���_�F��,.�Z6E�Ψ�{ߣ�>�o~�?��g*t�߿������w�ܿ���.����CLlq�,�qw����ǟJ�jUƍfv��#U���ʷo=p��%KTĉǂ��jS	P�ǹ��
-&��#L8�Z�8pA-$V�	瞐V� .fLBR�����Jp�'����>Ć�>e9����3&aa%�6X���=��oC8�y|��P�����UK@g���^�j�o�a�q�gݧ�Z	�Q�t�:�u�<�:��Fa�}AE��Dܻ�h��� c^k�ZW0�>�c>�}p"(�sc.�+�&����W��g2v ��~�a���!��j����TBu�D��V1�CG�ԁ�Q4��#su}���KJ���2�Y�� �SkP��u�"���]f�|WG:뼱9���|�џ�	
��/��v�ky-�W�G�@H����d�̱oŚ؊��T-��y��z��w8׮ş�-�}���s��+��̹�QHfјl7c~g<Z�VHQ8q�-��i�ƇS���:�2a��ìX`:�Y{N0
�tT����Sf�'�f��G����#u�?��P���N@	�}�Q<(A2,��X���h��b�z�d�U	L�noko2��C��}���;~�y+������������������/������ݧ�J�T�� D� ���>J�9��8!�,lyt�lJ�gi��ܿZ\_ ���B�P��Y�����rH�Z,
����oĜP0Q�`ZՑ!�.V��p�45�`�i=�AD�,�U(A�|Tb�cj�TB+d4���yq��_��k]5e��2�׿҇]����gBH ��!��_�<`�̿B�[�nA?�W��L4VQERD���(���1M������q/-��u�w���U��G����t`@�j�U��[-_�B��ܹsu> hd�̗V�$�1���	P8L��̫,�&����= ��t�k��O�����Y��R��|yN	8���2NZ���jd�`�y��)���,�0d���ߑf�`�O�����D>���b�v�ʑ��g0>�X�n��x�B~Ф%����)�$a��],��/WW���=���Zw��0V���-͍K �g�O�,&Їk@y?�U�iÔ�G��JD>YY���F�iA�f�:@���D��*�^i�ȼ]4�R<w��?~�;�����[B?������������������y+�����ڋ�ϟ�mlm}� ��B=z�&y�����'��ZI���!��{O+��Do��80%�XO��0x��H�,����2������K%���B2jA���1����^�����l5��_i^;��G��,��a�!�l�ص��㕊�-(�C\ɯ�_M	��zZK�^�uY�|�a��k���
d-�r�6,j���AX����>a�>`L��5R�/��jq�
=i1���{��r�y����x6���\K���c���k��R$h���~��Ƞ�U�:�oKKt�#<��_@.���p^j���}������R����V�N� ������]3�Af���Z�υ���L3���� �+$�D�L���QRL� �Ç�~�#�glX'ZfB���` �*H��	HY��Gl��O�ž*(���>A�U�/-�U<�\��ItO��0~�� �ί��5��DLt^�6��k��7~E�Y����ZE�)���*�xśSK(tԊ���9 3���U�*A��ٳg�]K)cx����l�7�z���dw<�����7��u���苾hVW�3�Fw����>�Yx��~x8~���[z;q���֭���g�uO>����xj���￷e��
��'�&a"j���);#��=W �����܂����\a⁖Ԁd���E�o�G��si��-w�YbXxŰv�F����j�����9@2P\��bl?�ѿ�H�P�������Z�է���A]3��*���i�O�;}.BL\��E�����<��5�� ��bUtXK�f4m��O�U/)ҤRs��Y�� �֦�{���[��?�D).�?�x����T��c��z�!�� ٟX��@W��w_%U:Os~��&t�*�x�!PVa[s��ȱ�f5�ʒY����Q�(FU�Dz�m    IDAT��X4]w3�SBa�w�r�r�'k]�{+b�9R�R�B
 �Fx�=b<*'Ы~>�pƉN��j��r�_Y��٬gp�dDO
�3�Rr��b _��_�ⶇ�Q2���:
Ǖ�>�B �/0A <h���� *�UQ�����{U:�RRu���)���4��SA�緆t�J���It��I�Ԗ��ًbx�5Aɺy;
�ȑ�F"°I�-�����G�_y������ˏ>�h�x���
�_��/�7��_���p��s�E�������@���J Yr呇N֤'c6&�:HM��R��=����
_尅�b����7�¾�$� �0�����T�T�,��, K��*���*�e��s1^Z�������d�B0|]���ھŧ�� �i����2y���Uf����kX�$���3v��PX� ��O�먜��|7��DH�7KV��ޒ����ZU`h��gs_-K~
-����X/�o���t���'j���G)�z�K^�y.��u��~�N7h僸�]�ai�����%�A	�_�AӨ�x�B5�����[���x��n�V�B�,�Lk�\���O�h>wm��X�jQz�؅��ɤ�!�s-�h�I��ߨ�u1�
�Y�+ i}A4v���a��	��m%wǳ/�����TL��E��`�2�����u�?{���X��<G(��}aE��������Y5�=+��,����GT��n@<���P�/�Z�J�#p򊢃/H�,{Ӗ)-�EF*���B	4��������c�_��h4����w��K������ƻ�����?���?�������������nU%��/t���i)�����{�9N㕂0x�cA|~*�$EK�+�v�S�]48"V��l��=��ܷD ��B4	m�ϸ'H�S�C(�-¿��Ӳ�������)����,L�h$�e�3��P 	���Z�tZL�~6�S�v�I�|��?��ʀ�P\i���kŌ���&�=�E�g�[8���
������ߵ��9�(�.ü����
oMk�Y��c�:~������ZR��̦���R��~�S����>Zs���;q��
��EW_�����3)xY�ѫ�G4�>*��:�`]Ǹ���O�nVzM㓈_��W󮹵 Sxu�(�͝0���JSA��
��i��X����c�B����:�=>�`�A`��SRdV�6
d�1�#O��{`�>�)�(�� �3��'��*�$���O
4;Cӌ�N��� �GD �w�����Rֱ�h��h��(�E�"Ԙ#�y���(8�L8@ �7J���Xу�<y�=v85�@Q@G�[΢i	N�83�ͽq�"BE@��̙3ݵ��ϗ;����%���-U�Z, ��&s���?�����~�K��Kn��S����=���/�Ї>�n4����`������ƭ���s����h��<���ssݣ�NvG�.E�E��R��0�P��E�� �zFM A(.<߂�e���)�.Ȥi*�'tU��Pg�3@�����P��3�#��(��A�y�b�Ֆ�5rG녟0�Ҥ޿/BU'.>$;c�Cs����=ĮW�scJB#P�Eo��
� ��Yߗ��Ӗ�-�J˴��Z;B<��%:>�;�%i}ijM�wԘ�cג�A��G�Y�J�����3��իW�����3��Q	��d�<������Ɋ�4���ԨuԄ�.\8_a�07�[Ye�c�t��K�gHS�V T+Aذ��֠po'�P4y�E��ݓR��L,m ����+��@��5̓�!�B&��>$����+cg�U�9��6CkK_#VV`��ns+�/�@|���Ȉ9��ф�������JV	  ��P���"/�i����(�b)nW��/g��,T�Z�[����FZb����3+��J�!���\��Z���}� �\[�y1�ܢt�j�)��q^�~���8����V*�R.Q�s�ww�o{��~�O������K��w���Ї��΍�_�����\0Ņ����Ī�[���z����
�)C8,Qpe�4̒�;
Pa�@`]���������_BE|@J��yZ:���+r����2����X�n�Ɖ&B���y	��0WCo��	`�����AdP�$����J[k��p�w�8DZ5����#$̥�{q�|�R$�W���Y�^��2��[���!��D3l�����n֝U4JE��5�ż�������֪tl�E���g�l��x��ȵ����e_d�+�tj�|�С��>*?P�a݄F�! ����m#Z.4��`���v�x���URd����H6�B9hr}��� �<;�i�T�
!�id�\���P0>ׁg3n��KO��&t}
Yr�p����J��;�t޵���_"�RÍqno�z<��֍�E>�΀�,��%�+ ci�۷J:Cz�H�X�&{3~���U�?�rk��Q[Q=�p�Z�H�ù��	��������sdݩ�PѬ+�|���OEC+��	͡qo������|	�x�u��*�VQp9��p¹�M���~�^���U_�Uן��'�/���}������}��" �b��Mw�Y@��IVw��%ti�-L�P���T#��A406�hh��3H�Һ��xH4�]�����, BZ�Ts�1����o����-tS���a�q;�iH���8��A��H?�����\�о9 �Y �$xr�t���̐r.�ҧ#���V�&̘�+a|+㔙8G	T��1�s��
q-K>�V�j�2^>�!]9@-[+���:����LR�YQ�E�h�sY?��!4�QhQuz�'0@qՖ����V��y"	�@'�/���;��<!-<Ǯ�)�6� 20+«�)h��Rs_R[��h���w�0\�����N��j
%�K-Z,�5��kǙW!`�yi�xQ>�fAAOh�k��`aB�
�=�/�Q�*JeV��f	x
�J�0��.S9��TI���<y���t��Q|��3bI5�l��a�5	�@�]���S���*�q��ڼ�ݺu3��@?N�_�l���[�wɄ���j�������w�X��/�P0hKp&�����3��]r6P�^��G��3&���W9�08���O|�7��?�5_�5W���������������x�9 It���ŋՁ4]
9 �~�;|$5�"2!���5�-8g� ("�	���rS3��9 B5j���r!�LnEYŒX}��*�:�+fI�'S/G�(v����
��<���sX�6����_�h*2+z8��K�˽����u0��kp�f�LJ�.�}�'5ܾ���GW ��7�����M�J�R��(��8s4)1��(�2���Iܓ�	<`�������_F����� xk��f� �Ƞ���V�ZZrX�Y�X�2���@�5�A�%��C&��ZA �-\חq2Ь*�S9H���� ��~Z��T�1nֶoY)������b�~	�)�쵀�w�ᙪ�
/�[so��p-��X�AA����5�pl'T˖3S��e
��g^��>�?/, ��9��Iڔ�B�q �.]N�����{og֮��	�A��fw�����b��A	od�"�ȞD����<��#���-pa,FPha��t�Bw���M��u�@�� �n�pys��;��_y�۾����$��>�w��'�����}<��R�z$7L����ݥ˗������ �x^��CU�-�'�k�I/x�iV�K|������F�ļ�6d�<�z��kf[р���
a�~��qhY@1��ʆI8�bz�Ѭ���*�&��5���(���8W��1��|-������w�RFG��wm+���,z��Gߊu������[~�9��a�Ӛ]�����F�8��19N4�`�MR��Y��^����!]_��$���x,(�<�����~�1G�~�~-:C�ڣ-���Э;рU,�|��UX#�TR\�Lv[���@k2}r�ST�	I�S&��
Fj��6>�!� +Tm���xg�Ga����c��2?s_�i���B��҈�z�+'��W�!�Y��ݸq���{j -�;����_��	 �HC��;�JA�A����+�JUɠBCK�����$AI��n=���!AR7�?���b%Q�R^��W�mf�@XAM'����g���"�{
 ������?��>�{�U`͸\���������O�������z�O��?��������1P@6��ًݕg��Z�p��Z�=�`w�оi>���ը6��P��fP�TY���l ��D_��s�@�藓�C��G��x���L]�JA��`�J�������%p���I�s����D�a�ѐL�$0[�����(��o<�4��De)@�NKI!�6XXnӄdj�2V�2J�#�Cڷ$ЄYG^��׉��������Ȑ=����&���
{�1�K����	��K�.s�?������:�YcO��Dz1o�K�9CX8�o��Y����� ��a��µ��V�K� 3�.h�Yj���R�byVYͭT��$�Ja���F�{
3g|F*�T\L�p-k�2҇P�z�w��f`Ri��PI��̅FSe���V�͒c/������[�
��<�W 5?�\���%\>����g� r��2�����I�w�+��,������L���c����_,���*]�<]tU0���K@eϒa�3��.�o�)(�#��}�(��U��������3�k���^��\|�	 �����������hooﳘLɇ&��>s��VI����P��=Z?9$�����߈x�(ZL�ﷄ+6��� R��(���8�@��.�L=�2�HUT�9� L6�� B5 ���s}���W��Qp*̝9��T��-�[v�s�y���g��(�A��0�SWC8M� �Z����X�QxL���T��~��y��6�j��Q_a`���@�s!8��{Fر
y���j�-J	���G�Z���]�F�h�E����޹?�g0֭���i=r/�9��/��U�6�r�J�Y\)�8V��R��5�m-��f	�
�šeN��cy�����S
�$��``�B��	U
�2�md�Ʌ�.+�9��|'g6{:��I\�ɞ!X�����뼟�QeA%a�ތ��������y��Ԣ�z�u@g�?��s��J�=~:�)�4��$��U������i�Ҩ��u����� J�{���u��E�����~6E<J %2�h���l� �>��hw��.}�DOHx���A���c,7 ��ͭ��w}�����y��^w��(���G��O=��[���I-.�]luO=}���N[�D�M&���8c׺��$Uiq N?:łe*�9��})�7��oL`, ���~�f�I�J��G�6��K��8�h/�T�w���@�	�d�)�Ih2���荪�h�:�c}V(Hl��H��Z8$M�H�6�s��M k�@�ZI!�n�R�a4�S)��w��q �Xj�Zi����$J}Aj�2-���XF�f�?��W'�������+OFA��?gs��z�g|����m��XհeDB��$��f(�Oi�R'��a����0H9,��P��?�>K�f�e���;
,�� r�Y�1���i�҄$��z�>І��V�s-4���
�h�
,-%iG�@%���@��'��}ss�%8AG0��9�_���KI��i��YΡ=>�"A������
�%�9�XV�
�5O��Z���,h�r٨w9?��Z�EA���Q�=C�?�E�o��E�U�I��!���m���9W(b.���Y�S>X9j �D�egwtk8���^��o��o���>���^s�������@#��� �y��b�@��z]�8q����<�E��B����	�$��K a��Xd���2p�"��@ZKF�s\�&�b��
�Z���(f�M�D���v��g����n���B��շ����?0c������@��>�
B�K�����6�YBe����@���a��}�cXƤ@��v<�.���.�
�A�9�=|6�b/<@
{�S�p.a���O&�O-/;��\�戄��>�D�}2)��[H��M���'�_�п��iUn.A����.^�F��G�\kd�U���m�p����B��:/M����e,S*8��T�s�J��FQ���L-�.�~F������g�sC����U�
�k�d�**WZ�!�Y��7�ŷ��
�7]�UP@Z��Ok11G�#R�,���9�"YsdMF�Y�m��V�0�hE�����0�PE����u%&@����B�\�b�<� L��;*>0:�b}F�	��<�0�A�%������x2z�}ї������8�|@�o�����Ͼi8lL{������Sg�[�I��w,f�\w�����D̐�(6��GRE��E������.��\F�bCL�@79x �F ���L q��v'���p��Rlr�6Nb��+X">��)����hy���0�STa��1�=����0k+�Yq:�k�}+C�ۦz��H�G�>B3u�ԨyOfB�|Ƌ�&<b~H_ q�#׹�2�I䁫�Ѳ��&c|��������7sa��A�¾L�?Bj(�Z{�4�kW�v�N����܅��������Z�~�/Ln5��/;����'��@�1޷�Ng?�_� ?���I�_��+\�U(�Y���2��cS�H�쯽��N��2�N+���V˯����!Qk�?C��0EP�c�)���f� ���q�9_�:S �<H��΃D"�P	B ��k��Pč5���Mr}6�UJ���ך�%�7�Vܸ���b��ܬ{)X#����`�M�7�ezJ�G @�	T@�li�$�
���*���H��3B�����<�� *�~�w���~������}��kJwע�&�������x�ҹ����{�P&�=a6K ݼEF0��5_����XL��w!J����M��>)A��3�
Ƙ�a���a<'AX@&ۺW�<65�5K΄�I:L���B����B������e�\#u�@�/�a+`@��x�:P���8�l�_`l�������"� 9v5վE�gx�7LS_������42�c��k�3��C�Aj�D8E��]����aU�X\�ykűΎM������a��,zyы^TJse\(j��t[��V�Bj��6hfG���D֣B����3&�G?��
Rx�^w9k -k���q��F��SM��u��Te�X�J�2{�-%�	#����+���O�I��W�d�%�Z+�"c	�ưy���`UT8��A�������	��>DH�Х�:,>��`�H(�������⡇*E�{V р���'�u����ř뤕}��<�Q�߀��^Z躹�n�P�Q�Y��B�"Z����ѣS�u.���!�/�s\է�����#(�S��s��Fi=��>�ݩq)�6��wv�ۿ��_�߾�u�{�Su���h����^}���7���X�ߝ;ݓ��.HPAp�ֺ�N�׭�[*"1��G�BB�x�����'�k��ڌNA��@4�ڟX}�pume*�
��<{ИD�p�!7U��0���$��vGe�"p@�*���i�N H��� 2����<Kg$Ģ�������S��}�@�}-�2f��{��Z�c������o_ ���~��{x�c�2�u�Ps�B^���2��u�T#��̥M�C�7��ӧO�� �[�u{}ʜ���|�+�}.4RJPS��Lm:�����'��z��3z��#�`��9%ꉵ�[V.@��L�-C���.������i>�;H+��d�3�8Z��s��Y'����O �$P��b���cޱ|#p�1>�u�~��a����YRh���CW9��J4�$E�����OXE���y���blZ�õkGtZ#    IDAT�L�AM6݁CGR
�Ap䵱�ˋ��2{{����щ|huV@֡CS�D�.:ك7,=���d(
��2��w�¥)�Q�A:�įŹ�;����{ߗ��K��h�mo���r�����F/��Wy@�6�'�|�,�jF7#�k�ݩ��vGSn����h�,VEc4x`Zm��ׯ����\K�W	�֌n
�Ts��a���Keq hL��3�����_�S���}��z��D�D�!
���9$�8R�v��+�h1����b�-u+�Tî��� F@��8�ul��J�H�񊧛C��^�V��R۪��V�J+��y�4鵲d~
J-��ȍ�c��Ȁ�Y��a�N�ɽ*�vx5U>������1��'0��쭚+[�`C��X_����H�,��%as��+׋m��4��A���b����x�r��W������a�M��:á��RE8� U�V���K5�j�������Pdyu�^���%Йk�\U��St��=�}������(;	�)T-��}�ݨ<�0��'�Ղb-i����
�T�������VUXIQXi�]����}�S��r��Ү��ځ��e��[�%����z�'�gPڔ����>V�,Pd��Z_\)N-��>�bY@��( � �V@�C?�p��1Ͻ�_�e��m��mO������i�����_>{�����/E U����T �ߤu�|7 u�W�f��Xwω#u(p�A`�¨�h���k1;S@��n�l����" Mi?ۉ�)���|�@���RU%ط�1Z/z��q���Y�����d0^Ni�`��\Ħb��(8`i>�y-��� �I�k�Բ��V�l3��0fP"�"��d
m�Y���&�����1�Y�J�	X��իIk�u��w54�V��	�	�<�{F��:�݄��7'Na!L�Pf�	����#y�Zn�wD��?�M�|�W �{�Vs�t��$ha+Ʈ5��`�=�p����׻��{�����ܲ*Q�Pz"X�c��
Z��b#T��wҏ�֠���{�:����V��j���Z�|2���
��Z1eI·�z�s_�8��|g߾$Z�߮�e|�G��j�!�(;���3QV�y 1����D!��3aT�k�� �b��V!�
x��ߔ��w�a�h	�;w�J.}�j�Ʊ��O
�nnT��Zs*���Xԃ�M�/E��7�XY���SO~� �(пJ���@�م˗��N�k��
���cG��0.��w����}/{�˾�y�br�x�?��'�~��&��clZ`�AG�'�z�+�-v�+%�V��>z�;���I6+�.� ���/�o�<�tILsC8��ݮ��̄����]���-Q�ku����L �qZ��0cKѱ��e'n?P��*!�	!Ǽ��Z��U��� 	/n4jL--���-�y������}g%��QUiph�AM�{	�c��{
 ��X-�A�eX}CkH)���Q�pp���o�0M1�%|�(6��=�8xO�������
Vi��'�����CU��=���p_By8�Le�j�8��M�eSXS`=�y���b$���^P3����a$G�'�G�2��	*��P�eI��GƩP�[<�R�-�Cr��.c㿖�B_z��%�ƽ�vm���S�>ҟV��r��;����;�a�&�d!�  *>(��� �W�]lwX�^Z�]�ޢ�\����-��j�I[������W!{��f�IP	>G �!���o�ڤ8m
�z����z��P|��Z�+k�����Z-T��۷[ؗ�O��~_�r�{���%�� �a��_FX��n�F�����_�ƿ����Qp%���Ͼ�ӟ��?�LF��D��L���O?��X��u��na)����B��>ҭ.�τ�H���/������:M �N�h���d�ss}�?"l S��ZJsԢ�۝'�M/�00����"�J4Lg����2��J0m���	 EY{��@QK�T�z]W���;2�
��j"4�9<���/$��s��K�Z=j�V��tj�'#s��\�IȔ9h����I�����jpj���^B�&s7�e��G���>N�5;쁹�����|m=�ʙ?�a�������&���ҦS�xm�v�.��������RDnp-�>���v>��8Κ�|��[�rV4��z.�J%ֈ��z�*mh�Ms�*��Sq/�n���E�k�J�p�1@�ĳ��gSMZ����Tg�ub�&�Z:��gZg������Mb1r-��`���(�0� 4���U��kB���,GQA�/�:�N����[�ܷ�� �H:]���`\���i�*^�"����
 }�%��K(IQ$h��C+/�'{��� Cȹt����a"�P�O>@�����cg�����h����s���^���>��"����O~�?�u����ٚ��/�2�>{��z�f7��ԃ�u�����UD�vp����B%��@�S�L�n��� E�5&\�0ؽ���݄�.���oy�[Y�׍��]Q��C E��ƹ���K�b�_S��<�H՘���N�n�R�b��i�0��d ��k�q�r�`�k�I>2��j��DY�s@����+bq�q�- ���-���El��qsƧ�,���Ɯ�i���gf���O�!>É�{Z<�gj���>-sT�&�1?�3W��x=�=s�Fw�R,����.Ģj
A"2�bz��u�@����yA��C��F������"�	�ݪv ����W�HGE��Y�Za���m�>�k��B��7y@Z��h�hO�^�~�IQP>��Y�z�����^�A�&!_�u����+J�%բ����z��l��n��u��������)�;�+6�Ŭ%�RĽ@�\*|.*��b��g�k,� 6�-�v{#� z � �� �	J�/�I����D!��E �\di�P�OS"�[MW�m<i&��(��^����z���P�@��vwҏJZܛ�o������/���ᯝ���������菾�����xnn�y;;;���(�v�=}�|��;��nqaI���V���p{�{���Z����(XdY­���P�\¼���"@��2�+�Qp���_��@�,W B�sp��ih��l�������d�8������B�Z�]���
]򜵵�~h �B�h�샭5 Rc�[F ���/&⫬�NA��z2W����>��~_&�!�����RR�;���F�� b<�W��U�́�3� ��6Vqi��j�:�y�9<�&�=�@�\e��:&���kݙ���&���N!�j8H&�T�QL\wrѰL��G�O}��t��b$��޹����p_>/x��8��	h�]�2�_�ǣie�Z_��4�)�O}A���U"@��6�UuE��~}!�zp����pU�7��6l��rO=���I�87��Z�#��Z� �&���xJ�D�k�3L�e1w��Vu���"�9BC:W9#��^r��&)Jn����W�=ֵ<5�@�n�ۮ���56+�i�9������@�Y�S�Ln�x�����?�sYĭVc���9�{�*I������#+�h���� �+!4�����7���o�����ϿR<L����/������L�p2�,�s���QUþx�r5��tiJ�"���YE��~���"9��|�����NL�n�� k���B�J\4�@p��e5��.����~��}kt�a1�����4���J�]�����@� �TK�C����Η��Ҭ�`�9�Υg����h�[�Gˉc�K33��IeDq1^}�ؒ/�ijxB�p�@���_�����QS.ys`��//X�@�Cƪ�%W 1}2-�oXn�k�sh��2��_�#d�m�*7p5��|�\�y����K`���&yN���x_��T�˒������t����w)��T�&��ZZ����^�*Qh���[&Z}� 	������x�F���"��n�Z|�O�#?h�n[�2ZvUL ���5��i!z��;�Z�Z�a��@:�9o��N��M5!���NQ\b�yψ2�Ui��4��Z��9<�3�u0r�~2_���#����ځC��ʇ2�����-�߹��z>���n�_l-�Q$�B����"ܙ��@�I�ﺍ۷+�%ֶ��PG�������X�X��k��iWU�Ac�]z�>�,�gJaE 1ks�Y@uV� ��#Q�40�]\�;;;76�v��7^����y+�~�'�����I7����k����*�p��3	�,t��I��=��uG.��=�(���=k
ע��5�Y��@q)�ǻ�?P`U�A|K���2�(Z��'7`u�%����[l!�h�9K��s%��� м��EN7��΍++�#([���9���	޽�<$�T�u�����DJ�+����+S�D�$3�M� \�OL��狹�k)q��O,�I�3&����z?�S���	��A��x��O���(�c�z#��oig[����4��"�	Ip��G����'N?���u�=�X��sg����bR-��¬��Ǫ��B�1���Ҋ(�8�L[�Włb�bb�ؽP��RL�A/}E+�:̂�"�%T9?�c#d��S!CKO��җ��4T�f�״tk�[$�*(��q��JeɽU���<����t��׋��a��(Z-ZX�ꕫi�� �XSظ�g_US	�1�sV4N������.�ou}᷃��M�Y�s>�pŀ��u�+1t��6�e���+�׍צJHL)u���ѣǦgH�w>�t��J������#��hG�B0�]�F	��B���V��N�,�����K�����p�g�鯿���}�i�3�yW!����w~����������`n��C��йKW��=han�=�����Ǧ�EO�t"�4���ٟ�ډV�0?!���KY5 �cC(h5Ct�b|.�͌���V���U�^R���܄a���J0��V�|<s�Z]G�i4�8�v����*ٷ��Zh k��S-�v���}���]�*�H�Gb-&�p|ǭf�Y.��O��ss7*��iY�	�V�S�KJ�P4�0�058�3V8�kZ��ߝ�;�����\�E���*I��	����^%���z��C9���u�<�����e������\I��g?�YY����j��h�u�߉�,jQ\Z`�<�uPHi���q
�c�%}�.Tֈ�J""�e�`le4�V�r��U��ʉi�f��4�n{���hЏ��Z��#y�"T���͞����pn�a=��i��K������x�ݽ�{$��Phr���Jqj��@@(�����{�h_�t��O1I/4�8�?�0�|=s���o�Lm%�5>�a���R�+H8����s�K\���#�S�qp���s�� ��F� ШDhW�gϞ�]�Yn���jAp����k��f2�~����+���/}�����U��w���~�?���F�ݗ���1Σ�O*����K�-��I��e�;�?��5����Q\ez.��ML߬nK�"�/e��Xu��ʾ���>D�����@2O�_��6��+l�g8�!4�sY�����T h�m�� ��q����d�BS���"��c������{	�f�
��$@�)�{�W8�z%px��h=LOÑ�3�V�BѪ�B�C���X�����[�*᧡�2�Jv�6��/�s����3���}o�6��Z�'Ow���u/xዋ��-�p���b ^�w~�w~��?%뿺�6�2�͒͞h�wn��%���zt=�i����nT���q/}�ENZ�&f��ٟ��h;���6kF�(�e�]�~_�P��4�fY�gҘJ�H��;Z�AR�F��߰v-b���&D��29\��{0�h����!�x�n5�fq�i�{��wO|y��ȘFm��������z�#�pU�lEd�7�����iݾ4�ݦR��Vw�ڕRh��P�)T�_J`��s��YG���� �UPJ���)���{� :���j_��p�u���R�FI�&У�W��w~�7���}�W~��!�/��^���ۆ�;�\X��W�c	�cН;�;s�B���+S�詓��#��چ�n6�4�h!Z#����Qc���*sg�,q5fxE�T"��T a1D �v\=w>&;���$Ȳ�t����}�#�C`i�����	�=L� ���R��0��Che0�9x�����=9\��0���{���n(�y@j�2׎C�sU�#�A	������XJ#l�����Y9��/�PSu�x�ڶ��^2v栰��UAD���VV�K���:&�UB�%7�M���C��G�������CG������?1���?�OTݸ���^)%��d�Z��hZ��ڮ��8�7т)8͚n�͟z��D����
CM���J��b�k���L a�#��5�`��)�mv��R+����@�����/ZBZ�Q���b&t�5�e��#�b%j��_>�V�Mz�����x���[A_g�E
r��&@���>>��G�z@*qB?��0�����T����n��@p%�����]
�z���?d��/oH�4^Q�k��s���H�#�Z�@p�$7_M,�m� �,��*
�駁�Ӭ�С�çN���l�&s����_}�7��y�
�_�����W��K?�����-..���_�.^�ҝ~�l$VJ��=x�=�='�M%;���\�g���@}��3E�U ��R �#����"@���
�����%���U���)�b���uǗS���olŤgX�@ ������A$���c:z4a�s�\��9q�XE�!���_�4@P0���Np�L\KF�����3�]�5ctѴ���k0>%�Q�ˡPpT�*�V*�K�K�kJ;l�����
b(�`�Z�BP<���+qM뱣G~C�;z�{�;�ّ���W����j��>T{��'����oe�j����|2!M�5|��,pr�XB�k�/e��T�"�uѷ�^W�-,���Dp��=MiS0*H���W�[�60��e(9���d�X�~J(PҎJF1��C,��	� ��Cu]�S�V�B�j��NZ����s�UwE$�~�\�
��_�������\�[�x�{	�I���oa��I��T��Tp�� 0�x7a�@�տj0� �EEl��s�gn��
�@�3��s�����d@*{$L�����[$b�oz�;|�`!�����'�\��wa����o��oǟ���J���uW!�����_������;_���P�|�N/.�v�.?�=y�L��C��r~<��C�|�FLN��X)�>��`�����̂�zmS}{#�vŦ-N�Ƣ�!� ��Xt6LH'L1k�A|D�8j�[��6�;�u���!ҲPvr8��;I'X��7�=�G���ߘ�	�$�A�ȳ!��К�gh}ᡓv
1�����<�_!PB��S�y�%G����sʚm�ٲ������1���Fۇ�����#|���:�=�_������\/�-Ѣ�o������Б�ݑ�Ǻ��8�f;Z�+ �N)#y��1�a�Z�T���D��'o���ӽ�?�5��ge�CK�O��\��������@G���b��$�SE�=5[��=w�}+l&4�=�������̃���O�5��,�Z����Ƹ�֓
�Y=�u���6%j�5�gYfKi���bǏ}�beB���e	�f�.�Tɬ�Ǻ��i5����`��2V QA�D�ӷ:mHG���%P?P����h_��@�9_�0x@ţ66�3g�t��[��nTHT��ml����w��������,����7~�WN��������;aii�(�X��ʾ�ʕ�U�tsk��5M��a~�='��N=T�R�    IDATX�ː+�q9ƃ���@�Ȏ��M7������ք{f�0˥�R�0L��*�q�&�fv0�C����}BFY�Ia}�6��"����������B�G����F�%�����z���6c�`S������^��E#��k�}��3���-85߾� �?�?�Z�
���z���b�}A�5�~VS&ˋt_�0�����?{����)����lu+�K���k��#Ǌ^�d����:j����گRV��A1���yVx����D5_s�o-F�M�!��ה�a0(:������SN�2�f���F�a]�7
���JT��bB��#�Boݹ]�W�R����!����B�"�^A�3~����e)��	�D��]�O}z�:
�ca/�!o���*iʝ=�����\�
 iI:,�l%�#�<r(����{��E�I���A����X�ԛ�}Xh��6� W���Qp\O�l��=#AV�_���R�X��ļ,b���o&���F�S���wn��G�I	�S�_����[���6��/,����~��>��n�ٓs}�n�}>�=���7nn������	qee�,P�f��O?�ݾ=�)7��r��ǻGy�0D��&�L�V,jb�`� }@B�Ah�c��/�,w�h��b7H�Бc�|�B�<�/\͔DrQZ�9&8������H��8�F!�Xo��QB42��f�1�d�Y�Ǐ-_�N9���[Z� �grp<L<��?���!S��1K�����G������C(noM--�.p	֦@�}ƣ���RH*�Js��̊�z�AKs�C�x8ܙB1>�9�|,aR�&�M�B��'���Pͼ4���NB �+�-��%B%���6�Y!ڇ*c��!`�jY_�o��{N--�V|��D:NE�(S�nk#!�TQ���bieV[�1y��S��ޓ��)��|Zb�԰f*����:�6� �;͵�<��jy1o�/P����2��Bӌ���\G�_h=�A�w����pŲ=z��sV9�kJ�B�:��K�"	G!
�`���k��g6 l:e|X,k�%� EV9�U�q䲴Z����.-_��Z� �^�
�������{Q�puP	���\�x)�D�U�����������߼��/�}���]@��䇏��O�̷\�y�o����s����nw�~�t�"A���9z�{��OA�Ư��&_� �� �dI`ܼ80Z@=�0�W�vy�[��is�)�x��	�&�-tC��gc�	�c���,���6�.B a�l9|�ƾ7L��=�$���&���ǓY��>�V;��U9$���!�ZKυ�x�ɧQ$"���Ch2�	�n�?ߓa��V��	sD��`j�}&#���*P�H$�c�?�O�4�:̓�(%�(j���ZT�ω���2���k|�����4��Ђ��I`��1}�ñɰmX�5�]櫣]�{q?ּ�s�����:����Ѝ�9�g�Z�C��Ư��8�:���]�1�<�_����>�3v��x��r|�3�෽i ���[ֈ����5�7.� ��Є{�R	
Rê!�0�롏i�7�!1e��V,��	� �������?9?�i|��c����]��Zu�[�{���+;p�Y��
���T(�#�B!��3a	����YJ�,�+��D �B�% �ƛ7��(�lyL�������������>�h�����
�O�������.\8��vwv��eSn��.n�f�!�X�#�u�>�H���Ìb�;��j�B�fa�5%��̼n�V�i�]0��)x��P��oI�<��4�
�h�o-!-�	P�ƬV�b?8����Ɲ"�f����8�|1�^gT�8��cǎt��oZ[������p��{�~
"hLY�ć��"Sg�@ɬ��@2U�M2Ʀ��
��(�|<�]�����E`�1/�g���A#n�u�V���H�k��x�����v9l�[t �-8d4� Q��/�2`�[��迃1(�c�W_�	�DU��\�����%�Bb�
�4�%uS�
�FZZ-�����6_O-5��
;���\-T}V<W�k`�(��Y!_g��J���b��.-�W��A�����_�z�:�q�
�U�((n;V;���>c�9�g����ʷ��uRAb��G�8� !ow�VR��ڵE��*Ee�,�X�)�3���$l5�چ߼Y�o��2��@�w�Ǽ�,�z�!2����bȞ�(���<s�$Jw ITea>�-4���dwo�����Mo}�[?877�u^wU �>}z����_���O�/�흗�9t�b�����^w�����5�ܶ*�0����G�?R%y T~nU����Y<�����#nM������O�� �H����M�I�o�e�&��g�	�5L�=�Q��&�/�JS��ԳΨ��-�jߙ�=�Tcch��8�~�O�i�	�3�|�0��!5�Cf�3d��ؚ?�C�{j��%� �
�h�姚8��K+���eѵ���<�O0E�T,�d���Ǡ�U �0�"s�����[ ������R7XD!X��=��j-�Ha^a�=xQ!^��M �L�+��� 	�2�g�����)@�,c1��AYM��˜R]bk+�4�(O��h<�\�V�J��*���>�򽂅[�w�Y�B� 0o�WZS(�>�^�qw'QmZ'��SB�WC��e]2��񺮌G�-�kg��]�>-┹9�mWtڰ[[IaC���^�nY^���(�a�AI#hE��Z�P�?z���[7�;D���D�x@�a���(���=+*���(������8��Ecfy���̘]_�ťKWJ iq�ȓ^�P���0����pwo���{�oy�[~�.ȝ�-� �L&����o�3��~��p�@��!��{]����˗�K Q�#fҝ:u����{�8K �`�.��{E(��3-	\�/�����хշ�JPmr@)Gm$#-��U�63yu�	�A3��l���`~h�94������M�����Ҳ��C�~B$��(F�6�����QVi�D	�;�����4�K�aJ��ڻ��p����T#ԸFM�/@��X-~wLV�K����)DZZ�|_�B���k۷�������IK��[���M�X�.kZZ3-?������i�ܳﳒրuy���L@�	H��>~"h��aJ�0�~�B�+,�R�3	8Q[��4�AߪB��V�]ny,�X�@�U�Z@��	�i%�,�~0J�,t���zT�L˪��l��\`M�?,r�m�{6C�(�$��5��a��XЁ)cm3���R�f���f*�S��1���k-�l�Ҙ�ܩΦz�U��${�T��VJn!��TB����;E�(�(�� ��r@
W�HP���(.-��k~-xJ�`\
�R`Z��������/y�K:�,�?�'뻽��5����W���������
 ���������G�:�����}��@�@p�n�;w�bw�µn�2�����v'O>�=x���t��z��/���/�<�b�!#�4��N+�a�W���aP�\��Ւ�U�� �~��0��� d�a�J�$EM���6��u�7��⼬�v��:�󫿗�v�����ܷJ^�ku�Z��ڪ�1�Q���y�YC4�XS���!"��V� 2��]��w�#�v�<ZC��ZI�L-�9�ą����+��%�)M��jȭ�e*�g<24>7��]պ��"���p�c=:�L�ߵ@ ��;F��
���'C��?c����*X3!�>�P�78H��A�&�N�C�Y��ڃV��	g*��c�UR��t
�Ğ蓱
�BD�
��&:>xdZ="4��8������8�PH}�=`�՜�Bp*(<�1���+���=�F�s\	�m]�g��$�@�uʩ?.��� �.�T�W�"ڭ
/,�0�i%���-%�j/(�P�yo�b�Ql@X@Q�[�<�<���Y
�\�@���34��#�T�?����b>��G��/}��_���/��'���g�_}�G>��o���z���`���w�K+���rw�����9
���"Qcsݰ{�����(L��� �r��n+p�	 ���Xj��ْ	�S��()7�4�nP�b�$gu��*M���/aҬ�b�s��/�YO�\�{	_ݟ 
+2T����2���K�Y�}��c��,� 
Q%��Jf�Cu�-�PPˇ��Y�V����*ӖIr�͛�-<�jK
��P��B[W�Xh;�n
֑�LhT�ԢR�������V��Q i���j�ZuB9���A�@1v�c�i�M���X��q�����e|?~�0�(!�0�X��P��~KCma�j���}�˺	�1�XM��iME�I�k�K"�R�Jo��6��*���4M9���s��Ώ�̕�^��Z��t�>h�����E��ik�Y[�?���%+Y� �!�X��N�ZyNu�]N"6����(���jl�ݷ�
֝K��S<����2f]Uz���oDAO'�sn��ۨ�k�'���\�J��Xgƍ @�5�������4�K+Q��q�˷�zŷ���$|�� i��#��T�&D�g�*ĵ��/߹u�֍�����[��{��+��鮽�*Ǩ�������}���ۯ����O�nY��ݹ��3g/&{�(��ܨ, P�)�M�H�RYk#����̕�"��i��YP�g677��^��]Հ�'U���	�C(8폞8>M��v
z����u�����(����l�U�&:�0LFE9�k�i��3�(����"J���S�J�cń ղ�*hM�XG�RijM���F�D��C�oGA�3dD>W��uD�$xnBK3v����Qu8��C�%����<Z�Z�����:ML��J�� Z)Ee'���Pj`�(�MЕ�] �Пk)M�����~3O,�K��ܼ4C��((2m��q���h����,��@\W�T63�C�K�g�$l
L�}��͠�(Bj�ªп/��{xM_q�Z�G�8/|@�/ f�OA ����3<�`4:����Mq��$�����΢�̂
���7n�s�#��
B|��dxc��
�ss�ݶ��
�J�۽���-+b.A�u%��F��S����
+�RV�k��E��������������9c�y�J!��'�;w�~Zy����(k|�:EJS�w��������x����_�_p�z�|�(k7����Я��������]^^<S����v�Vw�����
N(�0��l/|�#I�Х3�E�0�� ��F��|�(Ă����
s(��p��FSX4�e@v0/�z��Y+���p���iv6�1K�zv��.f���ӜJf��Vm�+l�eJk*Cd#�����YZ��i<�CD�1����ؤkg	^��fY�<���������w�
�2�[X�Й��՜�Zߋ���Le�V+�4.O�'�d��\�J�|E��x�X���l�	�M[�Z�*(�p
Y�����Im׃��J�kT�q�Ҏ�8��H�k,�ﱬ�F���1�\���������M�"$��ڹ����U���O�.aW�IB|y_˚{�C�2�`��Ҫ���:�e�Ф�缤@h��9O<���{rNu^ZG[�3KH.�c\��,�?��Ϝ�{�C PByq=�}��.fG�(���g����ό0�-��S��?"G�n���a�7yf�7�	�7}x��!�ڇ���9�нVe�O���K !%� �>�(�	Z��j��0W�d�9v����{˚�Ba,����ή���׿������kU�@��������+o�y��7.-/�@`aЊ�ܘ�t�oou�˅�#��_+���pڍ�`�a��%� �s��0��L@�
a����c���DY:��r��G$ȁ���ʳ�����ɶD5LT�+cљ� 2�SfU�0��0��J�T{�1ŗrp�Vp"/w�oݪ���Ik�ȴ���X{Ʌ2��)|���8������h-�	����,�T#*�{v���rly�3' 
�����*
}� �ƸP0
�
5Sg�kV�(S��#zL! ���� ��ڦ�Ap���c��Y���ʐ��'�[A-sQip�e�
p�#��:����z�<Z	�V������|-��f@:IgQ�)���o�WJ�c��F�LU
~����l2�04��;�F��=�hpK�Ă�A��jٰ�zw��4칫��~�~C, �y�ZY�q�·��W&_oܾS��S�����Y�X.��h>qƵ���M�5��u���V,��,�a?�b��A�(���9[q+8�}�(Os�� �j�(	���cG�Ƶ
����F��������������/Ρ����Ї?��������׾}~a�d��^]��Bwgs��x���͍jJG;@r���B%�A���/VtY��d�{���0uK�Nb�2� ���Yx���?�AFp�@d��I�������[���
�ˊ�kP�	}jua��0�܊�b\�5p#4B2s�v�1O�����P�^@j��Om��#�85h}!2G���;p��������EP�t��;�������U̬�XA��\��.d�S��|�c,��{֦��r|Wk�kU$���V+D�"a��*^;~�a��T��p>���|��|B��%�/L��dܖ'��)��Q2%�?����$���A��ZcL�Cr���W�@���82�\�4f}W2;�"��s=_2����B;W8	���´��~[S��y���Iq�&g��h��H:���^M9���bw�_[�`���B��nԵ�ީ��kT�;���������"���������,"-�d����-�B�ZR*<����=�RLЗJ�����OO���}߉�Q����M������|�����|ӛ������}�
��}�c�����_���շ��C�T(f��ם�p���hˍu�� �Q�g�~@q�� 	���lY+�13~��@��u>�-��;Q�@&fk�PC5 Am0����e��2�!���BLܻAY�2j��qHDX\��Y5����!Y�Js�b^]hiTWU��J��C��22��SA"\�ג2�8���R��C3&�DL$���Vͬ�����f��BǱ��9�}��F��4-�MƦe�X�q8g�BYS�
��3{֬����fyN�Z��f���(ƨ���(��s��jҚ׊3���h�}����-M��`��4�� Z�S��lE@*��\��w�{d�6�\A�ƂL�֥2[{y>��F�I �%w��&=@�;�j��t��N��3�^J��;J �>74	�B�Z������5�Q��D�Z�>���gZT[h��,:#>�L���o��S9��5\
EC�©\E��YG��mY��VԬ2�UD 3��o1������籦F�1����pss�?�꫾���{��>z����6w��L~m��o��/?w����M����d�w#�.]�ڍ�������꾕��v���O����j���X��-s�@���J�3�:`MH�9������d��{Id!�̈́ )>����&@��g}�Yy�}�}���hf`� �$Ą���a- �0xׄ��d�XN�X�`�Y�0��B(t�ѭ�}u��Q]�]Y��������o� �3`oFTTU��������&K�Κ��|:l (g$k��r2��o�'0�Є�Q�����y�k2���CJ3�F�p�='��h&f�˖��am�{����P9̶�����ִQ	�I��r�k�ȷ��If�l%�������U�Fs.����{V���!0�i߅aX� c�`�p\��ʄ��'����o}��o^o�/�! k�f��n� �s���f�+�c�f�/��ܬ�S���׋�XPQ�G4P���lR��~ 'D���V0�`��0	��/4�2�����Q�I�7=��i��    IDAT��ݸ�+o�],�b��E q֬L)\}l\�p;{��` �~]�fl�ٲ( �~#̠���dk�V�����Cح�mD�v����:���������jɢ��r��E1c�pKh��h)k*G�Z	����(���@ +>́*�!)��8�'��|����<g��k��[���U�z�4[��-Ѹ߯����e?��/t{���ΐ©�8RI�
�Q;�X� ���cGӡ�sjQ�Sȃ,�0@a~:�ǌΚݵB�&↼��f$ք��GH-H]1��M���A��̡�"�F��#/j�vh?6Ca��r9@ U@��K�`8T\˽�����bõ�J<�C�ș3�/�����[����"�2|Q��Y�e�ApX�H�(����ǂ�ϱ��3w�	G.C��+o#W,`�X��ǂH���J�daW�51>���>G�q���`Xk�O��L�(!�q������5��~�X��=�J�s�R����K Y�2^)/�R��Eǿ�[HZ�Hf�@6��p>��YX{�,(@"�(�iE�B�)e��fKԊ�֢|4�.�\,\-,-<���6Lj�������ڲ�f�ʾ��C+�1��Ỵ���f�T9�^� �Oe��OU͕=:���06��:$�Rt_H�Z�Pg+"�P~)�c��v%t���W��b��>�����
��E(JE+X-^ho��7���3���~�g�*�s)l�����#@"�j�yw�`������?���^�����������7o���?�s���ΰ ,�t���V��KWS��%��r����(�Z�,��S��1�
>�>��!���).��XLL�\��V�?��'�~��ff�X�!�0�C3�sr{/Z-�2V��23������~�=Ui	�d���	��|-�U���*�_IM�y�QPI�v�!,3r7k��,�1l��]#�Z��=ssB�����k���X;6�d�εpTh�-�(,3?ߌ�ա�No)9ühX8�1���fk���և�{�1�~��-?+4R�
�kt����ϴrb������1�d�̖������V���Χ�N������sc�ݎ��Z="�<WG��=�`Bf��QT|����^3[�0k���l�B+�W�	��M�*�o���q?Θ��̉gca��j�V��}@̇3��!������r�h-��(
+�T�熐�=���N�[[Q����R$(#Ϊz8e���	�T��q/� E����y��S�=��3EHY)�(Z{��i��mXk�isgwqlt�?~��}�/>�yϻ��B ��]p����5�v�q�כ`@�����._U��F6XJi~n6�8qD%g��{��փђ��&Ys��!��V��$P0��'�%�B� ���)!T�}p�`�:WĈ�&���`m֎���#��9���l�}Nnqo<p?����
'>}\��t4�kw#�3`���d+#������5I��>���e<
��ړ�VQ�5no��k��ߐ�a)C\���%�S���wcg��ɠm�5Sk��|Y���`��܃�yܶB���Y�'-i+ ���,Z�a�����g.���G�����{���v�֍�+��r����`JU��S��\ϴ���E�v�<U��A�g�#^h~ǚٲ3-qf�^��]X���u�%�ʴ@�s�	�X��9(�0W�5�n!��<��v_!r��/t!��������%j�M���˗T����R���rX\�]ae�y9�3�Ed/�C�%"��:>F��d�/a��ؓ5QP�|X���KϦA��Y��i$>��	h5���n8�}�`�o�viu�����/~��/o�B��8����}��;��]���Z}u�R��L'�����9	��G a>#��I��8'�ju! �d�#	�č� 3�ڧ��`�Tq�@���vOᏵZ$�NLLjS�0>C ���J`��  ��J+*��
z����`�u��P/n쇿�pOX�.�E#aHG���K�z���S:����{�`�!��5�ᵳ�����}P�u��&�>7��;��]*��6c��x>���OXTEA������;���.�fٓ`�Uz�|_h��M��vhAaX��|X͜�tf!pЈ��m~3;������ *Z`<�c1�������Pf�6��ER� ^{[d��3�H���M�K����裢B��L�_Q �"�\H(��y\܎�t�����BC]�[�V�|F}?�7�y*9���W+L�
>�`+�5�����Ƣ�;��
)!9���q�������ں��U ¡�P��L{	����U5��b��Q���� N@
3�q���LFQQ�P1�P8+dTC��u�1z�|�k�"�\��O�v�m��������L������n����}��q�ԩ������ z衏������W�m���r9�T%9�i˰�._��66w	I%�Z�41>��M��(Ș�iR���H��u�$d2������A���P͂�M$���T��p�yMLMK �Y��r�4��'be�ڵ�����z���OWe���i�;`��6�]u��0=r$��*QG�_�=���E����ڨ5T3��}B�����N�G��j����ǚY��4�Bm�}����yV���mh���؋V���G�����33jk�V|��e�s~S��V)�6��ϥo�d(Ǵ-vӏ-�k���>����1�i��,
����p�h�`��_�JL�J ��ja����=�54��Z�;?�t��2]����0Et��&���rТ+�5���=~���H���R����"QV������q*wg?�ZZ[YMW�S㠓Z�*�貗�As?5����g��ɰ��G�A��	�4UT~|W�
 d�^��1�p��T?�;��i�ʄ�"Qq�M�;��:u�M7����������l�Z��_��7������(w���.h�����?�����7v��� 0�GupZ���p5-.�%���3)�c��#��b!s��R7�>�"�D�Ѡ�o�����Ʋ��'."��ñ�>,�XR=�*O��`��ƽ!�8���FCEm)�5X�u�!G�� �&a�f��G��j�cn4���pDY��k�Y/F%��[�`�`��p����X�	���-�R�������Wf�f2�͂-�����q�?3"���>�o����B*2�"=x���Җ��[\![,0�t�Cf�@m9h^���	��:Ch���Ng%_�7d齱?��ڂ��G�t��V
���fL[�r*
K3/���V޷���̸U^�BƸ-�������yQ�{/]���<�`��|�\1��Z ��J���D�ڂ��&������A���Q�NJ��!�i�����V@ĽQr���M��N��R�sI�@@g�c�*�
X�ùTh�Կ�� �)J~���ee�D3�B���Y�X����ȍט�S���իR��:P��s󟝝��v*������7��:�`k��C�і����_|�Յ������+�h�GRi���Eq�8t���Q.�^�� �cG%v��9�ʽ8���(#�R����-�D����͈�S�@���;zR_��:"����|�����b�À�䇶i����̐�sp !�!���mE4].ziӄc�ā��!f�li����i�ٲ���4a�[F6sa�dI�i�z��>f�����Yf0��-�,c͢��"��d�.k����䅒>�S�R�����$���"�5v�^9ڿ�f&]�+}?�U)BnEK�T@��)Z[�z��d�V�lyΆ�,�ЪU	 �Y���#�*�����n���"���Z[�&���U����E��ʌ*��L����5$�����
q���
4կ��������}מ�V�˱��ޞ;EF��b�rY��N�o��H�J��cQ� ?s���J�vD�*l�Q�ዎκz���Z��?�xV�*����>���$�L܇u���OF�k�afvJ��榧����4�<8X�+���o��|��_~�zȊ�"�������S���ϵZ�K�[�F������'ϧ}��N�L�v:rd>?v$�2eM��R0����Į��P��y�,� ҭ�m-��f��Ih(4���r%MOϦ��`�9�B��Ȉ�#L娊�s3,[fF<O�KQ+���D!k�>�>xf&�;�"�����kf��!�����\G�Cܓq�ʱ��֘[��,[Q��(���κv ����<ی��ck�cw�O75ks����I�/��53�p���u)Bl\����b����s������]+���d�J�)[�I��L׌�϶���0E%Y�F���i�kVJo, Ó\7��󜘘�ӭÞ�<Y�ۇ����Ŗc7�4��LG+EVL��}��������<~h-|��;i?�����WT���3G�a9�)�Vvv�V}_mV�.�!hV��R�z��v�r�<'Zq��I������Q�7��&
2��M�����KH4��h5�!�=��~/��c�2�Z�aL��3��q�S�C�ӧO�j�$���(kP*�.�F�~���o�������W��}�?�;~�T�}c�ӞF �@G"����Kik{7���T�H������I��,���B���(�D�@&t6�h3�com��3T�rX���劬��`������<`8,���(�����G��L4��\ ����4�DE��1�� ��_C"���В��r^����ظ!)b�� 4���7�WQ�YXX�q_�d<�a��-
&+f��is�	?�'�5T�I_�3�Zk�Nr亢 ���Cj��gۊ-j���#O�h�q��5�>�#�+C��`�ް�YXY����s���ʛ{��ۂ�P�8����hbe���n/#���ڪ�LH��}�#d�	:��̉1���}��5��C!�<P\g�i��i��Z@99f�~�~l�Y12}Y	u��:���	7|nA)�6��g���L�������$�RZIO�\���j�d�����E�%	��*%��C;9Rsrt<�Q���ֺ�3�� ��/z#�.W�/"�1s���>���o��FApL�S��r��ЉS�~�۾�;����??��~�_��z�ӟ>����o����n��SN���+�/\N+����	�D ���T�gzz2���BAb�L|>�ȟk!�X3�qrd6����R{�h�~�h��a[ �2��`�
)�F`����p���n�S���G�x�׆G��R=��rjTk���:�K�O%� �@��l2Nk��f�~������=B��&n�a&n(Ȍԇ��9Ҏ�Z�i����H$[Ef@p�\����>*	�Z��>Ӊ��m�9X+��+
��3Cu�/ϱ��xMLo|PQ��Z������a9[}��u
C�o�_�s�ѝn�w��=��A$��@��m훙�FsX�}I��>W&0}�=[?�Cܞ�!<��М�*
t��34xƂb��.�V9����Y at����<�����^�2�K@e��1�"�5��@U���B�pͼA�{�F����-�$�$�"<�a�RXe���
c(74,��R�紐a��7)sd�j����ޚ7�фN�͉� P���E ��{4�v���ė~�?xÛ��)�J�/��	��/������^����C�N���p�ZX�/\�/��J�jE�y��g����ic}��\�6_@A�Q_)�x>]b$g"��!ӄoB'���H0F�}8
��>�<B�!�ad|�F��D����dM�M�Nh�a�RJI͉H�r8�-��[8|��-+�X�����$a�i����k` >��o�
��0�a�֊�|�&�Z�;�"̰I�E�d��|�y�����L}fzD���}_���l����H[�^G[�<ߌ����-�]Q�D ����I�B����B��[���4�(Z����/c�(v�ET������ذ( ��2c /+���������/B�C��r�KP��]<�* Q�}�,X�B�WE�ǰ�����2��9{��a���ɟV�9w��i�gP5��	�iblR��Hh2��;<��6��m�Cs(�NM '��I�S"���G�څ��Ù� �� �|۔�!��֛N���k79%����'q~��vr��]BVZ�]Γ��l*���+�F�!V�	ɣ���v;|�]/�W?�#?��g9v�������~�S��7�z��A��BD�g%�/^N�Q`�Xꥣ��3gN)��ֵ�>��V�}`8�)!�8��m�C�2�o������UR<$l.AԭC@B,$ˎ���R�]Օ?0&?��Ԅr*�, ��U��>�zUJhu�Q!�0����x�A4�5[�g��x �!��=,'r�̈́t}�e�t���[�B��3|A����w�V
?,:[B�����J�
v�j�R�:y>?Ĭ��f̧��7%WFP�c���F8�+s73����[Hr_�f��ڵ��߳���B�B&e��{�&���������q�><.C������u�����{��([�\cX�gcl�@�oP���r!���<�M=*$���Յ\�����/����'FǕ&!���Y�2V-E_���y�$�r���VM;�j�4̼a��,��␛�y�a,�/+���xQ�+���T�&���f(E�$����e�Ԗ�W ��~�Gµ�[�i�h7b��쟕K��P)�m�M@)�V>���`@�
��LDϚ��f�2
��F�XY�ZQ�Rd�@(S����u!����c���˗u�ၠ[;볳s�u��%?��W����hD]W��w��?��?��Je襩W�������چe�թ4�X�<u���0����Z��Q������������z���ɽ8:"�:L�0}�C�-$&��'�(4�S��Wh��q�39��KӀ �������5|'s=�,$G��c��yX�N�@��[L��!C���m�W�~_�OQ��؋�D[�\��1�
3�2Kh��Ǣ��c����~��[J$�A)k�4:>�D���T���'�i��}��آ��f�\�m�/��A�b[}>�&b9O��k馯���6M�7�,:����:�@a���]�,�L<?�A����F�<Et���q[&,AmZ�TTӌ}��^K;kr�C_d�sow��.>u9]�x^̊��8|B�:$V6�Qێ���3�Q���X����yך�׫>?h��'Ǝ����;a��W�x"؂tgk+�]
�ʂɑ�ܛ5�����Y�3�`���ǟ�9U��p���~3�ސ�V,�@Q_m@�Q�����-sr2F�|&J���2�	�+�9��g��-�� �u�sp� G�JGV���KW���r4~�ʕJ��_����K/}�K�l���*����'���������Z��Ag��}	��B��k��3�N���#i�}��>����W,xTJ�`�:c��F ��lTl�a�0q�á��&5�h�#'& ��c����G��@���u��k�f	�E�$=�cf�f$>2fa�ը�ˁ�ϐ�n��6D�3��ۂ��d�@N������R�";���a��DI�B���ѣD���>�ψy�p=�����h�E�9�Ahbir�ځe[H����\��i��\l�ʟƱ%ɼyy���x�p{d������� ,�L�E��ߦ�"��k��0%��a�EZ���<	���ܻh�H�K����Г}=;{!��;i��T+��sn�9���i��"��4�21*(���L�!�Q)��2�Ph|���b����D�cGj���C�����3~�	�e�{����~�9��w}+�.�0�dߢe���:�xs�,����h�3Nx�,9��H��AG�y���b�����wB�{l����2��p�x�?:�%W{t��V��,
!�;�M�lQ1��'��j/uӕ��dX$��G&�V+��o|�o�v�m����    IDAT��.��*��ﾙ?��?���W���P�3@C<Ԅ[XXV.���.�-�
�����-���<1�\%ۇ�TTU��0�[[�)��"�!Fx�+���Gs:,��؏\�4�ZSJI���0�͠��K���6�{�Z8v�c൱��h���X��VК�o�D�/c�����@v��92g(�CjXɐ��p����Vf��`�A���l2��KӇ?�ᴽ�#�x��p��(Ƹ�!& ֍ B �6���c9�a��#aOZe�P���ok��L��.25+:>��EKz�s�&��R�OQ�fQ��yѺ����y������}f�3t�c��gE�@�GsW�3�t�Ūo����)&=>P�Z�h�N�<vN�@�ד�3@�A�� �_f(�6���Y�9e��W�r_�c�¼FX@��*�A�3�w��̛�pD!cbm���ΧE��:���@�8��Oշ���ae��%�`�og�֋x^{PӮ(��JkXDɂ�XyB�ː]{�L��؜�üX[��Τ��ʹ�H��L�e��r��x�Mo�����_������<�@�{>����܏����P2!����~��U�" |d^׫
<thN���8�q}���t�)�Di���lmm3��,b�����y�P8(�xk��bM433-&�^6�E�7���Ղy���裏�#���N�6�>0��E}_Ҏ��֬ �B5g���=���0������9U$ߑ�dXt9�<yR�vi᪒u���$����ǎ�*B[^Z\��\�V�`Z�7�{|�
��9rȲ���_�H�<� �a&f+�����"~��|c��b�r����[+��2�"-"1s(
�"�hAc��1z~��f�������|��{ˌ�~BYc�n�Z_K̓�4=9�D������#���%�_��fV�Ϣ����h��i�:�?>�4��x�<}&Cl� �`q�4�uԽ��r�ʊ����$7����̹10�1EC����&�XC�w�>��g�>Z���`���(+S(]<�q���*�C�;���8]"|@�����Xӆ}x�A��5�q)D%w�E�Y��YEdz)
_��?��c:�xK��p]�iccK�e>�Ngcc{������M���W?vE����P������|�g�����ry��T$W���V7ғ�.�f+��z�'�N����
"˅�� �@�96��3ԇr?�^ >���P0"�959h��ʻã�(eH�y�����ٟ����5VB�����G7w�P���e&����� ʰ+�b(����E��z�f�^�"Le8�L�C����� ��8���GF�0.޳�ŷS�o��v��>������{�4/;{G���L�։�>����?�y�P�Ṭ�k�k�т�ր�f\��"�a{����iߌ�k�B�{�=M�����x_�iM�ڰ�xF^�5������V7׳&V�mQ�bg+=u�\������鴵���|��t�����V��xs��z��:4����t���SRJ�}>�N�p���`d���h8;�Gǣ�U�~��a���<b{wWK������� ӊ[�EzfK�6(��듭�P2��R�����2<N)�y�BTU����8��o�K�[����X	&��E��H����x�-`�9�� +JN�(Z�>�>����z衇�Qu<��o�1�z	����[k�}ego����˟�7����k�����{���ol4�����r���j�s�/�;���
�����,F���k�A,���������fK!�t9�̧�kH� ��$O0ǈ�A �� ���W��"�����A�o�q)��֙/���bx
�xD�S' H�R
����_�|Ɩ��jgFĽ8H�y�@���\���Ŵ�-����#�ê����z�io;2�9��k�H)�ʺ"�s�s�`���O��-̰�DѪ�&���ܭ�y��Y��p �!
;��N�B��v�DT�����5�1�ϸBC�Ӱ��c���6ڇ��2���9�5�t����2n���Z�E�M�)�J����\�?�}v�#�f�&��'���Zz����sO�嫋���к��E/'�
d���499���tSz�}I:|��Z{?��#J)���T�G�{9*i ����d���tV��C����r��	��arvXO��"���S�+m�μ�o�2�_��Y���͓?�CA���<��R.J���K=|��k��o�Z�E��{4>оk+�u`ĸJXaE�{\��/���2Ĝ9{ǏW��1��¢�t;��OL��yݏ���h�P�u��x`�����onn���l���L���+iyyU�\��q�-� ��M�?�3!��xB��:�!��	g���=[G��2u��A �0 D�� ��k�8��0����q�� �qo膤S���pp$Q.L�> ���-Wߏ!, 9Uk*����X�=���hE�����ȴ��z�i�#o	����J9kA����腤�ac��-�^�w�-�ܢb��8��p� �uu���F��"\b��)��В�[������BCzЋ��� �,j���x��W�`^��fd�h�\� �W:	�7M�0�^���5cf۷��ɘ֋#�I��L���Y�Vs?}�ݞ�F�ӧ>����{>�6��S&���s�>�j�Qq"��|%�k����+ҡ��ǭl��K����'�[ĚL�h�Z-��"�ߎ�u�`�fܗ�B'
{΂�u�ܸ�+&�_�β�<��L�o���t>O����y����+B�]�K�00���^Nh�]X�5	 ��r�BQ0�x_��DR���8s�/�A@�h��i��\��|P{i8�g�Dl������	���9�t:���x������U�T������τ �}��x�SO=��[������ҪV׶ӥ�W�a��F2�ٳgEX�O���>�EP=1�A��h����8�H���K[� j��%��"��P��?�ʳ�E��NJ%�q���A$����M2���#�f,���VZ���#�#���g�ߑ%�òK��泖�}9^��5�>X��w�ZA�@s�k��F@�<�9<�����&�	�]�,G�ܡ�~��\\Y�ȟv;�r˭�Pf梴%Axfkk�
���fXX|�>DЄ�k����E-�g޵p��}�dfM��5�����%S�"��Yӑ��� 3C[�����>��^���`�6s?CF@?��g����:�CpfR�XGj閛nJ/]H���'ӣ�<$�m�R��ե�t��B�b�%��c݃d���ӳ���ܒ�MUJk[�i|rJ������W�U�ܫ��,���u����d�k�h=噊p��K�q5ď!W[�V丯LӍ��
�aM��\g����"����ע�>EHCQ� �(��V, �E(+����]�;���^+D\��;pf�mp�m�g����\֢��ĺ!���X@��m�o����x���{��ɿ�h����u@����[�}�ޟ��X���k���Ԅsw����pIZbX.����̙3}��iqcȴ�և�������B|,:?`����c���ب���@=Ei��*@�VK���Y3�&<�7�B�o͉�ԴS���j��!,;D,F��������z�53QG�����~ZĐ���$��#�,�66ה+��-�S��TZ���I��(
i��@W�L�I�Kijr&>zDf?����s��Z� �'��Y�Kfߏ-">c�E��}���6{Xp��m?
 �y�����-x�
��`3�:�ɵc�@�U�������<����i3B��0s��;��{-����*����鳟����=8�Iiw{/�{�I11:S�F��g���X���ʮ�CG�'O��cG��Ҫ����O�.ǆ#׋*Ҭ��~D�!��
��5�!���� k����%���Vf�ʳ@6�mX��Rbh���/��,~�ݳ5�}%U�:m��O�[.�}mE�<��f���O(���\f
dz(�/dV�)*����2�n��4�Cٳ��=PR�����Ң� E�l,_�V+��=����K^���:1��@��{�}�����5:�����X0�t{C�ܹ�
H�!�f<>)�pl;l�!��j �!#�zsqҰ��/D���J������+TX@�y���i�5 ����8=9�{���Br*DLvQ�6~�3��h����+���L���� }Y�0?�@l��cMI���s�/���7��s�D��&� 2�	t&z�-��H�y�{ң=���R�faP�emY|}s#���j���Fu™��+���� �X7#� 8k����7�f~�[�>���,�X�3�e��̀,$��I�|ϐ����q[X���NU_[�e��n�;���!b��ڱe���p���t�o'c2'�ge)��,�{?�Y	�����YY�p�vz��E�-	�DyQd���3��������t�snMgo�%]�� e��ͷi�Q��'�R��ZD���9^w3R��1g|���sd�0L�E,��Y!�s�)��W�r3<��T����QH8�O3p�A�Y�!����|��$^�WA���V�P�-Y������\[�X��E���!�<��,�����!���d�
��
)�%`}C�gŮ�h��Í7�ث_���y睑s_ψ z�ON��]��e/^z]�Ի#�65��*����i��r?b�ONDÑ�kS�͠k�L�!Wd����#t�HP��xzWo��(��@����#���~�ƥg0��e�¿A�_C��P�>@9)���"��e�����׉�3Wi�{��kz�$����x�k�֒=7;��I(w��D�¯�D�!1A(�9U�����ieq)��}������c�j�z
���/�A�ZZYYKӳ�J^��n�z��c��,�D<.3M�KQH~���/ﳖ@Ƹm5Xq1�h����ׂ��-�YbQ�sk�~���h���u3B��l�0&�|������^+P�1��=����X,�mY
_N��������=�j���{�zM�+_���./��������r���Ո� ���x:}�l:}�������QP(]��&�x����k������@�������kt�b����v�W{=̀�-�|dDף,)�'W��?ǈn���N�`��x≾Eo��~)��@�N(�*�J5�V�/��Qh\�&n�Т`���P!(hhP-�Ȋi��DFx����'�ce�:��R��mm�~�k��_��7��3�Q��o���^�W��_��_��Ï�\��z���P����X�reA����M�t<����W��D���l�OL1ȄP[��`S�YY��G���6U��롁�=^$�*�Yh`ccQ=!4�`�n���-3�[��b��S����Z$�J�#L�M���w�̶��gjbv��H� ��>�F�%b�{2G�Yۦ2�quYZ#j[E����L�tNW.^Jz�e�V|�����{�~E����c��C�f�L}gg/UjUi��e#���G�������a��d�b����ck��a�f�Eh�hm���l�Kݖ�׉��J�%�^ v�i+�̢(�l�-9�է�D�o�}'���h��0@�N�ܑ\��̧�+���f������Ғ�]��ᴱ��{�Ѵxu5���T�4UB �t�ؑt��Ar��S����Ci����$md4�<}6�!KҶGj�!�B�U:궢f�
���z�ab�
� /zO8���@��|㹼oŖ5����=[Ԝ=�>e�]�S�,�VS�8k��D��xVt��C���"�3�&s��l�p�LV����wqm}��{G�%��\\���������v�������7�~�u��Vlψ ��go?��e�������J��,�m�>���1r��n���,Vh'Qm�5֬5�N��B������X2&e�ʲ���H��uձ�(��`D�β��
�< ^��W����<�> ��!���Rb'�1(�3WS��O���(�Ӈu�E�I�Y/;=�=Cp�� h(�-��H ʤHs��±#��Mg�����#M��9U1p���O�yX�����|��t�]wImR�^Q����P9���	���9Ճ#��V���f�s33�C��,Ru�xq3&[f�&��X{�|�-��W9�Њ �X��fE������5s3W	�\<�1���=+���d����������9[h�?��243=��[isc%]x�J�`݂.t����{?�.^�,�I��J��SJ��"�/9k�cSidb2S�jr*=rR�?|D��r���k/�W����2`Mm�*�,[��g����@��{�^�W*�HZ1�J�nМ#��3�+6قT�Jn]@�����Y��w?w� �x6ݗI:1{�І�}N�q�A�C[޶���0>"W�p3t����1ʒ\[�hW��mm=q���_}�k^��w�u�ZQP\���1t�}�y׻�󽛛����j�e�e5T"�luuMP��h#�9��,��.k�2yi�]���!��8�Y���������pLF���ҞSNy�aG?�<x.���
��ġ$ڋ*�6��a��[�8�fg4G, ��qPCh&	 �1��B���{ۺ��by��m	��2a�W�2��.,��?�6V�� ����JH~�ӟJ�s	|�B�W}�W��>��"r�����wPI��Si�y�@�d3}c�afj�/��D�U`m�(�̬M#j�\�<�Z�J�����K�3��ᛳuceư-�j��q[@��k���⿋�̖��-C�EeI��f��cfe����ur�7���Zu(�ڍ�����,���E%P�r<=������j��o���qE�?y<��N��P��If�S�ZK���4{�p:4LM#qnk.���P9�*Z���d��������mK�P6�+�'%][�Q-�8��㳯�p�����g�پH ;z�0~��9���:u
�A�f��C�̀���22+����t��s/���ߧ�E�|�4d���q�s�����ײ(���s��k���~������|�W��E���]��zɞ�����z��/��O?}y��{���J�:6)7�7��+�K��c���?)�#�S�����Y�9@��>] a�B��<5[�t�Յ�~��Q������42� �R!X08�g&g�����D�
��؍c�5�aA�l��
��I��A��ҕˑė���
�ފ��\k-_L�n���>p�p���������$�n)�][a����h:����ӟ���D3��O�Eb����Ï>��7���Ę>c�/~�����~�[ikwGi�S����ZU�������}B4�3cu0�
ma&��5C��kʶr��}\
�Z0�d� ?�QvEad��V�a��{�lu��֛UruG�!�*g~���k��*��~z[o��@6hڋ���UDjC+�L���?.�vmu5���%`����i}e=mon��7wh6��Ҋ~8U��� �n�6ұ'����z:y���Q�F~^4�r�/A0b^���2���|���zq�5�b����l�k]E�MN����AZ][N���B���r�DT��u�9���
Q����!���)�	o��h% �ADnS��yQ�ǰ�?sض�>��w,XY���({^���ʱט���t:[�z�Ͽ�_��_��_���3%�x����ֳ����{����^�7+M�cI�Ͷ`���M�5�P*���C�NGa�A]հJJn�hF�R����TdӢ_P0n1�^j��OpG������n�Q�GL�B[brB:����	p:�ʽ46<҇Hԛ� \;�z��5�p�Ü @�|c[���( ;����lo5����2����;�F�<����Xi�jsĘ}G�~X`����    IDAT�}'@Ҕ833���ΝKW�,(B̾�Q"��w��O<��:�T"�{���E/J'O��\.]���
�������*7Z�̍7�r:��޲�XSv���#��Cc��5�}���0~s�\m��ط�=Y���i�E�9�k;�����W��ueV�������!!4�PЉa9	���,[{>���L���d�頱�֖�������'{\{;R����͍4>:�v����3�����4��tl<�`�=�R�ܑ#izfN�;j�?�Tt�E� �PL3 9����l���@�CD�	�4�k"�t�rU� t����D�R��ֆ��@���p�ΌBK�9k���􈕕��O�p&�gO�Z�9��p��e	 .@ѿ:@�1��AC{��+�P�`V���{�LX��Y	�o��²��[�s)A��8a�O�y&����'t��줨t�Z�}itt��_������g��k��3f���~��������@co��C��,�h�
�lR;]]]VU�{�Ve��7�|6��SYf��������xo��M'��|�-�dD����!m���%�RyC]�*Fd�OE�91���26=IFF�et� 'B�I�ڑ�ȵ0A���T�D ����T���Q7�>�]3:�W+\TӮ��F@�І��7�+0J�ǧ��r�e��ʊ�����~@"�J9MM��ť�
͆�q����w�;�#4áZ�ru!]]^N�[[
<���N[ۻ��/��N���$h�`�{��d-��5��%h+��?�CXX(�Gd��u��3��4Ğ:��}Fh ��Qffb29����Y�o��6��=a�m��;�P|���S�4Jf��.C���='�+�
������tu�r�������҃��_V̓Z��'�h���<�n���:��:$nׇ�����ɉ42:�Ν�HA,#�.L<�0zO�wA@4\$�:H!����+��P�����Xv��b�����f�������7�R�[%Q���=�4� 3Z�0�i��g$��@hR�-5"ꍂpX?Q�$L���JcQ�_�xA�,��@
��� 2�3�K����a�1��pznV�"��py���O?s����w��/����FM�g���
�s����w��+W�8T�=��lW�G&�I�a-o��K����Zb=��l5�6��r�]"ȉ����6�Llε��1|��� �-"�(�፵`��2BU�s^�p]̔N����B^1�Z�f�߃�[�`-	��|=A5� p���_;�+bc1:�f��y�0�r9���嬦q�/�Hx������v���_Ў<���������u��Ç��p=��� 6D�G����������464���鴷�HG�MG��:��h&�o��~�k_���lI03rC�H�C@�b7&����}���Զ"-lЈ_!4���)���Zr�� �5ͳlY�r?��>�K���P,"��ϙ/C�|�m�=Ӱ!H�g��>��YJ�A#���(�ϖ���/�./�����CigsK�~?�O�7�
`�*#�i|zZ��"��jmX�*�wQ�X�h���
�[�3Ӷ�hK�N�ZP�JVD�d��)>��9���4��ŕ�5���E�-�	p�>w���X#��-JC�(��P($�
z;8�n��@m�v�B����ǲ�*��n����˳�A��<˼�0� ��r�~c��cRZ(�J�����G�/W������z�W���_���=r���gT �T`�O|�3o�uZ�xpК������BW6��)nwnn&ݐ{�ܓ	��j���Uf��x@ֈ������l%g���?Ƥ9Lq臅�/)(�8:1�F	)�!!2�?��\�z(r���m�9�2�sS���\~����V4-�~>2	�k���s=���q]=�k�����9���d��^��r���BD�֥EI�Q�t���4\�ڋJ�j�ґV6\W���/(�2&�Fk[J���%��MF8�!�/�CQX�'�݊{f_���!�UdK���w1K��{ô,`���;��:0w[�|���q�N|��U��/*C�I��<q`#k����jk�
�AR4
շy��K�.�cub%­���>����a��]�����7R�2��j7@�F��)::=8�OϤ�q)�($�r&P6X7��f�8ι�bd]`ƶ�x�������r�P�S�<X0�������ˋK��"ZD=������y3�m��)$����,q�m>ӭ���{��XK��J�����Z��9U��r��A�f!g4���=��;"`������5ڽ��t��;#������pN/U���z�7|�[^�W\�oZ =p�=��g���;����+�Rꖕk��ۊ�YX�lD�٢���ʽ��h�-�0��0e�lJ0.o�ӄ�.��y��niS|��kB3S����8X���QI�ѱ4>5-�z��G�P���#�zQ�@��B7��u��s+ڡ,�jE�c��w��d��P�we��4�[M.��h�E$/��no��)<gn&�� ��<�����*��k5uO3�z���<����>��{�i,k| �s��t���M�B0�6�`@;g���51�b�}(}�!A�y�-p`N���A�:����a��a�n��u޻��D/��k��r���>z.���y�{�ŵ�0���A��k�cx��,��m��`�+����JZ\\��Bd"�������:w>]Y���j���b?��sn�=�O�	B��ʙ;> ���N�0|[��cC��mQ"%�G:�CnG�6�g��N��i6�~
L��kE�X)Kz>�
����rL����g�^� ���þ�����@�մ���cWG�C��x�������$�Q�j�tm�ee��i��}�!9�B���B�����Ƌq�g��(�xymU9{��?[��n���?�]������/�n�O?�`{�- ��~�~�+._8��J���Vw?�zua1-,-�� ��"�`~>�t�A5��oEcG�.p(I@s���gAe��`6	m���uB�:��6PDQ�.��<�:��|1<F$Gx)�����a
�>�|"(��Sה�z�����T
��}@�i:�GɌ�����V���N8ks4 H��}Y�Z� O��K���Q������]ѧefJ��:CPQ����Z.�PlL>,�L����~��tT�hn���[P^�6َY��\Yx�N���~��
`[$�s ��l!�A�!7�C�e��w-��v�>�);���;��[�P<"x�BQ���3�ql�S]�Qr�Р��]�i)e9���0E���ڀ�|uuY�k�+�/G:D+*��ѣ\�V���9�I�&B��1�b�5���m(
����?4G�26�[>>��Y�(ه�{1���s���;�Hy큔����}�8;�ee�a�"��3����*�/��v�2����^�X�*RT4�^���=�]�z���'�,|�En�����<��^]ZV�i�J�W;��>u��)I�6gpkc{�w}�~��o~�}�OH\���q�d~���z���뺝η�+��bd�GEօ�%1^��*;囹�D���Im�&�W�k�y��(�`�3kEm(N8��V�8�=�C+S���PtI�������^�4���� �~�W�27��)|Ea�eq�{�en��C1-��:"����	˺��(�ҲCT!�A2��A��\e�yȗ���"�vx���Y���!��^\��������,kdH/ɧ~�g`�F��$�D*̈��m��u#R�V��������4�M^3CC���s�:a�D�j�(İ���Z`�}�����{��s� Cl<��m�K[����6yO_y��p��P����?��f��a�"�lQ��di�Vџ�s�s�e"*o�F�O.�����#�Fc.I�HT!(�cdl�,���#�ni�,i Z��ܜ��}��/W+"Θ�����L�>Z��3�6����������Rȓ�ނ�X����{ƺ�DT�a�,|���V:��|���
-���^K�V��a](]41ն���{#Q���4d�辢E)��Nf�B�q݅'�	u�2f�Υ$�5y��9�9Y�ʡ��������_��g~�_O��7����|��;������������T5Iy���\���.-E�i�p�?�;<?��S`��@��یf���qQ������Ђ@��Q?h�>�m�	�;�@�JUa��軡�áU�q4M���9$��xB�)�6G�):fr�_a��˳Z��ϹN��bi#��p҆���+4� =r0�)��&t9/\d�Ky����� Q��6��I{[�j�g
n�Sv�Ֆo��E�#̍p]��86��f���s���A�s�,<x�5R�faŚ�}�L��˫�_�H:[AbT� s��S�H:֒�Lc�4lU���w1�4i�`�
fg��g���S����%[���h�yXPRn��,e�� h=`�E1'4e�͘�g�S���HX3��uAm2u���a?;Vۡ�C��M]ǑZ�y�N��ι#
�ya��<��$an,ȵ�9ʋ�#���^����ezb�F�D�jX���-�
�ӝ����E�W+z���ה*
����TQ��ZX`��ī���᱀��'J�� �=0���J^��Ζ����J�K������HN՞U��j�~��ٟz�?�{���7ˆgE Q��~嗾������^��CCCc�k∄Ѡil�3CCiw��Te淓2	���$4��	�u�����|.�S�Cv���0�`�^h)�PT��K��zQ<U0V%����֚�v��j\��>�
���O�`n��p���pAxXfv>� Ja~�$n]k�ٌ��L��>�'�i�G�����,d̰�3�@��Y����t��#��Z*�zr�ѕ��b�k�*�X@�������v����z��ٰ�Ckg�Ѕ����~�+�9b��s�=y�i��i��Z�b�`�2T�>��3C�,�����%�l_�å�����#����a���nK���N�ж&���������)7Ux>+����mqⴶ"�vRDt�:�^Qe�j����Qn��,����Z����R}$��Uȹdܛ�;�ڿ�|/Ci���eMX{W��Z`�0�<4C�C�cj�����V��G�����M���8o`�D������h-�kr�t]A Y����o����{V,�cD0����#���,��Ҏ 2�?���~!��Py��n��7|�7����?�l#ϊ b�o�ۏ��G��/���++��	�Z)_�����t��i#�,�����g�U[C'�/M}�l�"(�}Y�COe���=ݨ�U�k�^ M91�u������g��g�vt\%J�Gd\%jn��OXh��8�<_~��1Y�x.Q@��		�h���Z~��E�>�I[bDQ��@�8��Qr�!83{<C:ۛ[�`O�a���ȖQR��reW"`ޑ#5��gg�2�=m)���ܘ���8H���f�|�k��2�cxΎZ�f/�T�`��L��!=��GxQ[C|n+D�d�a��0"��s�������w�������#���~����Sg�\G2��-�#�u�Y�ّ/�ъ��udlX�L9�ձ3r~#��q�9�FBw?�h	bR-�����p�a�9ֈ1��5f,�c#K�C�rn}=�m �,�t;6���S�2�fL�Ie�܁^[>cL���9E ��O^�o勦� ��㾯xA��gg�\<�m�-�xv��h"�u�zRXX�Kwqy5�O
���禦����?������^��J }���w���k+oL�Η�J����㓊[^YV	�5�Ç�(��k!���	�Ֆ��LXD�	���(�$��=�H���,d�	�+ఊ0�f�ĳ��F��a1���8re!�H:G4�6��w�|s'*��9�����	�haPJ����f�Ta�C�s-z�q_�-S�����S���gf�X@�X���Ef�c��b��-�h1"�"�0�tf�[�7���0L0������~�>g^�3���*����E́�|���B"JX�L��p_���f��>	���~��e�5u�a�Љ����H�8����l�b�����YVs� �u�q��B�-�(Bٷ��7�J�i�@��#B(V*�X+����0&�����4�[��f��}D:�����
2�7�5n���(u G+:��r����D�P�A�p�6�c�g���J�נ��^�*�#�}���s�-Zӝ��wl�P�al|$�7�er �abK���آ�@�p��5��2��J�{Z�{����o�C��SH>%�5j�����'n�����W��?Z*���3(��5�9��-�|�G}S����J��4L5����T���B�	��̬j���G�5G����ڤ;��}1�ޠD�4��� F87�ř�B9�Lڍ�����L��u-�H'%J��[�QZ��s�l顤�J���h _�A���ဍ9G"��1��	���!��ʃd��ɻ�� BY��C��_�u�!���7���[cmͶ�dA�������qF�?�������p�2���w�]���g���K0��}�]h�}eMXסjvF�Zn�[I^����g(40��s�a�:dN��0\��w�n�v0��5�h7�^NEan���,�����tZ��P
[�׺#��q^�@�#k)'M�RR ���~M��P�;p�RI��\���\�� ki(��D�FH��H[���?�V�����L�j�ʊ�J9�!ha�sh�b�[c�T���˳�O:�a}[)��??�3����pTg< %�S�CQ��Bq���������O�]�{��"\�~@i3�g�T>8{�fY<��m �}t:��J�����k_����z��9O{Գ*����w�/��k���k���
:�G)�0&���j�eT���D�����c�������W8�y ������ۅBMHT�CM6�"դ�/��b�G�H���P��%��b��s���*�8�ժ4oJ�p��~B�@'���BF��r؂�&�2JFQ�?�!ub�����7��ָ�E�1@��;���rI9���}��0��=�+D�H�x.;$���D�傱��ns�{��,�l5!�<^���~'p}���4�4�ým9H�!�:��`����� �Ƹ�.'F�d�i|���!?���y��غ���5���[L��[��Ȑ<���i���}a�׮�!K)����c'�#��hm�<1�N�C���?:���`�8܃���H7�!^3�s�he͟��X�
z����-�QzF�|.�A�=����h����n+�ŝ�Y7[z$�f���#lY׃���Nnw�8m�y�����'>���:C��d +�=��$I��%(��v3�~ԗ�wx�%��ly��V��<*r��!<�h��+���;�S���霖"hgww���'O��w}�+����p��KDi����_�ڵ��o��k_I*���Kb_�rU�C?k!�k?y&��M��h�"R?Y �ɡ�v�Fwh�\a�Ձ�mX�ߔ�a��v�{C	� @���C��NP��R�@vu�ʲ�t�c\�	���g����5����;���&(x ��U!, k���r/B�@��g���v
`|�Ku�Z-%�ڗ`x��!����<�a8̛g�q�4� ��%8U(l���Wc���z9��L�g*o$�T�3��>��ͤ��lb[	\�sG��|x9 �kl	�Q�c湌�0���X�A�V@���'�~?�4366чD�!3w��pi+EK�̌zp}"+@�]
uf��{�%"���W���K����_<�U3V���t�|�b�����YG�B���֟�s��Vd�u�����P�\��j���������q�{=��,���He����fDt����!D!�sr�,c�O2�E��Br    IDAT��|��+�5�O�f�j�L�M��2Υi���n���e�	+����ކ'P��`!�z�:�(��M�W���n����_�ܟxӛ^o�T
��Yx=��}��~��g>��n5�_^���1A�S3���W"�>���􄠈������F�1� w��%\�{����v���<�^aSww�_]���&fip^� �U���A��pqPԂ��Q�D�3G�Qt3�����@�X��Q�h���94�sB���"�gP�;׌"_Ț6ױ&��3��6����F�4���vB.�Mr�f�cCLQp_K����t�ݡ镢�H��� ��[�8�I�_&����6��`?�a2>�
�Y���ɼ8���>�]�K.�h����ʈ-��#��q=ϑ�\g��u,��ۗ'�*[�́u��kV����P�h4�w����}������n:0c�/�1#,�k^t��3`��@T���S+E[�HT�K�sGc���
��{�+Fx��Ĕ�!U���O�&�(�7��1�r���'|�?*X�N�=��,�L����Q���ؔ 3t泴�؇���a�oȏ���ʸ\c`���� Pµ�ju�7"{��YQL9B���֗7�[���1v:�Zx�ZC�i���(�:_�梲{OT#�S�
�Q~������[_��/��t�keܳ.�x��������.��V��Y�׆ \���*Q {��
���� fg��M7ݘff��.8��*iKPX�VvwF��2�������������L`�ƚ�
�D@��O����(���)4� ���3�]1��� �T~����d�L��8M$^�r�Rk�v��<W$���F���Xa�@�nX�����������@ �<k�EV��H8G�|P3f�Fz�(!�cp}()�-zkc�"6b>�g������b���'����Pb��y������?a�\�hA�C2,���g���a���eOTe"7L�\�����(�v�sO��^�w2��׺��>*��Ġ
9q9,	�m����vޓ`��Qy ����Ǡ<��nT��٬�=�P*xQP��V�:���lq��ʚ��dX�<:����AO�MB27������,��n�}��	aea�k�� ��RT�^�7U�.Օ�������~^C� -7��V��|��9лQ�7��%dskrӀ��;;[X�|o+���c"]���7��R���Yj�gKK+R@���˕f���ęSg~꛿�?r��w��~�^Ϻ b޿��z߃���N��GGG�p�� ���-���J���^K�
7�|c:vt&�RK�@&FVD�Â�,��q��@s@]�h�*,�8�++k��3Gw����b]Dą�&&x�G�Y�9p(�[�Z������$� \�Y�&�sင�.�\s�� �诂Փ+���Ag?�5cԴ�*�����Q)�l�-A�Iԛ��YC[(������a�yU!��7k�\P.�MJ8�5�A�4)r�sG��T���(����+�.&kJ{-�naA]OKeˇ��s��.��T�2�!3fC&���ߖ�!3�.�{qo��a�p`����������ϲu
���j��(k\<e+z�}�����h�A�5~��!VڤP�6,���LO�o�_��R�N�7����5�jo�dֵ͘�֜��L/�߰�%|V.�}CT9_]^�χ}�iP�]�Ky��M�E������7ί�K�O��&�xX(Ed��IT�0⢾D�OS�Պ���e�@& i���2gC��G�oDeV�}L�
檞b�����M��5E��R*�����?��7���gI���wB ����>����W��*?���uc��	���|eaIY׵�h:�ǂ����t�̑419��!:���3Ж��~�[�j���ԥ=���p`�,B�uvttc� 
��2�d8�`��V��"Iw��b�!����r�l吘'f�#���{�@k==�A�P��V��-ƥ!b}FE�\=W�[��q����=|D�� �"@��C�C24f���}fX����(�7̃��k[�~6pk�6�ߔ2!O�	��5�c'UXc�N���PN����?���!x�J�5�ä́�Pkš��݂��(ӕ������B��΂�=6��3���=���73�笠<۹3f�̷�s�Dd^b����2�y��0̓�N.Y���(>��(�ϙsX��\�d��u�di�AF,(*jHN��a�N~�מX)��b8��0����i��]�������|ùX��7f~dAJf�z��U�H�1�]!9�B�Rr�>'�{�(�Vz����Ͱ(��YlEkր����.�7>��SU�ߍZ����bFF��:���W|�|˷�d��@)�|���}��wmoo�������&��R����FZ����p���.�n�g$�|��t��Qu6d�1�!P�;u�r�"vd�g�����ELW#�q�Ics3�� {ISi˲��dI#�������U!����˙��fE;jE!��O0�3����Wh:0%��FT ������A����0B6��2�j�L_����,.�9��6ȩb�X=}�3��PX��7Lð������G�+�˄R�)��b�́�1�{;���zis}S�'���q�EXP��0�b�B�#"�}��֚��K�lo�;�+ףU�ѻ����u�.�3�����ks�Ge�ps�5�\11�������|'CG�V�,t�'E����c��}�|��"c<І��恢T)�%�i$��v±�uV��aAuTq���{!���@�7�¸���$2�m�"�� 4,�@C����VV��A3�=��u@����PX0�<8����PJ"j���UXytT��l��ދ���P`~��.��K�g$kN��ϋ58u���Y[��[F:��{i����m����?��?��R�{�$��	����w~��>��������J���P��-���zZZ]��TM�.���Μ9�N�:�*�������$�H{�8|�����@r]���
M(Zl�7�:�e⁍pF�P9!���7� �C���щ>֎��,��p]QaX|@��N�>j�'|D���뛩MQ���Ό�N�!g�c� I�QjDI��D+p ���e���R�r�W�Ҁ�	k���|(�R�gˇm�L�V$>��`F)h.%����+��p,s�a&�JX�>�<���+j��F�Q�"y�i��~`�EM6�ܹO�{d����։���>������� �\�SPP�	Y�J g�ʘy!�l�@�
���r�p�U�G���2~���9f(V�^K�ˑ0~��)���˗��`�:�|�����_�&�n�u�ڍ)`',J	���8�b��ZL�~ Y4�}��51\Hc>�����7|��=Z�-��F	��7���*�9J-,x��!��iѼ�{���ס,��$Ou������n�gxAL��͵��y�_�%���|�$�W�F'Ry�|aye�������W^��_~�d���wF �s�=#�{�{��X]��V���T�9�|��݆�4�l7R/U���͎��'�����"Q_�'�ڇ(��8������F��044|@����B�R�#�h����Ю""~�?<P^Ԉ�#\�ϝȊ�4>>���^�(B��c� ��G�'FL� ���β��-f�]����Qg��B��,���������j/2No�B^΍�`)j�0��e���ETG��I�{����tZ\Z��Є��`���}�~�wb�5����rH�ek1�;h^�u���$�j�d?������Ck|?��x?rNvs�3� �`4�c�������B(:����k��!P)#YIaޞ/s�"�9��Ba��������'׳��$�ѹC��+�%k`O��Ë������1	�̂��Eu(��Y��^���c��C�r@� )�ٟ>����h����7���,�|��v��9'�IrҜ��$`�V���BI)����Q(�Z�Vas)W���b�J	W)�����@	J4ҥ�s���v���=���5O
���$Yc��^k�9����{��}���wG�������GA�/�HzV$�s9^w���̼ţ�<*p��?���ʾ�2��r,3����^����J��+��B�Gq�lvn�������۷��~�c^x�Y)_��)����?��^��O}�?��[߻����b,wm�!�'OT����66���L��^�w߮���U09Bcmy���t�-�K� ���Ū%����G���"���6ގ?d ���$��\dK���MP}r�E�Rw�� �8E��dp.	�z]I<;�O���N��/���9Y���ιVx҈a���k�t%�̪x����iZu�%�Z ��g�c����K���<!�X_
>�XF<��\S�
�T1�3�G�9����Q6�����*ǈ��k�0b�3�&��j�mRI���x�^8o�n<�(��W��E �ۊ��|F�1AG����>���$��@?a�q�-�|A��ȫ��s�N��tj"��Ao��Ih�\SϿ�d���+t~�?�^8>ժIi���+	������,���׉����6�b`���]����E�K� �3�.$k�:^O��T.���+ø����۱FmY��?k��^�es��$a��vA���?X�Ryt����5?��?�[/y�K��������o��g�߳�������+(�Rv�^A��������3Pg�.8 (��.�[ƈ�X�Y�5Yo���Sù'��� ��͌�/�*��i+,AeC3�Z�e���QTxN�3X��b#EH$Xl���4r48_�&63}�;�X�~JEY�V�r68��j�s�܌�z'&6j�g�K�t�919c聛2�]�,c����(*�z�����Ff�,-`�5���0�B����9x?�-���2gM!arA,զ��b��'%xbp0��g�N�)%&���9S�/tn�
l�\!4�^��yNy(�xG�lИ�Q{����XI��/����+�x&׋��+�=k����H�2sC/�F�y�}3(%�7J��B!3-B��e�H�TΙ"x��oH�g$X��k�dĸ�;��\���G��-�k9U�UZ���5���a���ްq!���(���<P�-���fDn�ISD�)t�$�B�~*,��C^Y�W(���۵�DL��ע� 1k����jzzj�ر��8�+?�3?��S����<U4a������_X^���Ņ���,�f��U=������U5�U�q�1U�%xN9b�]j)��/\�axRx@y���|�t��Y�(���]mS)����ѹ��]��ڮLftUMOQ���l|&�P �6�z�ka����1��W�+5�(���j��J��6����W��� �amź$X�k�ԭYj%�X��\4�����4Ђ-$A�e�ϓ�K0��^W���T-x���<�w� ฦ��D�F8EQ$�ż�`>�
#����0�b��3�}	�-,J��e�3dL|��}�J6�s=^����8C"k$�'s��-E�1�6q�/8���:�n:=���f���Ro"���b���WnҤI�,�]�����圸{"��b_�t0�o����Q�Ā��_�b��`br�f�t�[��u't���J�'b�6D]�41��b�Ɛ��Ø14�F#�L�y<��O|[���)�ZSq��y�=w��y�袋T��uFed�ք!�CG�{��^��_}�K_z�$�O9�����3�s�_���Օ��t[�"`�^����^���^W�-7�.�iL��];�?�����NrQ�]�
��6ژ���}f�%��4�3>�V[�&:x��J�(�Ra��\T,L� 
�\,�x@ސf� ZP��hZ*̚�y��)���Ѵ�+�'�Cl)��@�ly�*��)�TJ�`m��c�|7pg��L�2v���p.�K�R�2�?+���71�)f*xNX��)dʽ���OL$�q�&<x$���7�������}����n��A�����{'�Cj�3�ё�oB�MO�s���ښP;��lX��vi��*�SZ!*>5fF�&��9>c��6a�dL���W�a�-/�։�5=,x�[�4�+����L̆�n�Pb/y�yyVb�=�ۜ�������5s&Ϥ��g�C�xO�sHQo9��=#�i���d��8�o!4-D�G|?4���A�2&����1b2�I�Q�v��Z^�<��o����?5==��W�����+�_�y�r
�yy����7�S??6޽�·y��1�z��?X��o8`�,̎�{���%�%_5A`}�Z`2Y]bB�����rz, ����Yj�%�^e=D���cda�A��%T��A��U'�1ɚ�ɊY�2#%.�X�[2�ci/o;�
lbQ(+Y�%������a��Pi��&�&��6�'���&|������97#|ZY�[��"Tc�s�x`�ٔfp����T@�|��&�oM՘Ǻ���rhƣ�B��n�%
3s��E~H�J�ň���#��
�+p���x��\⹱�2��S�lr�2��߄�2�l�e0��c�R�W���d_&�,���d���c\�c�<{�;��q^T:К*�Ѽ���Q����;�s~�]��'�|�p,Ͼo�2U���?�4�^��O�Uk������Mp�O�ɋ�j��e�|?�d}c�5�|�D��Z^?yV1P)�8�3a�`�}C>ˑ8�瞫���(�V�sx||�=�_~����u����;#yy���\����{����p���n�
`.�!Aq������֥�����=���ZHgDn� �2a�.�-�J�����|Pӌ�C77�9X'�	7-�bA1$B\L�;�*��xO��	\p������* �Ʃ�_���!�ټsS�tn�@R�Zw��qP��W���;Zq�Z�^�Gb�yN��v[,g�v9���������K^q���ʊ@O|+V��0yTf�����R0�M��SXH�cyN�'^NSx�S��iB]|'�/�j�Y��n����s?�G������F@�w�g�@��EYE�s�-����o[������K��jz}��x��������t`� 复�9�9�f��y��k���i�6�J~m�5��ƎeOm��*��%�:���!�@盥�+�Nn��X�����G��=���l���D"��}3cG���/���	l��̼�Z��iw:�P�������$sT�Ի�-k)$���/�/�y@��s�&cܹc��7�#%y��n��9_ZZ�����w�?�y�������q��S�uJz@����.���[v����Vk�S�p���<,�CG���"=�qbAg�ۧ`\P�!�b������S�N��
-�RM;�绱�ϟp�eC+��)�z������?���cVM����&+J/.��f��Ĳ��+�Ŧ�Eb�ݹ�9+��d�!
����T�K!H,��DV��bʒ���ͼmH-��H�"�cu�~��2�gD��W7bBq]��k�9�2�"
(�`���ce�Gp�w�f��o�Wj�Ei��@q�(�^0�^W��(,+e��;ȸ��8�IC�Z�H͜����������V���R�]O�E�D���'��\�1rl���-�����r�a��(a�=R�R֥�B��i�jXr�`]J���Si���aO���Z(ہ[��lYY�XbF����E���4�M��T]we�=�s+�xa��w�j�!�TiB��!�(�N������m²Yk\�g�=_u�Uխ�~�z���'&`<8��E�+��;�6�<C�@�nll���O|���?�5i���t�)��n��}��{�_��������������+�Wtn���u: �����(xؗ\rIu����*��dh��֮���4��B	^�T@MAk��Zg�Br�K�C��4�l�f̬�8    IDAT���ui)��K�@l(���ǜ� r�Wt"�G���	��%���$���rg܂�
Y�y�K��� ᜱ�Q@�&�E���,0�CC�2���Ɔ�ѐ6�Ԋ��yt�=Ǻ�	�>E/c�g��O"i�z�� ��'Vb#�40d<�Ĳ�WSh�;w���}K��	�2�I2����K�-���Q�5_�8�c+3�c,��x�( �%�2O!��Q��L�}Bb������A��Z���R��*����"��fHJ�0ޭ3ɞ��1Pd��͊�L״6���T��T4qo����G��y�j;fH�s �9��r�6c0/N�5d�9��H0`�E��m���<���p8l�(�<�TP�2K�쳔�ʽpmH O{��$#>��n��&����!�����qҌ J@����9l��A���b5�����}������WR_��OY�d�����+����2>1��յ�]*m�� �C���8�X�MYD�,�o��oԃPB�*����b���˱�~��P!H�(��f�:l^6!�Y-��*�%\?��|�2[U�i���%b����}��h]�cG�SIFc"@6X��U�S�l�m[l�&jZ��='�eCn��%�Ƣ$<:�s������$��l`�(�4^!ǣH��K��K��w:K<�_I�ܵk�h)����lQ@�����"�%4�Z������s�=�}����%r,�//���9S 4�1��(��ܚ��}���wp��-�����X���[M*�b�"HL����-�_6��YgOA�I`��C^aޗ�O�i	ϡIZ{�nz��M�͊����$�b�f-%{��2'4Jd��Fh�l�0��4�ٗM�����<kb>��k�q#�&lc�
(�wvv�4�t�B�B���Q�dro�W�,�8���)L^��)��1�nY�W^ye�{��{ս�ޭ����<|˷|�������5d�n�O������W>�~���g��嫹�)�����w���G>����?�j�.SYJ����#�����j�d����z�%�
�
��B`����Ud�B���R� n�ܜ7�[[ʴ�=&�5
#O,O[ke��:�q��B$@a�z��:�c���#Q@S���r[^�]V��~�Ӌu7����"��i#�L��\�@�N��#���[rޕ�C��$k6��(�XűL#851#����v���OEem�	��
��o>��e�̵�x���(hj��V�1&�Q�s�#7��l&˼@qQ(����ʁcC��yVbQQ^M�( �	��ϋ�q�d�@�#1��uw���1"�L�k����Qw<����j|�y�mk�db~U�AuƜ��栰(�,T͠(ڙ9zY�i��Z:�iqn%�.�BMY�WW\\4��
�'$��7�C��ۘ�cR1�{b�Q�R���T`K<2�{��n[R*��J��(��k*4t<+�RM�S*�&m<6�Ml����(:+��'<�	���r�m.�5R�����ϯ��������E/��S�����j����~���s_����MO�����!T���~�զ_�3���z���L�u_�uu�47����d��?�h�Ј����&�"BSh5a*a��.w��	X��l=!~˭��r) �#�M��p��4��Q@s�����R>�����Yc����HXV�jya��w�Y��9�>?��K���_Z4G����⚔�O|�k*�YB](���#G�]�wjr�W����&�!O�B�F�����P��욚q�������Y��]�����T�:��ToUb?��F �&�c����+�#�Ϙ��R�넌@e ^1
8 ��,��ԹK,��&c����TT�Ԇ˳����Qx@p�#�1~�J����B�?�%��&�����T�)�1W�槙oeRYx=����	�C졽�c<~.%��W14%9qR���c ��#�B·`Oɢ�p�!4���\��>/
�5��Luv�J�V@ca���%GP]�J�+�J,��E��q@����'��n�M��9y6V8 ����ÂJ�Q:~�ytrr���\����_y��|̈́�Wq�S�b��_�����{��jb{ؿl8�y8I���nU����xP�k�����.�Lt�$����,0�!ի��c2tK��I��B��!��-����ݸ�����d�@�{��v�|��
�������rB�{�S��@���@�ءD�`��.8��-���9�4y m�x�BaC���/%PP@|�{I!K)����Ԥ�J��T)r��*�w]m�i,�mu��ǫ��jv�g!((��(��'sa�xO���y��隍ܢt����r�4�f^٬�ӴMv��s3帜q�,�P�G��0&�du��	K�ss��x��W �� �(��x.��Fk���k�N���ⱅ��8���S��x���J��#ǎi����M���9���u'�&��Y0F	�ށg��W�=�eC�44-��=ƕ�J����1:[��9�uʚ��Ԋc,Y?���&��&��r��qbs�jSe�Q�5�g�ۖ��s3����Өƛ��s��j�yb|����1WI���c�NLb4p/�5�`<$�;���������SSS���׼�ڧ<�)���sZx@�������^;66�����>��a���}6K�	��p�d_u��^�X�\���^M�D�Ҳ@����YД��,��yV��Vg�p�a�Iec%�^^P<{B��Q�l~ܥ����+�C����8Obvf�����{��̾�**ֱx��)̓�I�:BV�Oa]�~B�B/�7���Qi��bʆ�e.(�wT�d.�E��DA#�����9�5猐����$�b���#��7��K��y��)��Z�(��@�M�bue|y��^]�(�;p��{t�e}q�e����HC's���U���$�*����!S�oW�k��$s���F��<�SݸM���X+�+�Q*r��SoY�g�"��+Xg`�<��4�C��4,�L<wl'YӸ�����i�l���)#{����G�q:f��r�72�������vMǩ	��"_���a�����*�7X{�C:�V�A�}O�x���^h�k��5ʇ���Ҽ�I�p��ᕕ����'���^��/~N����S�bvn�ᆝ����_����c�N��[�VO�Uo��OH�R���5B�����:��T&���±Kn�l�Y(ڱRk+F�ΐ	P/b�|���AY	�B�y���_�v��u�h0��t>���7�#ܰ �#��ߪ�ݻwU3�a�ݘ�}�H�m	؞c+�+��&9�@[�ϡ��vc�5f���4��UKC�.�'�Q�E��w��,����bL���rL�/�B��;
��e�k'�K�<�e|'�Jϯa-j�5l%��L�L�)ǂFM�b�Ȣ+t�3
���r���/��Tp�x)�"���#�LW�fY�k��y睇�)+8�c��$?��5��b�	b�l���K����9��W�%�!o"
��RJ'0'��o~� `.���o�Cσ�h�7�P�����$KmE�U�{2�UC�^/���^�l�5cS6��MrB_�Zz���3cN��1g#�[�"TR�Ɣ�O��^�AY�kC����5�"ɼ��ko�ۂ�a�RΞ�^H8~�ENЉ��5����5;;����7>�����S1����P@����>��7�d�������~m��S�MN)�b���P^
�(r��W;w�a�LP�'����)��'���FX0�I`��גk�b���+#B�b�@V(
mށ�"����L|n��:�-~ $~�wD�k90?=i�:�N��#/�Na�t|�ބ-��F@paߤ*Aʪ�r߂7��^d[m���3o`���b	V"��4����Y:��bmZ��_,�-�&�-����/�G�&f�5
�k�|�)ϓy��(�\�q��{����x1���󙜬���~iS.c�@����{/�:�>53S�x�g�?�BYC�ϕ|>�z( �#Vg��W7�5�θ�<�$R�*Sܴ@TM%K{ƞ�\P<Ʋ��\�@�R��w[��}�����j�L�C�tF�1^�N�\�:��8P�=�����cf����V�c5��!!�>u�w�5e;h@�����lD٫4!� x>(!�M}C�1:�5������0>>��������g��5��ڷ�~���R��6
��[���?����p8����K�Q<��1'j��a� @���?Wns}�Uza�5�E(�G���sJ2a,��x�x��������e%�K�7\<As��X"h2��j��I�J����/����O|�ށ�AS3��Wg+�~�]�&��l
�Zq7�(�'��mZ`����B��{��-�O�s��c�e���z��$c�s���<��A�Qufƈ��,����� �	��Q#���ł3�20^Ss��&�"Iy��;��1�x�z(�u�Z�}�5c_Xr�Ԯݻuo����1v����2&�2J�m��"c�Q���X�Q�1�8cӳꏒ�#p�1�u�g���Oo�(r4����St��^�Sy�U�-=����f��7��g�#*����ڥ�X�Ȅ��L�s��Oz+w8��oƉ��� ��|J_��6(RC�seDѢL{� '���x��B8N��Jye���7���7|��}�߾�/X�j�����F1Qo�������?��?���~���nq�z�]w8�c�mX,�s�?�=K*Tc]iq�m��S�;$ڢ1����f�E�s����)^�1Г�r�7)�9W��X���32�{�^H���K)���1ſP@��֚ ���	���qL��x�gB@��2�x��6���K�z(+�QDX���qw);Ju�D���*Ȟ��<�x{��F�g��C�p@zU�8	��7B�c�n��x@R���(2���+q,c�G�wr�Ĉ$����Tb	,GAEqƨ��B'k3J1�� �	>�y�)��B���a�5��@���g!S�}XxI����#��X�B��3O/�i�xLd�<�,�Z�!����=�o�����D�1Ҥ�5�h=�Jʇ���=����f�#+�q���z��k���( �oU1hU;�O���;,�z�51�26K��~�X�4o؊�4E%�f��y�$�r�L��=Ŗ�s
�G�u�����;'&&����=�-/��O�~?_I��V
覛n��p�u�t����vsm�*�4Ԓ�R۹í�>��$�iB�Νg;ݳkO���$��b��T�g��:�L������x=���l�������=���X~4�o;�Ђ[�	%f���ir��H���q�y��Jn-���pϔ.�T��TR`�P@��4������T��6հɕ�DBb� �V,x���ʪJ .Ɗ����_ES���a�Q�_U�E�];	�H,"J2
H1��Q��\��ɂ��f>B��C�n�1���
ˎ�q�(�f���f́d��:�����q���'������jK���&#U�m�q��*�R����KQ������y�I�Pd�T��^yR����Aa4��?b�����x�x�q�&��(�i�?�G�E^1E`(�>�uR���&'M�a��rȷc�J����Q_*Z�z��
(���9"ƒ?n�b�r-�B�Q�x���$'�h1�؈%mnn�X^^��s���Ɵ�����W\�Ev�N+�|^s�5{?�����������v���t��<91&+���9z��(��-Ύ�e\t�E�ri�z���"P\mI����C�6#��� sH�ܐ�~���,��r�34��R#�n��EV�[S9A�^II>%GhnzJ�P��薗�ep�X���a)�`s���� 84�����E%�a��"�M��R��d����D��X�>?�ڀY",���0dN��|,$	޳�go+Vo�J
�C1�u����TNa�%~�o��*I�|����5c\0�y�.\��ŋK�k<�(&>����K��R����4��(1���(��}��8�'�( ^�Ң����'y�Eyq�{�Q�QЁ㱣�B}�{B�����4�#�Θ������$�I�C�j�՞ZQ��C�N�qZ?}�1
k�p�$* �4V��������d���sx@Yk�\�g��l�k/b�/��[n�re�/�����!0��f/UU������={v���W?�=/}�K��&��N������o\q�?���OL|G��˄C4<�ӵbI��R����=_	^($A%Q1�4����ԟ�p�yʃM�WߵJ��(MQ�C����`T?�1�^@�xYt��)L�M@�q_�hK�6&Y���j'��N�"�v5M��M�{>�`_���N ���ZC,�3^FY�i`�s�Qܚ����@5��R���Ҳ!��>�riyş9b.xNQ$|a�ϦeM�(90�+1��rH|(��i%z$˳4Y�`�	s^ދQ�����:ɍ	$˽'����VÎ���s�XΏ�>��VD
�k4$d��8S`�ȣ@b1 `�E�r��m.B�	��gȹf&GPYb,Q�wc͔��a�+�Bǅ���\.H����뜹:z��sR����Zw] >�bI�*q���1N�D���&v�uw��V�sӥʆi�$��U<&'(�9��qi��;1�@��)�(�j�g���y��=��S	�:��spia����į��_��_>�i�Ջ������w����?�ݫ++?�괯X\�o�(`����,��G������Tܣժ��w��8�,S�1��& �C�J�()9��
{.��'d���98���#c���h��`���E*H������0�ͫff��]�vH����ah�1&o<����Mq�(�S�]a,'�U�4��O���'�A$�~�B��O@���Np>s�gM-���9Ϙ�S.~�
�Gh�^�"�9$�<�������MJ�:��\��1P��B�:�=����P(�ʼ��xm����@AY%��{'�%I+�Q�759!c�������7������]��x��%=�9��?�/
(�Gͷ�R�|�1Ϙ�V���Ş�@P<4X�̝	#$`71�J�P��U���2M�(�e�SЋ �7�����m�=��o�pZ�u�5�W!Ŏ���5eU���E�m��y��o��(x�����פ$O-(���ŵnw��={���^�]7�.ă�:-7����|���O����_X<�/V�g���pBS��t6��M"hj�x@y��f�S5(0�����1��@��B�e�P���F�%�/l�6_/���@>V�n LLO)�던M����E	�j;���'L�$�q.�	���@�ʌ�n�$/���rߣ���Bk�t��s��.����<��c;�k%�����T�W̭�e}?E\#�26���t��8�7�����D��w�M��#�
�b�zKs��@x�KZ����|���DV����S�~c��1;WMͨ׋-u���z>��+q���qRJn�k�(} �{��� ��{������3(�1��Zy`�k=ϖ5ЄF�����O1�3�
�/,EP"�=
��vխL�W\�$��d�R��3�s���x�Q�2�񺦥�x���-Zǥ�T<*�p���������Xr�Q��^wL��r;�5�j)ƓrbxFĆ"�
�⮩��w<�O~�O��O��P��t���U@������������s�v�Wז'����sF55>Q;~D0�l���~53;[��������ĵ�㨃�%����d	��h�P��N)��Px$�K*�2�����f��zO"����N55;UM��&!�11��
�bٖD9Y�X`%�M*��e��ù�̉ŭ q��cEB�^Y\R�nb=B�[�9&
7-}�se�Vz,���Ba�ql�;>�o��I�廉�2�0    IDAT��<����'Є�@)�J��s�����d����<g�ϸC`.�H3��傰�@��R�履@�d�C�g��V�%�Q�U��&�tXZ54W����=ྉ��C
�G1�b$�x�ļ�;��6!ŀh�_�!UU"�0_y���V�6ނ*r�@��dEĞ�E���y�1.1!��#��	�6U<P*�P�Vg�ⓥj�g�e�k6s��ގ�B!.5�A��G(��ﾻ~��t�~�9���/|���8�V����;�+����{�3��L/���u�* ����|���G^1��xss�� (�IS-,�����g�.���: �*�,�,(Yx���ðj�q�Qʤ$��7�R�y�����|�R9�U[n�P7KQIUy�%��v��b���w�oF<��ii�S�
krjr�l|o���i3��JGƞa��*��R�ד@�\�2Ă�ӗLs�@,(&Q����5��I�ae�|���o����kM=�~^I�"�i&��`�5�D�=�"�#T䡙'_%�ik�z�YF!:���Ey`�s��d�7��|�$��=��X��d�O��'��8_�\#��BA�nG�צ�:ޱ'C,(���.c��!���:^�,O����6��H<�GLP���=>����j�?�?ӵ��C�d`HOSS0�׍wC�ӄe�J��Cw(���`@{e�����S�;9�!HL �Z.6^�@�SĈ��q�Q�*p�n��872,Po�n���~��ߟ�����_�r[٧��V@7�pC����o�����;߾�����,x� ��������
���?�|)*�i�tCx7��Y����
H��T���H��U�zĞ�<IjL�%��$%$k�g(P\3������@Ύ6E�R��$��E2
��aũ��� 7]�^^�w$���rMƇ�A�6��-�QQx�#�.p� ��F"cN�U�G6��$6[�g/�+�>�$��TJQ�MV��&��y�<MI��{�:M���1'���<7^��xyމ�`�D��pa�)�\�n��R3���˹9'�E��}ړU����y���&lƵo�0��q`����3�{^^��K��Q@^W�:/J�ω�'&"�����(�ŬXݬ�zĨr5{��
w�����a�O]GZu��༙�(y���X[S���?����ɠ�I�z�b��.�^�����_jm���6��J�_�E��(ׄ	�c�Ć�Yx��Ν;����<淟��'~�E/zQ`��N��
�پ��kw_��=������孶��^`6��p.��L`c�;s�XqaK��	\#AWh���n5��±�]��1
�%(�T��æ`s�a�0�3�Io������e����0�:j
�!F�����ELI�So��Y+�mb\�l\'A`< >G��c�6�WVq)8
�ͦH�ny3���|Pr�^�a$6��麉�K�Ik��HE�5-X��4O<T�h��K�J<4��;����5��lz+��(c�	�Q��k���%J2ރ�m���BVM���X���k��3����b@m��ql���V�߉b���2�@�Tpbx@�����mC�yX!Q��5_�G��V'��)7[���'V|�3�=��i�4��{K-9�/խ1���U*�:f]��c�b��܁���V#Jv6?�Q��@t��1�L���i궵��Yυ$�~ѫ��Bl��F�i�\�\��M܉�a]��P,w�}o��/�⥗^�=�ڒ�懘��������?�{�����}:�{�rZ�W@�������C��{��{��c��%��M�w/]9I�jW�?��Cx>���䒋� 2AU�e�AIvC^��R ��Ɏ2LS,��A��|V}^�������'Ă&=�G���YM	N�'Դ�I0��V\�	�!-�?�̲1ܦ�-*�;Wj�`��i�j�cnN
�{ւ_���rs
m��$�i�ž,�9c]���K>��#T�8h����F� ��9I@-/7 S+3h�Q������>O�O�\3g�k3W+0
=j���2ś�<y�y.�Q�X�n��yQ5�qǈ�h�� M!�,eQ�v�W��@���kE��t��{̹������FؖyM]�g2C`�o�W�E,� Jl�x*�bz��b�����H�u��Q��s��\��d�C��/ib>v�d���F��6��J�	�r��y2�	��P����T57M
�zS�/#Lˤ�"�'ʝ1B�	���f�fO�3/FK ��}�s�d��]�#�587�>�{�A�Zڽ{�����x�S���׾��|9�~:|��P@���g�������'��筭�����Y\i���di�`�4�^�� ��X�,�=���T��hT�`�F�J�l�(����FY;�����h*e~
E�	��B\/�U"$Pn#!NR�H�<۾N�; <6 �{�L�>p#?�r��`�^ ��b]�;���g��bH��J�Rq!�QP�X����3�z��:�g����#���lnQ&�dSqͺ�&��2�DI ��Q2ǁI/���W�r�=��|��`溬�EA��(��Tz��㸢�;r��*1�x�k�������R, �2�Y �@q|�{� ȸ�Ƹg�D^8^v�GCAH�Q��@Gy��X�%O�(��c�S%iE���b���z%��D�/Tsap�D/�� �'i��t)'�q�IV�����p��Vm�o�{��p�]H	Q$�.=�\���������ڛ�g���(sy+Z���6R�:v`���T^wJ��H˘+@0g��V�%��k�Jϣ;�y��)�e\��u�zy��^sB�$XoȈ��Z������<���������L�Ei�����P@<�뮻f�{��_�h}s�G���/��1A*��z��5`:����l��Y�]tau������֬�++5Hi�]Z_:B�1$���Ve��#6㉅�ژXuY�@^X�ҼAFd�T�|��4W��cR���0�ڈ�4�����R0|�R&��DA07X���^`�p��Њ@�0l��0���*���	����	�����slG�C&	�����8Wi|����>۹k���ƺ������R'q"��E�G�4=�?��ܳ�w!��{����{澚�̜C�/�\�(yE�bx$w��0c�F�1�xyYCM�u#0$�(��>�����,�-�U&��G������H�ed-�qO��B]s]�i����2�'�D���Ѕ:��s���]2.ދ�9(qKߡ�A&*ڰ��<y������(��R5Bk��y~��-��i3��A]��F�k�q�i�r������8(��3��ܳ{�r~�=�<)���G�O�]Z_߸��s��o�|�3���/~��[�x��������c��_^Y�7�V�l,��{�����C�fSG��jX|���Q@g������j�PXǀ*CV�t��:��?Y��Sɂ� ���Y\^RLhaz�sfl��<!6 jkF�Kp���(�	M�J�D��*$8+ߞU}ـlp<��l�T3FQE �;
(��yl��pm�ܦ�?�I�X�͍=�s8���O];�L�S�$$E\��1��%�� �tlY�5�U̡�-Gs�-��s��E���b���~ɤ�+Wg�8g(���؎�Ψ.�����4��:�7FG���HW�O�ysm1~���E��R�]oK����h-ʁs0&~��O����$'��CЪ:��D� +d��U����/�q�A�����s䜌7�OP��\�0�]:G(�6Ŋ�^�L`Y�L�0e�f>��j��w$e^��̍�P��`��N������]w�#���s*N;=Q]x�Eb��Ͽ��/JAEN�������mSS����=��?��?y��JJ�a���󆉷���O=z��Onnn<����b��;�,m���_�\�c����^P�۷�j�F��W#8c�l��������E�߱��hY�(��G�k��,t{;������n:�������C���8y
}�{��$L��.��ː�XČ#4��S�~V�Wj�|[�lN�*7Cl*�(j�<�ܤ|�jhrB��6!8�,�mCY\�d}XW#�cu>T���6z�C������Ez>!;�M�P�(�>�����f̣_�������p{k��/�1ǈW�H�߄�1�����#x���G��s��U�u��4AS��3�*6�F�P�ݕ� Ɇ���%S��4��(��א�G|��<����^�L��z3f��cA��7��	��Br�:e����Sno2*�3�1���\��RVRg��Ӕ���%�Z	�W��A:U����b0�8r�.������\��ȑc�ߣ���S��LOO_w�Yg��K^��\y����J�����a����뮻n�{��g�Umo�juu��^o�E�&D L^ZY�C^YY�zc��
��ݻ���@��T\6ld�&x(�����X�Q����t�>�����vu�%���b��2��J���yY����Ѣ�dS����
�z�]���x��������P
��I�$젦b<���nK�����+:coM��Ĉ��`}	*s�/b�/ek���s �<U�ê?ܖ�bC$`��&�Ch�P���4¨�9�<Ɓ�d#�P�p�l�x( � ���n�ƽ0�5�a��K��%ɑ���O��k;f0���4��2��L���Rk�Q�:��Qj��/s��PX�σ�	J2ė�7���i�VJ_?^Aڀu�=��'l���\3����9n(;^O�c��֊v��c���-�{,�x*B
��Z�<�3��vݧ��&$�4{׿���a��
��c�=UJue<���a��>�dRb_�����3vT�{��V����!j9����233���������x�u����y��W+_�v
�[��x�g��������~��K�A���c�)B���Tj�ݩ�?�1Յ�����M�e�� "&"��E�T4'ǂ���q 4%���n,�@�"��"B ��<��U1�dя�ȩ�V�Q^H�	����.
��:&Z����`�����ML��Q&��QB�>�1�aO g{�f�� �4qМ�a���^�V�uPb�!���;z�Q��Sx�n�$,��撆{��FA��'0��C��k�8��oY�q.	�M�ŁiC����pl�z�����ɚ����̽��*S0�5�{��*nbf9'��y0�@N|�*�0�P�e��b�;uݺ܏����w�f�>����H
E6�(�/c��bKIϸ��K����y62 ؋C^����>���.�T�<���s��}r<���(���xDQЩ� ����g^b��2�&m��y��T]�k�K�^����'�Hb*��o����v�}��핯|Ż^�<l���ɇ��o��\���~�O---=���I�A^�S3*�Ȣ>t�"��Z�X�G��.:�zqa��*DB0�����o,�թ]҇�Zp��#$�tTMB^��H+���pS��J�QH	)4�gf���"�,z�u[]�0�zdC��\�߁d*8�{RBe�J�)�j�GH2��UXu)�/����΢�S^&���;l0�	E	bj��6J�� x�&�G����V,h� "�S¡��@���zjC���;1N4��v]z�y��!�5�c�8jɝ���0$n����.6�-�y}�@�b�ǃ�&�^b\(J��a�g���C�p�X�0����<k���k�T�8�����K9��R��_���T��X������l=�Rd�6 ��p
g�g�ikkS�.<_��*4�MB�g5�|��d,Q@�z����ݬ�n���Yi]��FGVPL�p�.k�.�P�# ��<)��꾱��k�����7��M_l=4�)~�~X* ��u�]7w����6��f~a��'zs,���~EB!���:eޏ�����+
�~�="%P-��X�]���t�Ƀ�G0Xh��c=EHh�v��p�#8m�l	�Kݸ�~�A}�Q]C].%3>f�@yo���:�>"%WlŶ����[u�;�4����є|�Xt����M%ĸ�XZ��3���7��V[)�;=SM�!�2^��x���w�SP��P�E�^a�5�<;,v��,`��VQ�=��x�Qh�@s(�@�QBYR��H^�DbG�U.���g:y}����e�v<�G�彜#m���2��I�d��9��g���۩�#�9^��M����(��`�"��iNt�Ĥ�����O��0O�5�N�@�fI:zJy[��x_P�)V?`�&�N��(�x�Y�|��R֝sg_����j$�����w�=?�J�)�J�x#ߧ7ޭ�8_͞�����v���{�������+��Җ�����U@<�k�y�9����5�����%]��eA��gw53��Z^^��=^��?V +�Г[uV2�Y�c�LVWM_�3j*"	�bQe�4=w^;ȕ ��EaE��Ř�d�#Љ���."l+Y^�t��;,jA�'���[����k��C)pN}��Љ�QNA���J���̞u�ģ/�[�o���x%Qn|��:�c��NNy^����X0'��0�ߕ����*Vzq�&�ԄD"d<������r.yr��# ��s��ܒG��-��/�MK���9ʚwp��@n����m���xt�{��j��G�MH-[�O,l��Y7�˽7�]b/"N��f~�x|̨u=k�c�R��)��=~�Ք
���])Y�/$��_������sM)*H4��V��s��_Zi��R-�R:�A���ބr�2�1��7bAi8'DPe5���)M�D�q<�n�n%��w����AK	��}X�:�|���������?�k׮?xֳ���ӭ�����V@Lį���.���;���z����)QTu���E����{��%c��fEa�Q���d�#��[�;X��t���(���)�3Hµ`�#���
J0�-�R�91�Č�0J��,ˆmw�2����OI��*v�=T}Ւ�f�G�O2���jZ�\#�A���)
#�H��E�il�&�@�����0a3�Q2�VU��ݞ(Тmo�	� bCX[7ۑR�[���斠;ƞs��DqmTe�Rg\�*�;�'˚��1�6���+i�.�x�Q:�"kT1����Q�"��FSI�'16ʸ�f��_�G�øL,��k�>6��|~��4�E��ѡPBx>o��[^�n�0�V�Y'�3��|(2�Y��y��k�܁�(v��!F���	1@��A6@�ά��A�-c��⽓��8ب�v��|�s�B{mm����i��DH����+d�0?w�s�෬������;;��;�����?��?{��z��z�+�{?���7���>iyy�G�O������R2�c�[v�J��c��hH��A�O���_,w~�d�?T�$�C�Ϧ@������;?���(�( c6B�M�O@�-/����rt�TBl /���{Y0�P&���f���~��y/J)�!�(��-Eh��s	�E]7�7���%&ؖc0�+��R B1�0#��(�!t�Ғas���(#��A���ՖA���ƒW�>u�J�ZC�Eq�j��Z�7�����:���u��;
�kE��(�w!W�c��k��0��=3>��	��ێ')"�$�ʺY�t+)�����z�yU�7
�8S�ġ�M MƜ �cG�z��P"�8�w\���E 3ڀ�>b��h�'/6
�c?��WC{&�sS�[P۔s��~���}{��;wX!����}��X��J�����#F��Biː�uQ���[!��M�Zk/-9�]�`�v��\rI���R}������w���;��u\�_u�U����]	�a�z�+ ��_]s�����O����_�����n�;[��7�eW�w�>m�t$̂e�����G���	e�K���O���/�b%� � �w
3L�YIV���l��TЯ�@5�lDM|м��e�=�8��
��)�� ,�@{��G    IDAT�L8>��߉�ȃ+���r,pf�}!�⼁��.l�T�Kɗf�1X�\�J��N��(�8�]��\~s-�oG���~��;���1��5$V���P�x��č��'Z�"�EF(q9)`�ᨃi{��f���^��F���#`Y+��vԥ�x�����5�|OJ���3>t��|_�-��
ac�׊���3�I�	
GD��=sWO0�	b�}n�n,1�(6����[�1v�����e�ϾorL�����>SĒ^#�Z�x�����wU������%&(���zc(<
C��-�d�w�{���ު>^6�(UE�kb?|��������&�T���N�cg�}��Ӟ���K��/�;
�	��mo;��>��.,.����������;]�~zfN.1��yyeQ.{6��Ņb�ب֛��!9Ci!�j+��
!�ϲ�����6	>��%@s C@����
h�){�k˚n�`m�6�����w�ݪ�.�=�A�9�2,U��g�<���E8�Q}�zZ�`��t��P�c�K�no�Ag�W�YyS���:�+����g~R��p)��(ă��v]�3S%�߼���ܞ��w`�3
(
�1#�Uu���0�jQPJ�-;�X��"\y�a�IQʰ�g�c�;V�|"C�����RL5�G�R����)㡶/*[��n,�$�G�G!=d~U�x^��_���u/��x�h"a����YYYֵ��*��P�ǆ+Y'̀�~��VX�צ�ɋr�ǐ�J{[�^tyX��w�VWIT���D���Վ"�k��S � 쩬�%cb�MN�!���'J�q��|-�!2R;�|X�Ԙ�8'9��V���>;1�{��W?��/{�˨��=bO�����⭷��j�^���u�)�^W��� �1��ڪ����i��1Xt���!�\���oH�@.�J'Ҳy���� ����ȃr	 9�ce�olRtJ2!�]�E��@��Զ�WC��T�R�
��r�]+�"$v�u�N�,��hař�-
+�[���!�X��C5bZ�q��0sʳj�â�n8�	��C�=�(-��_\�s�r\*�����A�$�F�������3֍�P@p�@�lB�K�
]Y]UM�x_�E�S�X;nU]<[�9��7�z���xN�LK��f����HWW=�-ӕc0E���҆��IB@�[bIڝQ? y��ik��T������[�zMH��r̦r���%��=������V���!4a�N�J�O��چ�@7��
EY�5���x<Q@ڗ(�vG��9���o���.�@ ���#GU��z��y��5Cbb⎵��w_}�3���W��]{�Sn�������?|������V�����%����"9R=��5�3��F�&������Tx<�C� �U�m�������/�M�8D�@����L\hqy���BL8r*o�R�6Kɛ�5�k�8����`���mb�u��|h�"��͉�����wl �������l�Z��7�_���C���4�70�ZI M,kei��GX�Y�܁3����N]3J���AH���+�2]���.T
����dT��i8��P�б�gyk�b�Ҋ��'.�U��CK�EP?��	��	�o;�h�{J[
��}É��R���Źk���|��')���[���Ҫ�H�z�[��7�#�5��V�Q0آd���pq���ٕ{4�����8V�D֪�g'��3�E���}�������"���QCP���.��}�� t[j.f����e���˝��S2-I�M�[�a�^|�ɖ#GU��u��T}�ـ��ڵ��;v���x�篸�
c����#J�<o�ᆙ���/������姍ML����=�x��8/,T��s�eb���!���K��[m�ˈVh"EQBQ0�,,L}�P�7���4���Eiml8�om�Z\r	�x@o�������3����ZA�����
�!,;���̝�Z�Rɬ�5���kb�2׊�:r�u��������Q**:
L��^���I �r��Y)�-y������+�;n�A�$)�r���X���ư��B��Q�:97�e���1n0S�g���O[�Ą8.P_z$e��',�x
�tXW���܀�\�`���p���1>9�VT�X[��(
[�k�l;�q!è/�����<U*[a��?�ψ��aa�'�	� 豐qk�����Ql<!��eK�����b������q���,�"�4�0��N\C��l<��Q���ܣ<�aխn��6)P�S0d���%D�~�������͚���v���������7?���^x��q
�;���kw����<�������>�H�,l�s�ݯͳ�`�Yҁ2X�{���?�<q�Ib%�*]6�j��kb1�Tq�Q��l�f�)��I���/�y�/���R�&��Wu6}�:�Z:5�R���{�4�B,?���d�Nj�֘*r�'p��M��66����hAЗ�7�)s첄���l62��5Y�w"��;�灼��d^�T�'����s�j���3�D	�]�v����?�R<��������3`+^	�3+��ĵ�x��c[�bi��xl� �=�PmD<>2Tx�&z�X��1T���ٮ�R���>J��G��(��w�Ε�� �ԕ�Y`��=�hA߭xk�M����a�%6�x����Rp7s����C�F�|:.�cvG�:��s�X/���b���z�uQ4��#2q=��a�����|�f/3��>�"�o�u���$�����<��������z�3������c�$�#'�vù�w��g�x�/\X^�����ݩ�!`�p򂐀P �*����hP��Mޢ(�A����Ž��Da�廉Ȃ�7Be�Y�J��p�Ҕ�I��J�E��P���y(-�n���	h1{j! %�#)q��(�!��s�.�48nzzV�@�D�v�5�:(0�r�� pMC#�3��J����x��v혫f�Q"n!���� ^�TbkK���s�?�T'p�cL->�'܎!sj�b/�����11B�M\�c�++α��Zѯ)^Sh��EYr>��A؈�x��L�p��8�b
���T��#��*6��~K����r5��b=E2.JD��3��]b��3���Tnd���QTb&���c>�c;
)B��*x�2�@�x���»��e|�<�q�\(ey�wHq����7��t��x��~B�qDg�$c�F��#�=z�X����CG��AÄ�#��OaB<{��ƥ�������ë�z�_��G��������7�����7�l8�����E�N��`da��}��PY�d4S��D%�`�,P��pz���,LeIo%S����rCE	�J���u�l��-�~bFIq^'�P(��8T3n����'��Ͳb��=�G��du�Y '�/Vc��s��v)ߟ⑌Y�PvSi��D���m8�֬�P2\C�y���'PA�������Ee��tL߅Gca#��n��H���R(�+�b#%Vb�YΓ�9E�U%��ŋb�;`�('u?�r�S���T�Xƛ
�l¶��WW�&�Wbay�<�����i���)�e˄�ԸZҺ)m�?6���^M�Lk]3n⟉3�5s��Ƽ�1���r���d���'s��{a�1��E|���d���2��W֔�no�SÀa^�����gt���T��/��������s*ϻm��T@��K��R=FC�����;�Q�N���q<c�>�3�><{PU�@��z뛛���;o��o����5�y���TG���n����7�|���s?����݃��y
T��L[��3�ha�\F�2�5�I
g0�Oh}Â���w�V7��%��Q� �+���+�M,%�*�ZX�����Vɓy�$��G����#�Q	�Zq�7(���Xr��I��n���R~�2ˎx��y+$�[%،��f�a��9�P]-�0�dM��Sr�]!p�щ1�޹K.q�Te@�"�Q�XG��CP89_��CKN:S���\;�|r�l\7�
����T��	ܖ<%�Pj��i�mI�68W����=�=I��N��x�Q�ǅW��`�������B�����DoB0�7�V�E(H�3v�x�)Q�T�V&���X�-}���x8��ƐB��f,s����I�>>��ZY������=��g�qF���?�iU��;��@��R.����MP
􇡆�!����� ����.��$U�>����̤��N����vn���|����������w>�+|%���V@L������r�đ�U��U++KgG��YP6L��Ў�8�M�r<����#0��L�|G��Ԃk�o5�TJ�D1��mH�k"lQ>������)�)�^Ȩ���Vjv%�C�Q<�x�V��p��x��\��(+n��C� N!ARJ�KO�c��fP[��>dеaX�1z� <� w�ځ��8�A&�F-��L���0�7ccN�BA�J�<S�we�E]�ځ|�/�_<4���1�P�
Q1�BAg���V�[�|��yN�c*��Y�=btD�����
����]-�-W��C�qf�Ļ�G�g��k%�NM�(���I��J#�xG��㹦��I 6����'9���ݖX������
�?KuvvN���J���⦇yn��m�=Ŧ�w�o�&r�{�4���޸7ƌG�!�}���~04�\__��;{��5�wџ<��Ͼ��}�-�G����x���w�͇>�ͷ�u����[�����֨p�j�u�RA	��[b,P��}���o�Ǣ��6�,$��Yg��b�2p�Q���æ��{�wT�:m��:An�M9[�T��P�(V�=��%up|(!X�t�$�ނ��(Ұ�ڥT�Xu��=�O�@���<��Kͮ��1ѓTY�(+8Ӝs��L����B�+��.��=;��!�K�q#�\�n��\Y�J��"�3
�%d�g���u\FC�!̹2�T�HcC+�1d��9�gƵs�����yk�/O��"�Cx���!Q��fMX�v佯���<�K+���Z`�/:k?���L��ЌW�Y��V���K�1�qh*q�w;Ei5��P���Q�9�cE�b�^���%r-�9�����1�5@_���m2)&ʳ���b�V֥=C
��I�����0����8�:CF �3S�����������u��yρ�����{�^���;�m?���T��}������G}�`�b���e&�PV.J�ł�ʦBh�rO�,06*�F���-[��K����3��5�&B���6<EO+f�ܛ�1.�]\?e|b����2���T4r��'�����L=����6"u�bŪ�q�a�ôL�w�9��s1�E����Η�\ ����ͱx��9��QQ����b�'�C�%�SX���5���oJ1>�,�!��y%a�Ɗ�-��l�l#GU&��EW _��X3�ɾ}g����r��[��(@��%�y��C�����A\���R��w�����,���B��rbL�w?��s�sQ���s	=��p�ا�G*m�xl���T�c{|[�A��p����I�x�"�s����n_��ϕ�#A���c5�\s�*ރ�ŋ�F�1>bg�~~��V�u�\����mO�痽�e�~�=����k�����|�;~��+����j��L��ȲA�! ҽ�EƦc���B�EQ8p�*���Q:��P$��c�1�7�M!״Je�%+�$W%r�p"���+ ̢�²|��s	$�T��D���X0�o:x��S���
��=	�|?_���)`���Û;�X�$m2�P��n<�(!Pz�s�	���<�x �E@.��C�V�0��9�0w��x{��	L5;�C׏G����µ�������kku9'������Νg�lʴD�q��q˱�7�ؒ1!$�����(6���F��:�kŹ�� ��J7��j�E��&��=�^y�9��0)��D�o�K��t�R�^�T�+/�zx�T�p���K^[���JT��yBRT٥E
J��������[�$>��{	��	T��M��cM��ٷ[����H���1y?F:DF:���?633�?�������G�����
�!3=�����.,,��`�y�әIL �vǎ9Y�ll9��*�,l< ������A�����%�fs2dд�ORLEql<�(o�Q��)�!~�3�=�'���0����EC=����'l->��m(#d*%�2���gd�#p�U$k�[uӺ3	���ƻ�:�F��d
,��Ṅ�fCH���<�C�3�c�� ���ü"���'_��qʑ���d>�����2F02������}��	Y!PW�m�-�B2���&7p��xd��V|K��:o�;#Tmb �1{���R�(Ə<Ͳ^��>s5�x�RСW��{���7Z��3.D����'LK)��;�W"��&�@��δ�*{:��(��9K�^Uϩ�%fk)��O1͒V���ybl��1�[��?�d��D];sdVbe��ssso{�s�s��_��C�p���T}����w���\����������t	�u�~:��) \O��r)m�˧7ȥ�^&�^���Ɇ�*nn�&�֬�ۄ|�w<{A��7�-�b;�'�G���K�'��7P��26��7���w,'�A�(�(����J�������7�˱7�9A�k g������a'������pJ�g��̳�^�M���[�� ��Ʋ�9�����\F�׈@a��Ռ��9�Z�+C�1�\/�Ap�Q$( �?�%��2�H��K\Ɣi��tO�B�.���
h��q��q���҉����3�sL;���J��(�E��й)���8��R�iT�$+�Q̦n$Wu#�F�2���1��9�_���	��u�;����!(�v)B
{��~jj�x�?��������<�C�*��U�>���s���λ�#���`𒪪�j'������=CU����^��ذ�X8�
.ʊ,_?9.��A�Q���VՎ"��Iu�(+P�`��(��ȋ��WyX(�[�+�t뒘��%���k�8?�慥�}%.�{Rx����w�5Ǉ�!�[+6��Aؙ�l���A��%�a8�����T�<'<�υ^��sn�ၕ"��p��)Z;��Ŝ����L���G�3bе���l
4�ׁu�m*�g}E�'Y�Y#9V�B�aHP��F�|��iOQ��� ���zrL�x�����E������G`�2?Z}����y��똎I�O{/��� �k�YS�I5ێYє��%N�����Do��Z���db
��V^�z�%�Ȟ����ֈ���s>|���X�K1������izz����ԧ~�}����yD����2�%�����66~���\���&�,H�����gi�;v�0ˆ�$��b ��Z"��� c�J4��VZ,̰�� �B�����(�@6��ʦ�g�=�3A��4�iṮ�7{ƥ�CSpBbC��Lg���5$Ћ��g�E8��n�	���@J�߸c�=%��D�8W�#o�s1>���(!^QB���s�KÊ���x�T*�%A�X(�\Jo$)%Bڪ7�)�����Δ	?���{�o�$Ƈǅ 53oYe��+�=���8ޙ�����ԥ��L.�O߅paoQ7N�:�<e�0��	��#���l'��H1�}y�B�̚���cǨVk�>G�觿�P�mD��z2�<�t���7�-��Pޏ�Z�b�#�G����I�{���ۍ�!�s��j���No�Z��v�檪���g=�/_��W?���2_��U@_ae��Mo��#����7�`��/��ڜd��dQr+�J��J��%ʂG(B�=��$�8GbC,l�Op��&�r�J	��ml��²-�O��s�����9qbA4�#��4�V�*U���LC���f�Rs��MN�`�X�E�F�2t���?�Y    IDATթE�}Wc�͜�����P-y4�w��p���&70��sV2����{B���T�/�e�B������DX��/%��h�nI���6�!4y����s1�(4��9V��-Ly祘`1hH^e���m2��@132Ǐ ��C�t�J���9����}����wH.kK_(�{b���s�xm��qn�?�F�X��C+�\7
�i��;y8^{V@���R4��f�9�㱥��x��G��"�ab�`L��3{��>��/T��SO �@���Ԯ�g���O�u�z>_^�>������7��>��7�����>33}�����	ʇ�lv�^Y�����ذ�A�$��U~�9���Î����X�+d����JI�x|�s�ȹ}�(6d��A�b�J
��V��H5oc�)g2�~P@�#9���v�5E=v�%��be�,��"�HE���$�0��;%�������?^G`h[�lN4�|x3($���3����n�M��s3�p�	Ȏk&�	�0��Ғ��'��s�A��`T�3�|yى�tvU�i�e�ja���i���H*>5I#,L~�?ࢥ�k]=*����tG	́��.����É"�訂F��@m샦�Ҳ���s�vV��}�6#������'E�N4�F8�sZ��T@3b��Z<3��Ϝ4�\��Wzu�W��~�������[�|��_��Ga�� _U@_a�ʆj��-o�����Ћ������\��xb����q3վ�g� '�����#��_J� �P@g�?SV�z����X��!Y��N�\��iZ���^��I�W̅��%6d�J�H���W�E�>���2���g񾼄Ψ�vl���u�T�F�%�p(a��f�u��B���&[>Yr���|�.۲��T����$��Bۉ�xqX�S�n!�9�rBJPoA�v9�!���3d�A����-���3k�߀��G;R�{0�gHm4�o1`h� ﺔ�"��i�`}�ejx��M�-U ٬�(�<��R�)J$�3��M�3	�Ȗs�"z�D�&����2pc��C�b��fj�9&�Ω��p�P��X�O�=Q>1�X@�a/"�cų�M�Q���؜�<3=���o��׿���}��ȣ
�\����7����?~����T���
a�p���)o��"6܌����d�ҍ�φ���kFT�/�5_�
��|<����l�c4(�6؎ט���@h�����i��%l�@>�b>rn,���$����+˾���A�ݶ]qxe�&�Qb��+)%^�}r�\3��b��YR�j8詥24q>O������_{_�$�u]���W��Ѝ 	R S���mI�h[cy�̄a�%q��c��A�����<�
�H�dâhRI� �$��э^��k��e���N�"8�L�D��":��:+��2�y��s��|i���q���� )���pA�!YMz�R�����)3R��,.Mh�F�V@�-������E����Q(�g�>/M�8~쳄4�����IV�W��d�a$A�x��=���&��j{ �[@x4q�ߐW��%��������%�����H �yP`��78i�����RUn|��F����ᘘ���/xH�7�[�DE���-�������z��O��7�yi3��M��o��ƛ}[��>����K�n�˾߻�R-a̰b����pv��.9rBHT�oma3EF���=o�s�N�fG��`���(e<����M��<4���KeA��J�F�q~����	��e	����}!n�դ��S��(=!�C�	5��}����P�1D~`��6�v؆�o�s E7Td�#��H4븺N�D�a�@�X@X��=`�α���Z$R��N��𬠷�Z����P"^�*J@TI������Ѕ
�ׂ���8.��i�d�-@�j�3��#��>�ܢ������X3��D$L�� �^@����9�I3� L��H��yI�-Ȱ$�u�*�\	"�§�+W.9�����<]��}a�j!Z�c�TX�J&��>W ��<;3��N���?n���b���� �׏���	�������{�˭V�KQܖ�狸I^s�Hn�;��/74 +'�6
�4VEd���Y!'l�:+����j��Y`J#�vL��P��|�j^���7��W�ŐW�4BR�h�da�\5�s�q�
���Ȑp��XO���L���r2�h<�p�,+^���p��e��L���!�9��9��H����t|��f�XN�)�艧GД���]���4U*2��0!tZ<��3[�`j����#����Wȅ�=���s��."��Rj���������t0��2T��L������	�L�wp?p���	�(���+�d[���O�Op|	w�����OO��ĸ�Q��ϥ蒄����)�K,R�xJQUs�� <>9Q���?����ww9�|~3���o6^�������+_���K�N{��yU�����fWUޱ��&���cb��eй�IQ$��C���)��p�ͤ!�T9	�`�mj"t�t�i�|�Cz0b8R�m�A���i�Ms@
�j�Rl���ĕ:�#�t�.�	r|.a������@��k�9 ����ca�J	>I�ߨ�۠.�=G=1�?`ʾL�u�߁W��;�(Rl�U��FP�u�u����8�<g^?V�$�����c��P{{=6zK?9���yN����*��WR�xB,X%����9�2��cN�y�2/��n8V6J�==��*?(}�`����@T�5r_��qL�A�� ��7�8!�s*qĀ�r.�{alb�Ƚ�؏��o���f!��̠�;/��B�������p�X�����;���H(�� <$Љ��73�ז���$w�t|<Y1"��<)�x�`��A֜	= z��(��p�6ܲZ5��h�lͷd5o�6�4���q*P��f��;��������f�zm`������Q�>{�>�U���3��l�y�SD89T�V�����C�87���sQ��KWUx:�_!,e_'��ͬ�g�4p;�g��[�!�s���A
<�
^[~5 MÝο�[B;�]�(��C�"ݦj���������6�4:I[�Ea���0��14�u�(CJ�y�����o��`cB���F6$��r�
�/	�|��t��5��f��˭[�~�S��Կ��_�5�F-_�?kU6��2�=���#Gr�Vk��~��/t�����w�����<�E�2��8t���
�7Y	��ݲE�2��j�SJ�sR�]kH��lO��*ۆ���:<�v�^�ch���M�-Cc�c��4e�);�/F]�^?���Nb������hX�($��������z���*���Q+"1'W���L����4�@M	֧L��������P���>���5	�v�۱>����{x~m`��lo��M���P�� ��?s^�~�EC��6�b8d8�<x��er���𾗹�y	��b��	?ȭ����y�%�j$�����D@�[r����NLL���|�3?{�ǲ"��`C3 z�ǯ~����y��?�Q�����|�#�F��3�Y«A�B0�=_�pY���-ƃ��jW�Y�m���BX���#�.JBP����b4��6�oȃ�(�$�S�K^�6?����v��sC��l��t娚q��
�������m��g*;��sC!&�O��Z�.�|';m
�4A��񒕷����ׄc#�G���$<h�j�=^L���xO0�g{�8'��τ�NA��j{,�=\{�m��8�XxO���>L U����޻��T]�3��ci��.P(�����=�}o��4�g/�0�xnpl�`�< P����Ƣinn��z}�� 6�T`{=g�����j]�}�_���������L��������x��?��n4־Z*�~kyyymŴ$�Ë���v�ă�UM���w���P݆n���?Ww`�1a�am@�5;>�A媑zL\S���6�I��$�����n��3�(qA|�Ѥwb�|���\7��pIL,#�b�0�y��� 2�1|�aM1l�4��nJ�=�Xd�_�� �C?6�/si̍�xȝ\/�H�O�W�"v(۰A ��F��!���q3=�lz�$��g*��^f�Λ���P�F޴jǵq,p� \dd8�������W�#�4�DX��|)��� N�<��C�aa��z���%��{�/	�7����t]q�����;v���?����ٟ]{�LǦ�M@�����ߝ晟?x��密a���ysZ��ȃ�rV��yG��IӅ��l��X��ش�t��z�*���s���@\��4h;d+��@�A�*`�\�I�T���x-��m�������'��nb� �\����(��٫~h���@�����G�[w{�����U�N���`s�Ǚs�qH�9�bHC|)��6��ު�� ��8l�N�ǽJ��y�A/MH�:O= ��~��xT( 0����m.��O�,D���㛺1M#q������B���Vz�86@�SS��dx�:]�赹��6m���|������Ç����Ի� �}���G��>��3?s��W����9����}�T(˃	V<����3>>*�i����6HD�ƿ��2��QU�J���uP�yIȣ����|�F���8j����^TZ�BC��3�g���U�����S��^�����1'b����ǲC�� c_���1�n�08й��=�~������� ��&�4E<.+�$FWJ]�X�A��@j{�lУpf�U�L�n_Yy�Z�?�c�4ZzԶcx�^�X@�����?OCf0�4�sJ�G�dW���c����^�bØ<�vW�$�BQ7��'N��3���� ߃x��K�!]�rU�x_��iDQt�X,~�С{�x��O���g?�z�MƦ�]@7`�_xᅉ��{9��W�����r��� �������F���̔ ǵ�E�;�=4T�ۦ��ók�n	�������)�T�rd�%�
OW�+�������0 � �C��
�{�~4|��yR�Y+Ü�4�3��Ƕ�enN��wh���� s?l��)	�We���
4G���Գ$ȠN&&��}�疴���x
ɾ���a;{\9>��a�Pj����0�i��mr�`�K���o�'5�!6�d�� d$}��T@�P�]�9H�ya���&��V�}�R\��Oh���C%3MH�!�M���D<7x� V�7�@��B�F����0\n6�Ƿo��������>������@@��P��g��<��S������h4��8ξ~�_	����{����kW�k�e%��FCl�J�X���ڲE�!�"�BpR�\W�T>�CM�`|n�p����sE�m�ڲ�����h��ǃ��s�S0UJ,��~�����K$ ؆��(l�m�rH/�r���* y��,��1���&�5�=���$��<�wz)�� �9m10��ڮ��~x�px���M�mJT,r ra68�������6�؀���$���B������ _$C���Mʽ�p�=����齑��A�b\'r<�zP�J�k.��������R�|�ӟ���f�n��̤xn��bϨz��w?�쳟_[[�b�T:�m��p��
TZ�%'&�Ю;��ŋ�%v�lllT~+sM�|w۶�򝩩1�!� �`����ӂǤ:�(���p���Uj���{��1z������4L#���;4�& ��M ���>+<�m�����9T���Z,۱�W ��3u>VmJl�!�
�%�J5�i�m8��Y�	6H��rE;�^/����è=�zl�y��AS���86�OS���pr�4i�l��1g�u�O,�" C��_IC�y�J :�����HC�����9�#$�{Hz��,�@ύu:�>8��={�þD(��U���6�1���뺗�0����������_}�G�w��!#�y@7dXӝB�����_y�O�9s�A�N.������k���F+"��T$q%	��hc�°�T�;vJX�avӄH��(�S��+P���@�3��&Î���pؖ+M~�F"/5�)�iPz��F���DψB��K��;�����0���h A`p�JA G�K�x�j�z K
�����&��\:�}�}xF)"9wk���@5���$ j��l@f���5ve�3W����eؑ!L�&�57��dx�Z��:騛�����~���m�q=oG�C-���<;��|fC�m�ڒ ����u"B �9 �� yW�#q�&J�E�[�b���������'N?�裚��^7l2 �aC;������O?���'O�~$��?�x���y�"|�$���0t��������TxQ��W��g�m�z]��z��{Q�C:�0 ��ǳ��0�0X�P�+R��K�*Zo;l��S;�g�$ێ@6A�Ǡ�e�6�8F��PB��>�
J��k��2F��g8�k'������?�� ����C0�2�+���@X,+����4���,2��u7z̴�)���l��\
B�&�r_ b�Q��2�D�H�Y���*��aL���ܨצ�N|�7�6"�[L[��>���1��tl �j��d���(���j��<x��w�y���Ç��z���#�����?�������W_}�K�+�/x����wG����#a����!��NKH!8TeC�
�n&�S�,1������@������5' fb�6�64�v~�^�s�
P�;�GjD�4�4�x/``r?�j��{"l��ojt��=�����I<Q�����v�b��4��)��K���J�$�_���W�	�X��~�9��Āy9h�}�I�FçV;�s�&&��S��s��i�m���I���\�n�y���a��A�"	_��ތ��'�W�Fc{ۃ�=|xn�-WQ5��u|��4֛^�S���%�	��f͐4�!�AEW�(��Z��O<��S�7s�4	��P }�� �B/��Ҏ���6Z���9�o����^��
M{\[9#��l<P��j�ݷF���V�6)a�((H�~�����Q7l8t��0�B��*6��ƕa����b·:��pN�\�SA$i�`V��I|�����Hp`��@��� �e�i�M�@4f��(QQQ1��~@" ۿ��pG�+m�Am4�5#��iZJ��4��ۤ$ ɍ�+
��k�\&��a�9&���m�/=�d;��&L��F���<�A���O�_�ā�B
���T�V"�;�:�;��369&,M��x�KB�N,Q��c��=�X���r�v�]���z���������|����ϗ>`s���Їt|������s/�}���?���O�a��u�"~į˕����`�`hY\��o<䶑��US�s	%�FD�^&��)~��+8q�L�l'�m ��%�i�Q�	]k1�z� ��%�5,���xU� CF��擔"��,���<����1�d{v�	�/==]i_D\Y�2�b�M�Mz< ��_��@�Z�W�a�w*��Y�+� I���H3gC�Û�n���}��p9_>�q�!'�aZ;��-΅^(�_<礥��|C���`jO%�G� Nd��<���C_�^s��@m��g8.@6
b'_�9�|IDa���z�Ғ�@����g�c�<�z��g 0��ˊ���_r]�5�q~x����{���4>$S���Ї8�G���v�?������tڷGQ4�ش�i�50Vz�ʮ�jr4R�-CUT,�զeE�<v<�B�Tz�T�p0i�簆�Ɨ�	��"�a� $��dJ*h��%����]HDP6T�4�S#�m8�iz    IDAT���B$>0�f��I?�.$�2,�����h��\R��_O>�߫GE��OA�u�FƓ��9no�7��ǟ�%�瞜g�ЪM'�44�:"��`а� ��m��4�3uR !4� a��?����	�[�)6I�$��qXd�7<x0�iϞ�,D�׺2��#\]�MH���b��s�<b>��Ap������{��<;;���c�i {}�#��>�4T�m�����v{�þ߿��h��a��E9��7��# ���5y@A��CIE�
c��V�0��	e5�� �����5�К�H{р����_LJ�3z@4�243�-����+��NE=a�b�U/��!q�R)����v(�Ɣ���3�c����j� ��3�~66 &c�x��m��Fr��e�zҳ�1�!>�\�a_���䔤�� ��#G=]L0��#���� ��7�HA�LT���b�"�1a<xD�?b�بÂl����Z]�}eW\M��  ��l��-�;��]������A�	�wwB�9�7���?��ګ��YUkm��_�S���;�p{������^eꥇ-���I�Up����i~����:�}־?k�2hX�3��T�� �d��IVr�$8�܋d�@^s�,P.���2/��`w�77�}�F�Є���`�4����r�gE�P7��bOݐ?X��@Lq�n	�f��5e���/�YT�4�*����`+�`��"s�ctJ�F��X5N�tK짺�}���.�j�E$�⴩�@�E�Z��w4�؄���_M�]���a~]����Q��B
��;R �^]�.��]��؊�\f-~ ���o�x�j�_�q���P\�>:�&^��m��Z�������m��b�� �Oś�ۼ���f	3ƞj��F,�aq��3U���edd��=�*�_{3�])r_u����p>���X> � 0��^������5�>{q>�!?����VPt��+�?�SV��b	�8�E��eT.U�z�z��QR��ZX�	Fe���!���_�R^Y{�54�i��,އ>b�X>3�u��j�q\� �a�T�)����D��g����뗞[,S�qE��ֿmX8X/���a��Z+��67n
O���a����:�G��-���Q"P�a�����bm~g���F���m�Z��T���*Ń{�0�wr��ҡ�&s���,�t�����ɰ�<�/�3K��4]^^�����������#x����V�t���{�������$N���8�+4�c�1~_5�ۏ�~��P���W�T��W��@y.�1���'�����j�Z�!wZ��7�>N��G�&X�KNJa`�q�I��RZlц�[<� ]%A��+��t/�|�ߝ�]פuwwf=�Ն}b��`<�e0HIN�8��K�	.���p����o�-��K�z��T�bt�B��c�GPjR�s���0����ҰI�?/
u�+�#�+S}J!RH��RQ'�t�U��>I�)��\��Zw��)�����O���9{�fěg�(C���o�0I��(��V͆����?҆X��=������"gx��&|�ԅ��/1V�L�W��J��
N���J�)��`ϙ��}��H	�)ZZb���1���*�{#�6���E�D��V����(�a0���F_�1 �� <����x�;ܖ�f8D���~��.abh�N��Q��]3y�m�緲$6�X���1 NƵ8MH�m�,�Ο���b���k���̥ �p�~��ҝu3�4����j�\塶N�׍w�$��n��B��8{��M��E�%���CS7u�-^��mF��9l�����m�nu��xy��m�{�+����:#:�-L��������|�"q�N�����X{
m�\�Q����/����e]~���am��|���!y�����d^���#�޼�"=oZ"[�!\�R����Ǒ�^��RB-�E8$������: ���Tn�}�]���WZrG����'�Z��]Ľ?^�O�(]R�Ph���k�M�Ϭ�ٻ����.Q7�y&���F�	�AH��@h��d��������od@���}s�}j=�H4�f���
@�*��f7G�V?�>�W����'Jbi������<�p��_w�>{�tߥ�f��`b�U��i�7���~}��=�4kՔ��Ѽl��W���������v�Η�mՊ����y�A�
��Er�\!=$F&#,,E�ހc��2F&#�Ƥ��aF�QU�A�1db�ͽ��o&��������-|3#���Ut���x��0�B���l��x͞�& �Ltʢ����}>�)˸�n��]��s�7!.J[�Mḃ+��]��=��C�~���;m���u�a���e����E%U�m�hm8#�be�����j�� (��`��8Hcf�M� �h��7P�Y��-�@f���}��7��t�'���;�IY�f,�}�LB��ṁ�ố�n��bJӺO�B~��ͺ���h�͋ܳ������;�T�sX�� }�'V�0
'��@ 0ُ�B�0�02�Ԭ���6��H���KB��_�c��rs)��̦f��:M��0s�vU����ǌ����Cn��Ñ3Κ /����ʚv(ej95���dg���?���Q�X.�ʀ,`����c�RYڴe@����)mk9BѴ�^Y-��|iK�#p�ώ|��Eܛ핍\U����"\�e0��&�\�5�5�4�(3
He�WC(��֚��u6�ْ�d���6�
���7�wD�AZSd�#�],ҹ��e��FI��������������:߂�@�c�JB�}��0���p����Lɰ�~�9����Ǚ#G�J?K5��|��\�2��o	�@�>��7�Te &�#���j~@7��R�Dz��Mދ"<�NU%�q���*7f�!e�����Qϊ��|:w�2ݺ���[{�ܹ�Գ:x[s,���4#ԇ��:���`b@���E�Q�9��^�ua�� �Ea�8;���8T�)qT�.#��h�g(,�%P�rW1KIF��s��m�y�C�G�
�}�=��uve�
Y�z�t��'���٪��\"� NP�Ƚ��^'�������I	O��SG�mb-����C%n�|	�UQ�������jF����լ�{`�裓�xƅ	��6�����;
�,i�Y � �{x�*�_�Q2b�|$�~���~�}�{Iul��J"TV�X�XogW@&�P�Ԫ�� ����X���Xz�+���T�����UDXW{(����WTEd:R\n�]��`'���zȝt��R�8ǹ'XY�@%�4R�d���?K*1>�J�3��ǚ��4s�@Y` %���c�����ûu�/���/����$���}�9b��z)�r����T�a9���W������(�����~m{�]c�8�J�-��;}&�?������Z���Q@l�I�n���15���1���%�L�չj�Q7��[��Fd�����o�e�
+hL��C5��j��/��vX93��+�}eWi�� &k�$�hK����H4��.���k5�1��Lgy|B���Lg��"��� �fy��%31��0�	�%�}{;��E8��y/�+D�h}�"l��y�	$�7SI�6Nv�1�k��d$���E������N����[�%�}�~�&���_�ދ>��cU�;#��~gs>-�غ�;�����N��>�77�g���y�a1���t���p{�ԋ������9�G����##�b������U�n���[����NHe�z;��� ^o���$O�c�C�2eb�"q�W �\���bL��9s'���0%=�Mܩ_��1g�F4�h�֊�rI�~֪4L=0�1E4�^��R��y�a��b�y"��e0���׫��l��� b��ɾ�-�Zz����3�w���0�6���8��.���MP�ϒ��Bx�
uD`�O@��<A�G9�u��+��0��v��U�+���λ�
N^�>����c���o=�w�u�wr���RŔ��#N���sfdS�k�q$ľ�����]�C�crcy�$��uM�Q��I���YYYi�iB�6'�6�8�y����ɜ�0���tP������{p��,��B�2��}�8��m3�Y�����!�cG�7�>~�E�¨$=���+�<�Ż'X�'&zλ�
�j�*��ȏ�jUL3eG�^[�$V���$���G^�b� 3y�K`_|BU�څ�L >5ǰS��Nu(ZA�~9Z���K��. :�@~��Ś����"r'�Ol΅������K�Zj�n?pC�v6=��?�V������,WWW�w�Bي��7/Cr?�ٷ䤏ӳY������ii��@Ǵ+H�#;~Z���]��N0�#\����z.�x�S*0���'�#�^S	s�F2��k��s�d�|27.�5�M_hԺ7�P�$�h��'y��<MH��"�o��X� �^�Rc�ja����3�t/AA
,� �:���?p)�*]�j[�A�UN/������7V��}R�5�%�1�{ڠ
�.N���xA��AT���c
���"����:�^@��nX{�����Eu����?o���q=EGVT�z�߿�l�j�{�$�3>�9ɍ�	+��J*n��v>c-��e��L��wg��EK��d�s���%�3Vb=�~X���
�"D �bdW��GA$�S/�-���X�eP�xH���gQɩ~��eu%���0��h��-�,�d�`�a֭8!�Qt�҉l9�K
M�k�Sq՚T��qzܺbf��܀��}��{$8zcp��⼨�vB����#�ģ5���7e^�o�ԥ0��b���L��" ~V�x�zq�<�qe��攇�: p|lGr�)S@��
�Y>(/w�aU�ܯ��,2�N����Sw��n~�0LV��X��=���P�#�w�������pES�N[�r��s��{�^�笫hy��mI�`��n��+�3Sݘ���-��1�rH��B��T��v-B���Z�C�R�쟍;"��
D�>�ʢ��|�c$���o��p>�rYG����O/\���Ć��a�&�&Q�|B�`|�,��j���H��ݏ��X�4K�H�C�W$�����n�|r�Z!���OҶ4~���f�x�7%�3]������t���]e���-^�����	Nv��h���{��ux�w��v�Z,۷�9�J�Z_�ר}�|��%�9���Mcc~+�ޞx�� Ɇ�P�blQ{�ޠ�Ӭ�[��P�m�t$�!��j�G_0Q%Uu�L_F�����cNa��D��1,��������=��z��tce�Fsgw�<�h�'�E���!�\�1�g���&�W/+�*�L�b�R4^!@�@0+b�Z}M���rH��fN�2��$��� ������״m�y\��ȁ�N\>�_:����r�q��qڽ��áe�ﵖ��t��b[w������_��խ�y�êD�<k�!]�B������r�����'����8���^�`ϧrMe��ߏO��*���N�����z�Cf��LP� "!�Z3���?����h��0�J@��;��]Y8���T?���B�9�x����4����с���Yq����b.��bz����M���?[Y�
���C(ܷl�F'(�Q��!Ok4�i�@Z(H	��&�ګM���i5���=:Kr�ݟΝE$f���4�O2��X*�5?
q)>�������NδlZݤ?uLk0����]q @�*�ũ�L�|Zǜ"�j�K1F��t�l�s��Yu��!��ha��CX�X�A����K\I��Ɨ/_�����r���6��r ������dU�`ʝ�b�`L2�'�d����E� ��D�J2q�w�h��ϋ�ay�����4���������+�V^ۻ4�j͂葠�n2��q���*����5�'\sR�.��n���;�L��kF�Z���i���,����L�FC�For?k��C��c��#Vf�Y��^��Fg�E��_k�'}I��񇃆�/��4�.�`�'`��3���9� :�5qy11�zU��L���1�z���fq�ɦhs�w�Tux���ӗ�Ќ��A��19�)+!쇾8H���_���0c�'�Cڝ�˟�#	Ufե�w�����
�c}w�xrr��-��ݐG1�~T���~�r�o�� 1��r�Evci��)�S���{:�ż$��@��%?��mk�ؔ���S�"0+�.H���h1�z��+��&sō-v9a|��V@��@�Wx���b���y�7����El��.w��-���������¤(��#\�>G�����}=ҥ�����8s�C�p��d��ٖ��J{p��������u]|�[��_�4�{;V�;�}7�D�x����	���i���е�)��He��:�$X�/)J���
쳊��F�'W���,oV�WC�+�S�0{���_�>�����HR���?���B��.!���XM��p�V$ȷ�ٱ��]6mk�q۳pX��E�����p�wE���y��߶
���}��ǥN��&���̳�1�C�+��th�	� ܍0B��R�K�U+YD 1��LC{��\bdg�������z��/,�~��q�&��%#��G$���82A>������ݧ���I�U�f��eO��6Z����#������Nl��ɗ5 � KĐ����������t[r��԰=K��G"�UC�tV���(�}��������b�4��;���[���_�>�b����2�AA:$jP���\�ںߢj���Ⴎ�f|)AtD�$��-�))4[^G�!W*�ue��=Z�[]��o��_&�����WB�i���q*~%H� ��<��)@��~�^fgg嶷q�&��9����IW�w8,e�$56�0=�QwK_j��l�ӛ��~|�3�f��z�����7�f�:�(,tw����#l8�TY�$p�g
�֢o�`3�_�r~wXDy:�����x�BDuZ����v����\Rh��`fd&ԢRT3�/�T쉥��`@���
jI�
��GӀ˥��܋���D��x�2�ٴ�#�4�����D���O��S���1��FN�M�5s��I5����Xr���XЉ�I�w]��lv'��-=�:Ok22N��Ց}�I��Fu�@� ��������#�

��M��x:��L����9]�:�}��=��X#;�� �!r�`�8��EuGd��1{@�_�������9��]�C��H��B�)#M!��s���[e ���ĺ�h#H���M���7���o�i���O�^��?�����( M,AA�X'b^k'@���O���ɐ�yV�L����»m�j։l�I����Z�YL4�J��k��Sbtq��\׃W%6�W:5\��o�q��ΞfӬ#�@��9^�E?h�,p�G«zxK���r�}:zm"`�:}�D
��>@f�>��TQ���6)�I��S�R������ҕS1�P0F�x��X�e��nY~"\��jc"}j� ���U)J�ۈ����t�)
s ��c�+]4b�X�O���7�Vg����ph�p{Q��iש&�P%D���+B,9q�iZ�J�p����tZ����'v��@г�Zy��`�:�����&5\�6�������ﲄT���߲������ב�<y�����V�.�G���7OQd�u�l���l�2W����x�:�@��03$B�]��< ���H?B�w��C�f{���5�i�����A�Ƞ��%�<]��}���&�	�c&��'��0��b�`�$�x�����#V���l }� Az�_(4+��;:����ƒ�_�3K�@hpE�rB�QC����q�B�˽W�L
.�v~��8�=U--��%f$�$�J�ӥ�.H"Y����h��_�ّsUU�-��[�w�)m"{�9w.���8�LjL�E �B*�L1��T�(j8I�,)?Y/�YW�7]�U�	}�$�W�|�J+F�%�[ P���P��Rc����[L�D��0��p�Bd��,�)l�B����H�M8��1�k	{�w���h�;_��Qr�t�f�WT_��$�pR��D!�7��U��
L���Z���!o��P�w��y��4z�X8���X~eH��;����X�{���α�Y��Μ_�0��$��-ͣv^Kx����ٸ�9o�4�ߪp�!��ˀpMW%Y�1p�I��ݟ�L��~����41��4��{N_1@�di�k��&[���:��Wr?��"Vئ�;�T���x=���E�^-����E�M����lE��+��x�4�����_�~�ͼ]]��j��Fߵܹw�GT�I�6�V��m�=��~���Z�5������ݽ�UPpM���ip��*��Ľ 2|k�{F��ى��t���)x�ܦ��Փ����׮��7yCO�]�l��֫�x�t�����(�ScͥK8�L�'Ƀw��E7NM��E<�k	�E��e��@J�1A+串�S^)�!}b+ێ��v0�� )9*�8�.J=�l�*c⢱r�ƽ�Fqp<�$�Q���qk���]ʕ)�Zc���E������+q0�<G��C̛�%u�1����}�gC��"{��ӻQ7ߒno���Ȯ�������ö�q�� �d�����+�2/t���C1�[����AӨ�&�r��У��(���IǴI�&Պ�a%��l��$�s�A�8\Al#�l�+�jQz�AكNq���+ƅ�P�} �ki�H�>MNo�+�]V
YLF��Ѷ�}2����$x��Li�o�[�dxB�ڮɭ�*��J?�@Gk�VV�jP3g���n+�t N�<f�Z��yS�;������D*��r��?s�=ێ�-Y��5++9�L����x[���݆?�������H��@�ёPH~ E@� ʞ{U�2 T�`|�1&����6���S��I��x'�����c��
DD��c9��{>�ۭ�j]���������|>�k�n�
I�l/�v���+!����r����kz�l��]����*�G�-,l���'�2��t>���)����\/)C:ܛ�D$)�1�қ�;W@��շ�D�%̰��X���Wζ�����}��J6d�qZ�䇩1��_:KTv�"]�	�n؉/�iA�}ҟ�Ģ�.���S
��`�0Tz�zɢ\,S����l$����#+�%G��'�"����[CK�+m���0�n��YP���MCB��s�R\7+/o3��~�f������d�4�7��1��x��m0�����j6p�i�Rq��;��m��{�_��9@v��vpַ��{c���݀CD1~��G����WÏ��g����ۄ�Ȗ����x`W�t�Z��ѨA��ƨ("�]�i��*��d�I���@�����	���&=��৿~�� ْ�?��\y�+�*4,���Rmqp�a�G͖���y�^�U2��۬��S�}#��?�L����5��%����uh��Z��F]�-]kJ�~,����t60i�Y���t��ϟ���M��Њ 7π��}���N���mX�T�e�Eu^�e>B9N(2p�O���B�Ò�'誽�F)0�6z�~<�.��O�A��&��}���rW��ˎ�����Tp�<��G��Fw�d:��ttIHIu�	?~�+�8�/ѢO��{^݇-���N��ƛ�sV:� D����*Vm�e��?U?���Uڻ�PM4�:���]j�-���N��q���K���bH�ڍ:�2��s���=N�ͤ̯�G�!�#�gF'(,P�& -�A/�q]��� Jw�hAJ{Y8�a���df�z���&���L���s�s&	��k���q����{�N���ؔ�v�~�:����v�ÿ�������g����te�� \���ǆU��:�`SY�~�ܼ&�G£|��F����{t����b��#�P~WT�z꾥�'09�Q��G�a'��/�>D%�)���!�Z`�u��'�1�}�׽H��#��!�3��Q����� ��L��Cɰ~����,��]O4444�x�N��a����kVm��}{a �����Il	d,��>��*�j4]��̪j�Q�o;�c�����u�����=|�`.H�&�g����8\�}|�32d��2jR�t���y��V�U�X��Q3ᢪ���;B��]������Հ��G�Ȍ*!����?ѹ��W���o���ʮ�i�v@��u����l',=8�Q�h�k\ݜ.�o^�9�μ�9��#"���A��������}��y���#���y�W�j�����f��%#���V�(� PK   �u�X�}�	  �+     jsons/user_defined.json�Zko���+�>�������+��$v�\�@\��&*S�z8H���e+RMR&mp`S���9�sv�c���H�w��*-�)Wu����}Z��y�В��WV�ܺ��������]����KΊ?qZ,���xop�t3_~�{'��:-�.��r[�7��ד-��#ڻ�r�N&�6ΆLC �iFdJ�IB���6(��YZ�e�X?�t��
�w�R���j"0�	$� d����E}��Ua^?<�LԔ�@L���2�Y�O�� vݹ��a�/��?�_g�n~��8��|��Ǥ�ܝU���}��g��	�%��	�m������3�U`�C��to���U}��K�a3/��UՀ�fMT�ei��p��R)�����%>������<�����Iw|h����a�#񳛭 �/{X ���z@��6�Q��V(9���^�F�8�(�� �^�FP8Z!�֋���A�e�x/�n#p�e�3�?K���hA)K��S���ШA	nF����[[Ѝ���@�~�B[ҍ��l�;@?����F�2c� �s	ڢn� �#f�����ڢn� A���k�֋�5�nUR*;Ѭ���Y*IR[ӏ��s;��<wH�!�f�P�/��� ��rUq��|>�!膪�[5����nm9o+73@�` f/@[����I9��t,�X�Jk��_�Y��̸(���'Q?KY��Ԗ��ph�QJ-�p��k֖���Pz�Ύ��-b����O=�?G淭a��	jp:V�Y[��O���ï��~�v�_|зj���'^Z�i����o	�żN��zg����;!��}q:-���}q6-��iQ�Ϳ�Ol�oh������~dpH��^��&֣�q��(�,4��<2D,��� 	�'�<�&&��9i�"��Gos̽�,�74�ӽ��Q���5%�i	%�\��{���x+<�φ���1���rw�F1�a�Pz���JQ���S辅'=8�Lilz�EdI[��-n+F^�t�Ҩ���Ca\m�����<nfi�r8D�\���G�K,PJ��ط.�3�P��*��h-*
�
�j|RR.��a���Dӥ���F*$+AX�N@`{*��v�G�c�	W��y�جGh� H��1���{��J�G���=�����/H�e�ڝ�!��4b�@����z��:SI�W�}ˁ��ꋣ_Q	߰�u*����Ӭ��P!C
�����9q�"�I���@LJ)H\�d��( h0Ae���a�9$C�<D�ց!���O�* ���R�Si�ڬƮ!X8.�Ocv�~E�'��M/>~��ߖk�~��^�	ħ�]?�ŗ����T�㋁�Ŏ-�= Д��BW��d�'�F��F[F|�E�Sj�[
�o	%�,����"�DK.2����D�،O�KN&�Lc�{��6�V�D���4�%��HR���=u�u�@��Z2A��Sa-�"I�C�^.�ӯ?C�x�مc�QT6��X*�A1��EJ*��ǋ���_�- x��&ه��v�}N�0����Q���;Ȍ���τ*-^�އN���Y��\G�����@Qt9P�RgiZ,S)�
MOJ9�!a�뢑<�~6h�{5ˀ�ZK�X&K���x���)�\�AK��D˧��c��/��1���������ߣ]�ʀ��Ȱ��Xxir2z���.q��tD�D��4���-�Kµ�eŏ�!�����M Þ*�CES����%�L�΍S2t�/(a�6��Lb�1T��\�g�gC��������� #�!���O?�h�� �NG�Cz<����e=��7�P{�U��$A�mV9:�}#�>����(�_>��.H!���Z���ȩ��p����e p��0F��v�3�;��}JW\,�oJ�ʁ����`�b%f�)�Vj��Ȁ�Zo��@�.����v�aL< �}���{�C�0�)�ch��h�$RnxʆX�4v͋���Z%�I��,�鴘V˰�����;?�;s��z�Hۃ���]�g٧`�X����2����e�?iITAY���9����H��(�R�W������)M�Wo�u$���
�����l �Y��F �L�q��ʨގd�U�ＸZ$���������0H)����P.<c<r�4�O�]v*`��h�]�&֥���:GnT�i�:�ج����-|L�����j���'+�@#�<�������:��D D)��4�8��o@�P��]0)��o����Xؖ{]m�}jiϖ�j�x��Hٻ���;$5ָ�#����w:=�A⼦�$����C���}Au����͑꽛m����H���c�������_o���ZU��vז��Vaۙi���՛��z�ܲ~�{]^6����晴z�at7?�ԯ?�PK
   �u�X��j�  �                   cirkitFile.jsonPK
   #aX׋JW9� m� /             "  images/0bb515cf-1352-468e-b4e5-fcf5b4434fa7.pngPK
   ���WX���� 8� /             �� images/2f18dc81-c63e-4164-9e24-83fe71d4cc63.pngPK
   �u�X�j�� 7q /             �� images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngPK
   AaX�34�� �� /             �t images/4ae31398-47d6-4d15-8d33-5c428753ae4a.pngPK
   :�-X�L�,� o� /             Z images/50816f02-2fca-41dc-8ce8-89c3cd37e619.pngPK
   ���WX���� 8� /             �� images/596601c5-6246-4a4b-a4a1-d26711181a9c.pngPK
   :�-X�L�,� o� /             �� images/6b34e9bb-e0d8-4181-9662-be6b7300858d.pngPK
   yaX��:4�  m�  /             4j# images/6ec16c1e-7036-4ea0-ad85-1b4c89c7aac2.pngPK
   ]��W�a[}�  #�  /             d�# images/7a3ae19c-2290-4841-8048-f2fb794005d6.pngPK
   �cW�����8 �I /             ��$ images/7e277f05-db62-4931-8fb6-9134226ee38d.pngPK
   �u�X	�\  \  /             ��& images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.pngPK
   �cW�����8 �I /             _
' images/996ffe1e-7752-4112-9b94-ba61923e6aca.pngPK
   AaXU4Y�- *- /             \C) images/9c0c4208-33ce-4eb7-a42e-8f166060eedf.pngPK
   �KX�����"  �"  /             �p, images/a8d700fc-8f9c-456f-9f71-f71b03bdd111.pngPK
   yaX���4�  	�  /             �, images/be3f368a-d9da-43c0-befe-16a00a90d491.pngPK
   �KX�C��z �� /             g#- images/cf548ed8-d697-4c12-ab8c-ecc45c0ca7dc.pngPK
   �cW���/�� Z� /             ��. images/d0383ef8-9bda-42d2-801d-b77fe86508e2.pngPK
   ]��W�a[}�  #�  /             �:1 images/d19d5e4e-12a2-4f6e-be69-d40783d16976.pngPK
   �cW���/�� Z� /             ��1 images/d30bee40-a8c9-4828-86fc-eff82b5740c4.pngPK
   #aX1ӈ~�� 7� /             ݖ4 images/ee71944e-6ad0-4091-985d-ee04a3ffb0a4.pngPK
   �u�X�}�	  �+               �7 jsons/user_defined.jsonPK      �  �7   